��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|݅o�@
�nI�֛TU�PP.�����+���u�Jf]�ϫ(#��$�r�jO!�Q%y����m����T}�R4�?/䃭0����AU�(�ƾe��������f�7�m��v����of� 6�{�
|)t�]з;�Y7�^�u��]]��c���Nd�e�@Ѱ��iw6���=uC�Q�׾���VL�����EQ<gS�Jdq���<��;^�<[0HFI�W�W05��p*x��$���[��l]/�a�a�U���k�bS���c���;d�#�{7H�2ŋ��J�3��Gqn(Q�¡l��uw��:GV|����J�'[MU��0qZ!��*T�P6٫g"���(�4s�4�f���_���3���=�3|�7�(�n¶Ē��P��ٺRd�Pa��vH�r];4�\w����F�XX��Q�AF%\�#�eM�5�K�5˧־}�G�s���P����a�[�gƉ��銴6	I���&|*�g�(���`|�G�d�q�jz��2��I1 ����׼ܲ�5FZc��V��\�ee�!�"�ĉ."�,�� 5�ݕ�?C�P��{З�wPt*��@ܯ����g�/����u��N��1P!�F��R��U��\|z���;5���d���Ȓ�w�}B��5�z�M�����+S�!�
��$�36%�f��Q�\�b�Jr;�Gn��Ng��6,י�����>9�x.r��u�3vڠ��M���/�f�s`�g����J�9$��6UGV!�ʟ�7�3L긚	*�����i�5T�rY�I���G�ϐ\�[���ᄯ81��vN�	�I�\	��W吟C�!�OQǳ��Ҹ�?��_���蚡�違h��v�|�v�E��n��=�������ڏ��ma.��<݂_�����y\b�V��p�f���E���>8� �t+�x"�ݷ/�]��6?�>"I�R���u�0�����%kĵ���`¤	������e���M�aXy�z����HbG�	������,B��M�G��]�d�X}��H�l��n sPt>����^t�����'^&�.�`XQ�)]�qX8O����O;��EN�����O�"�GCu�XLQ+`Bow�;f5�m �?#n��.EV^���#�>?�C�����̼�}���j~�����KC��W��S��8m��m��V��_�L�o��@Q�wq4ٛ5A4�Y[��YWm���#��������~��4%�v�6ܵ�}!>��(:�F>��ډ[��jLVN������$��n?m���A79���~�@���4s�HD�@߯�����`b�UU˭dj��l5��yECY��G��S�Ѫ_I�8�����Tn��}b��r+��#��E�S�G�s�Nt�1�p7�v%b��ݾ�;A�rŻ@��Yj�-%B���P�Þ\m�������9�wdTHo�)�	� ������&_3�oN��9j��Q|����#1� < _yc�U�x9ZFB>��\���}�q�`y�69iC*Pܩ�(X>q�s��O����Ln���9|��z9��:�u A�+� ~ȅ1��uy^4YHۋ�����4廥�J�?����x������j0x��]@�$��"������:g��t��:9\/���Pn�^$ aQ=xZrj;׼�1pi�Ǝ=Zb� ��JKq�̦�D��^Z�x��V��)��{<�H�Qa��L@���v�浽��o��Mf9U�||�9h
�?D���P����-S��)j*�v'iiP���ej��8�GX�y��ig%I횑�1�m�&��Jfue�a{ڞ-.f��ɇ��OY�WP�g�	�5Ёo��YM�e�Y�����%A 1d��c�#{�g:*} ��7�I\*�����P2R�e��7��*p��أ~�'��w���9��j�^X����Y�#CϿ<z�m�s�ǿ�����'��v��#r1��~�����e�o8����-<�~Z��Аj<F͠%F��]���n��*��;�ByC���9Ȋ��j�c`@
�OR͟�������J��љ]��[�+3�֚cϬ�ǜ?[�+%�rd�ԡ��N��zf�� �ܮ��
i���r���Z�=��w�?="I���tdQ�E�p�\�.�FB�%݋�7�/���Q���v�<����y��,�B�k����6�̣/-�A�����k_"Ij�HT�sA�_6dJ%��Յ�J�[q���x�t��J�ⷮ�0	�Rd�3;7޻:ak���hV�ƏaHA�@�lKG<<F��l>�����\�H��'����^�����h����ĵu��� iP�şkӶ�h�k`怼Q�Z�$��@/���S�m,�9�sEJ�.�w��&��	��٢j`��*�.���X�w�F���8�_��1�K�"X�$%�c,I���
�|c�����G&�[h�JS�PB����bbI�;01DY�f�=�w��n���_�����o\{��H�RG��h�]�=�^��Q�cJ�s��l����Dyy��u��y�В��eo�[F1r�4�Nk!�K���ߛ`��3����o'/r�Az��6�J�����sC[�<��/Y��ɽO+����M�i[�w��2�-��ԑuD�.lZ���p�ƅ���?����{Nc��8��y8ḅ��#�iЂ7�o��(ݭo�ܩ���S'�����uG5D�i�Y{�ށ�V��?�ގ��V�1TS���U�H��E>G,���%5y(P��cm�B����W����M�%Y�LH��j�
{ �d��5��� Θ�c��r�BX(ϲ5�9e��|��=T���v$�U�6�G��/�,������2"�R�P5ݶ��X��E��`�GzXa�����jEd��b<�����:{2���i�D�z�e�y��]3�+�joު3���ֺ�JL��C���# �jɥ����ЁTs\GI��b��h�J��d�+:)��P2X�Kt�2ȉ�B�n�=��BV��WG[�Ek����̘�D,C4�$���� 	&�6nm^���, �su�~�&�K��č�;�q��Ũ����|�`�r�_�^�"�f�xy��C-����������	[�F�����%V�ԧv����r̭�32����6|=�y[H��l@���B�#p 3r.������u���/�q��Jt�`��yn��^6���!�����n5�7[�}��ķ�h�0@�wu	�����z�K��|��CI�ƫ�?����(��C�������R���H=Q&h�Q�����n�f��\�0����-癱'P�%!���z,ԋ8jaH���6���Þ}+�t���1ƻ��9n�ֻ_��>�@�4����'9����~S+�9P��Ao�S�\/�,f��[���b�'"���S�_W@�j|���1�t���/� yl�(	�S�����q��J��$Ѽ�����x���G��R�" ��J����uaP��#Z�A�BR���D+M@-�^	a8��56�i!I{�+�霯FCd�*����22#��]���"�q�+dX�H"��Q^��Wz��ðQ1D'��=�2z�]Nj1��T��&B�N��"�x�3�ծu�E6�i��q��GU�ΐ���w�Ug<�o����u�u�'�*c���v� �G�2_^�~��7�L١���#1�χ���7/�w� Ṙ۲Ћ�-���P�.���n������X���H�t�����h�ź|���\�������
��u;[��'��|dRμc�7l��@��g?�?�Dv��W�656'�!�̡�Ȝ&#w��Kn���*�B[K��({kQ_���=I&:؊o5�8h�u����a\�<�_��C������=��zC���鯌s�T�2�����n��D���m��?ᮠ壾*C�1k��%H��=<Ըl[٤�GA����
~���� ��!ž�ɷ�
���=�ŀ���\��5���w�<��������9���[���N2�[jt)@�]�"����Ƹ�m�Y��^
M����Ow�F�B\�G�����0A�X�A�0܂<T�5��8���Ԭq\�d��;.^��vމtu1?4�;iId���OۥN�[��0O�g��\��&���O�[�g�·`E%U���e?ʣ$XJF?�5�k��I�-μ�W��h睂��ܱS���}^l}�?)en�uV��}��,|�p�˂}�ޔ��zF:ȭ�56P\g/�-����#��7qmc��bk �2���1�55�~t'��oc^!���a,��Sh]�������OH���<}Whs�����m \{����Y/O�z��A5�H	����F�q��Y��7�fnF�{�0��D9ᵚ�¶(]��S8�v׾afV����<*� �����M�r�*	8 
jU���(8�N������zާ�ޢ��??"~��?ɋ�D�L����v�A����.
����[0�k��"�ehgJ�W%i���HۙQ�������3t����� ��i�r`ع��ղѫڦ.���'�����lK�,؍:�Y�_�B�	�Q������A�@y~Z�&��C��9}=�4��_Wp*A�U��3C���o(���?�oX�	�b%�5i )��3�
	x���_.�Ә8ZVc��h���}y���U$z[�aF����@3��~���y�էq�Pr�佒Za����
����������*��*'^U�E��đEO�����sG?�;��yn��a[����vcZ����1hc�^b�D�]�ؑ��`HU\J\T9��%���U���\�8~ɠ��������(
-��KR$5�F-�:���tf~���_��g�a�ڡz�\�g�4GZ^�����q�ڂs��{wNΰ�w�v���@�@�n����CQ�R����k!�‬F" ��%܇t�0�?}j�g�\/�A.�'�#�J@9߻���1�� H����ǔ�*��> �a�[��)1Tpg��_��k�?(�R�0���e���ݲF#������k��]�WE��^�8xď�ϻ`�%P����f�����V_����5v˾�C_���s)5�f	2���E�ʂw�� p���r�3��L�_I*'�,_��YN���%��&=��G�iVJ���'��_��� �� ���dx�$y�
����!A�1q:!ԧe�a$A�Al�����4��o���$G�)��q� !I1���3��y]��K�~f
HÉ�c��|x1��l�0a�p�r;�F)Z7������ح�'���ί'�~�K�g�"s����M�p�����Ħ��7+~�n����C�k�ˠ����I�dL�����u_MЉ?SD:n�6n�|4�� �K=�d��w75��i݆��2�$�-���"Ĳ\.���]�Gd.��ft��x�6�V^����2Eկq2����ڙ�@1 a�m�A��S����+��([�.̣kP���i��Ւ�?,h㥉hyt�f��!v�75e����o-��s�VY��шt-"�8��$];qΌ7tFW��s��6�
[��z�}t?��ʝ���K�!�&j�����]t�E�W�H��?k��
{�oE:%nvB�U���j�p[�Q��5���ph���e!�>T�����DH����E���|��JE�}�],֔�\�������|�&���[��r��Z�2���i>����7�N�#��|�����mv�3$���9L��5�H�d�5-1~D6';Q��o���Œ��5��K��$�l<`���e�K�r��������4�ũ�:����rO�ؒ�k��d�03���8����rdq~E�8gu�t4�����*�z��C�ۼ�q��z�v��͠X�/�}��B�ނ#|�8#��RMɚ��I���"g�����*C�!��x��$�7�KO��c)QH��@����[4�+�VP����DHx��4�R��Y����{�������Ńa��*��������v���ۭ���Z�*�b�=
yP�Fy!�?��Δr�P���t�+�ja��H�^9+qVt�ل�g��@�=t:�ގlP������c�:��D��8�qa}6[�kw��Zn��>��w�}��V�S�"T�[�����2�0� �)L���r�f!�jSPD/K���㕲���L����5�q�Y�@�:�bU��5����6t�z�&t��$��Y�^�1�/Ep�k���'��u� ��3@F���̚t��jƴ30+sd?�xc �zѵ�9Pt\%(�e�˷��;ݔ\W_�ͭ�64K�b��ԉ��Vh40�iy���h/N����g7�(�S�����Ez_yq'5#��\*\��h��do�y�Ŷ��&�6n��=7�?¶t�T�0Q1������.cQ8��P�#&z(jC�0t����ƫ�i���&{�����M~�H)����R�j\�Q��S�i�?i�7����\jj���.K!O7��htr>��'[bn�� Bp�#�LK�Vd�NLƸR���[!��vzVbF�o���Yч�#'|�fBe�I(T�xxܖ-������3/ ���s��$��,�,)e���%{=�ky9��� P�n�,`���o���#�+|�>P��Pb�����>r����Cdp�M�ROÛ�"�4;<���.k���yE����Z��-4S$S�ɚj-�2Èk~���B�-s�%k���<O����}ǈ�h�|�B���pAn�JϏ������A���ON�r]~�}8�F�mz O�~�E��tb�j(� ��-���E0��컍�h��?��:�4U�4@�磂�Гz)&��J�G���j;�v�}��|�N:���g�Usm�������c�� 쒲
E�|��������{��2-n��|Ѱac�Tt�;}��so����9�c�ے�R����+�T1�-�!ɾ�$�u[1=�e�,�Q���͠�)UoއILʊUԧ�r�ǩ��ӗseP"tDUӐ�w2^MΫCmK�z�A�L���*w�9�������*0HCOݸ�#^�^˥av7r��L����������~ːԊ��爇w��[�`�a�4ltS��SBB�F���ώ����UT7�}�*���p댶�	��˝k���t(�4�%G���\xX�:E?�.�?�#36�כ6�����t��H�o�ێ�|{���R�?��j�ٔ����k*l����o�w��P�J��YɻU��i��O�������BS���%E"�P)��TuIx��n0sH�q���o6��C�� ���[Hvm��.XJ��"t�l'`��p������츲�����Hy�T���8=mGS �����g����E��J�1��˗�o��ʨ
H��X)iZR��7�hڄ:�؋����(sz}�:��7QL�({Hߵ��f�	�ԡ��5T��c�[�3+#���u�e3R^����^Z 2�`oճ��+_Fs=J{y�kDb��$���Tɢ1PhTr)����b�ت��ة�h}(fjN/l�&��?Y���bgO�ף�?U���P�����^��T�y\�\$�!��7��S<�exHNj�
��mø��Ө�D��Xia�FB�謈�$ɅW��nR�^r'Z�2��r_�\�7v���u{�ͯЎ.V��d�~�=/�3J]����(0�O��S�~���w�� n� |nzB+�,o_�ncN�a��,�*0�A��KN��h�'�c��\n�2`D5	�_��B�E����g�F�Tp��o�P������1� �ɣ��~[��OU<aNbf��.���=?�����6�	���F�uڈ���fs�VO�~��/���1/5:��^ukeEDվ���p�֡C�^ӣ�-?��uAu7�F�l�+�T07��,��;�(�hb�PP4/���M����`r�f �4���P�%��i�m��`���'ͪ�a�索�8"����4�����g�WU�A����-�2Ty;�ep�ڃ%�?[�r��)V�a�7!�TNb%����)��̘�/�Z��}���>�e��"U5�(��am�#��5�����ޢOqt���=�QU3�d��pi���C��Cƾ�׋�� ��$m���.�KD�������
Y{DE����H^�Bp��t�iz��2	`�-��:O(}�C�u���ް'�p!;��dU�BY)|��gg0R�yce1�g�T�g���xKaC�޺.�5I�-��0�K�?�T�܅�e�rmַ�`���{X�b�P`]ԭ��c+�w��hdE��%��6&���
��j�p2_�]�=��vr�s�q,uH1���j�h��̌@��)Uw,�w�{Lܼ��Lo}9̍9H���l�rI��d���K���И��ҳ'�'��ֿ��M-9⥱7<�'��ioNb �R��t��2?`�v�1C��/vt�B�Utݡ���2E�8�0^$˿!&�@�����L���48�ܰm1�Ͽ
񇶡�zˇ�\��B�>>���>��"�*���yZ�yE�ط��Q
�1UsH�% U��ʆM�Am1sľ��.�/׷����-"���>ܸ��*�9iR�?YsYa]�אꂶ:�aX��~^�m|�_D�B��/��y]���D�'O�����XI4ŀ�<d�7�k�fe�.�Tn�Ej��#���~O��#��4?-}'�f��y��	�<�i\Z�57����G��`��}��y~GT��u��x���0�/P��w�A&(�R��}����z���[������//��)+Ϫk1���`�������n%�2}E89�Oۢ���R��]5r�b̰��ʰ5�\����Dx#���C�=����;ԨCU�����
����4���ʄŎ��3Rk����Y�)���s5DH����?�i%�*�t�xY�
�*�>]�$L�pc'�[Z�/�~wB��"�D#�7A�[����1�>(+�u��p�4�V��Q<qrfu9�u�Q 	@nT;�S1�p[�]�~E��*8)J���St�V>���_�W��n�r�5���QI�+F���h�C�r,��Sh��@��0t�g\��,$AQe\��� ��n�5#Li2�:O�@Yl���4▃F�=��7C�	��aE�la�0�8��Տ�Mx�]�_�jTיZW����U��(�����jjj��.�(M���?	ߝG���̰q��XOa��v�q֮��P?��2�S��4�%2�ؠ�G�V
.����BX�$y����s�qK be/��xڎ��^IG4���4]��IL�6�PWf��f�w�fq��\e����d����R������x�D�ww�Mc0��oal*���m�y�O�짏��v�PI���R���q��"C�g����@�)ű)V6����j��r��
D�R��L`!W�`0^��^��#׷Xğ�խ��O�Xx��f��X��N�b���n%�ldXGS��a����:�!��*�K��:�Y.��2�$w������F�h�paNf���3���|�$I7m�C�<4�J�|��@ ƴ��ރM��}O}5Q7��:Uxݼ.&�_��\���4���Z�7v'6���+�����`Re}��렄�X�%niѺ1�͖�d�~#Y��������w����u�g�3t�ۑqd{��\ݷҤ^%DC�SjΪ��_4�D�K�ʾ�?U�g�{��6j:aB+6��
E2��Cd9��2.X>*�g\>@�/��;�r�!x�M��Pl��5/��c]/N�B佺hoR�of%0fԗBaJ����S��$�w�����S+�O��&�xp���ź�B~@��!�sy��z�6��3e�V��P�5Y����DGV����C�ŋ�M�;�j�d~N���E�7;�IA�͔�Q��u�x�43"8��_Wq����IK4�'�s�q	�\�奠��bL(��b���m��A��ņ����5�q3d�0�CA��O%��r�F	���-;h}Yc��<8m�7xR��4�_<�R5X��7��4\��	s8�P�|�{�6�'@_J�]e�adu|\��1h�*��q��vE\A&�TN�7t^��lYE���Nx��󸿖C�4��P��!�ˇ(X��(IbI�(�XhO�:%������p�5L��r��!�$��C�ţ�U�����[����S�xh��5�ef�s�a}�}p����S~##ǆ�Nʲsv��(#�`i*�e�J&���uyn�ȇH�*��� ��d2��_�hM���������Z<v.����^r�zY���q����f�v��~$�UqF P�q�.����>�\������/µ���k�'�3�,��M�b�J�G|��?����4�<Q��=�U��K]6�tϬ�G:�z�����"�>W���&�_����xnN��C��ւ��)Jθz9v*��t�]>�E'j�~i*#����q3fS� !�Sy^�����W���Z�˥���&��1@��8�����_r���]����p�Q�oST�'}����d���?u�����oxA�*@f<�%	�I|w%�\=����B�ﳙ�8e�$z���oh�<'�"��A�ie���v<�@3$׆��]���J����"��'�A/��,?~^�Rh���l�i���T� �>��,�3���K�h�J��\h�bA-Bک3��L�E�ǽ��i��r_�q:���떵�(x"��.�QT����(p���FV���B�����;;U��.��U�`�*�����	�0��˴V��q��p�<+F�4��;��ag�'ET͌�#'��UN���<�-�@/��yj�u�i8ܞ�����Q�`ݔ��s�^��jÍ��u�6_[E	0dǹd�N9?΢�������|��W��?C�:ðnϏ�fw�آ��%_E|�:�l.)�O��a��N�"��Қ.o�1�@̲86rW�����P���i�L���Ly�-�q7�m��=2��W��m�`����(���a�\�#�<`JW�dJb�AI���R��������%��C"Q�>ӚH}c�niC�E���91��sA]�����ƥyO9^5��X�*"{Z�L˿�섽\L��m��X�f�a4�x���� r;���q_�������ٛ����Uo ���o���zy���Rd�hM�2.�����#K���HI0^����Y������0
�c�n:��T�����¾j��
����u��/�8�G���0�J>'��u��r?�hZp{<N������bP��v ����������g���+�^簀LF}��r�`� So������B�	Z���[ךۘ����%���<ӎ�e��	wmw+�]*�K�-�����*�*�^�,+߫�����:z�<_/Z� ��CM;6b�O�S��*���Uv�s�<��B��Ý^z�S|pB���7q���{S4�췪���g����s]B~S�>c�V������4�W6j�׫�j���G���
pγ��y��oC����P��t�',GE�<���&]��.���٩K\���l,�/�r�o�b�\{�:�]]p��V@�tU������������kL'°�N^��8 ���H�5p��n�h���r��&�j?C;���`��Q>�p�r��X��{�'oBb<�W4��Gc�#����$����C����z���*�)��Ej���j����O��:*����8 ���\��5�x��&�|E����[��E��AA�����L���d�}ޞ��2j��_%���R����;O��<��{��Cb�>.�����̷���!�T��8�����Q�O�g�H�@�`���o��*��W]'9z����\�R��� ��eȐ]�,��sۇ�(�n���޲X[����Zԟ�q"LyA3�:��&�U30���Y;�S�Գ�B�7l+�6(H��US��e�NM�e}�F��s]�'K���|��{tI�h,N���Xe�^	ۈ=FSt�4B��fJBb�LC}
�M�5g�x���|,C,��L[�|�)`7������*��� ���ǈn�&>����n]G��#��@�*�g$w�ְ��S�|�X��'"�ue��sZ[�����qx˒�Ů�'���k�L�B�����2��T��\�tӾ��"�5Xw�D͸ �)8��#��љ�&/H/�y��&T9��>����5���;6Κ�+��݁G�,�-�܇h!$�����+(X#Q�1\#®��?�1�?�M���07��mS���՘=�^��Q��e���Z��S�D�`������\�2Ҽ:�5�'���2���n�j��H?�B�t|?{������"�"��4�%�8H���k`%u��j�]2��Ϋ��aW�r��l����w���	�W�2x��=��V��]X�aB?رZ����޿�ğ�ym-bD�`�Q4��Z�'���g�{�j�U6���K�i@���	��\�;����X3J4�x�p=�D��a��'	=铉Z�&;�W�nxk�"e��5� !T���3��𕁜Vi&/)ɳ�b������~�K7�zBv[K5,�z-e�gV��5n�?��DQ%�Z�I�L�l8��5����%h��z���|���oJ��2�v;�o�$W�[Ux�!�O�|u��~������ˡ	�nO������5��r�#��Wy�#;t3��V��$s�`�',�Y�*��έZMǉ5)��Q�şT��@|��_���
�� % ��B�N�n;��M\�ڹq��z��t�I���\�U|�72����ee%3˼be*D�Nm��kf6��	c�:!v��C��
�x똟D����?�����6���k�Y�K`�S~�N�gu��M� �p93z���y� {�"E�vʲAs�P�]D�߿VG�kF
WJ��2��a������m�Yϴ���Za������
0���Mk�p|�軯�:+�R2�M�~&�i�f��$M[� �������oԓiZ�ٌpN`2�ޭ#a!��8�M G��Y���*��9Di����o�\��K4=¢�x-B?�7ڵ�n�H�+ܫJ�F �{Dg,=��)��??�'=fI�˸�a|��ɻ��Yq����"���l�37^��ԁ�QL���m�[��f��gz��������ˡH<~"4(v���y_,���|�&y�U�Eh3�+�/�HީUF���b�A����F���O�*�3�-.�g�X|?�f�e��u��j����<>�p��h�\�fE�����4Cr��2��X���ϓ�������[��
jzC�<���#F.�v�}�*,�'h�5�mg���%�GV�W�1���X"q��:*�ܣ�ԓx���G�D��Y��{�<��c���
�?�2�<jK�TW�T6`0�K�P�`3�3ȶ�J�t|��`g���#�=�k7�D㫛�F��p!92��z��=�卟H֓s:�@ᛶ0h6VZR?����eY��E�b��1�'q��ID��}�]��������h��K�L^����'����㱶Xc����K���'j�\>k	�N¶H���=��W��^�$#��ޱ���"c�H�pL�<���P��\���%�D��d�=i��ܕ7�|�Խ���~�;����]M%\I����"6.y'y|Q���#Bhu��xZg� �҆(�8B�u.L���1;�s�f�-��2ȹFaw|aÉ���?u[Zr�)�'"�+0����^Aa��31?�7���c�ꍫ4��{����&�@��ڍFDk�`y��qn�.k�K��'��+ӗ��\M�ھ�w��K����<AG8�s���%�R�0&(*O�+�[�]!ڠ縣ݩ�scR�n]�A�g!='㸄�#��X��ʞ�e?�_�2C��:���ǅ�
��
�/I+Y�S�̭Qԣ�20�OX�1hY�j�`[�����7�o|U�߄�l�v@��r]�Jh=��GF4!z���|F���mx��nV�O�p�#u�!�$K���F�Q�a%#5�Ϥ��K�ȍI������)&��E�B1S��!ĳt���t#pկ��2v��aĠ�WD�w2����JI}�r��9��7=H������F�=� j��/:H�� lNM
�9�W&�����ۛ=��9��C0~�,�z�@
/��xa$	�� �|��Oh�ʖ1u�=��yk��g��P ��@��Ұ���w>M����Y��Y�M�6P��D����'(8��?�Ð%F�+f;bo/��Z����}����'uB*1�Vo�����
�|/ml���7��uE$�"S[�ȁ��r����������ً��2�f$y��T�9�;!�49E���%��p����)���x|�A
�Ϡ{���7����xw`�dv�wƏ"��"�$�@hA^@J�p��q�ܬ:Z�ъ�7��H�c�}M5uԇ�PǢWdە%�\V
[p���Hbw����剤^���.~	}c�&*�WD�
����_'��eޜ|7@��	�����+�[)^���U���K��*/X��@�f�*�gk\iYP����/�պ�k�d���^���?�~��B���R	~|6n������
�q����l8���X�*�(ز0+
���|�]o[��u�\Q�d�LM�^bƿ8� �8�����tȵ�LM=�{+Kt����=�bE�'��<:0�������K��w��ɂ �e:/���lU���3a�Y�/����׆ �qx
|��2�մ��	A
����V��q�&�Y-�Pj�Mn��l�/튶!�s`08)��m���ݏ��=�U�;�ٕ�S�O��Nm�0�XX$k+.J3�YM�١�L�+E4h҇��nm�V3}r�7�z�Ix�j��B��<�n.��d3t�#�:Ǵ
�Z�{���N�Կ�_�ZIF{��K��_	���
>�G�Q�𯇾T��-�E���� i٫d�!���O`cK�F��\���e�������ev�F�ݸf����Ĳ)x:����*I^�z���zo9�i8*�����`wS{���e�$UVu�n�/��c�^$%s���}�jۈ?� !��y5U��|�0�4�c�[��Z�q�H��	�{)c�#��ߠ�f�}p���@�/�E��Eml6�O�@W��(t��CP��x���(�a7���V�}0�_��K�ٍD!���A�����@��z���-6N�狣g��+\2�7�	?Dϑ�*�wvQzSvdV���I���u_[�DѧU�kT��S�!u�Y�K�����V]AMѤ��m��L��`ߧ��H��$����u�0�U�u�tb��9���ca��>^i�:��W���4ÂR�덀q�v�\���̬x'�!��E��I?�b���C������A�\DJ.��xj�=jߤ��d���d��I�f���C>��YI
]�b�լ���cg�3^��W3j�V�s�� _�PC��,f:�v��6��3����P�\�Q\+�<cE��Z���]�x���/T�;~@�cT�΄�d:i�QEDDao/��r�%� � �7�뉥�8��1��P��ӎ�S�[�:mI9�c�&�����mP�#�:m��\�Tz�(C���p�+kͣ�0>����G�(y��/� ��rm��$ǥrou�<��n���]�z��n��j�������]N(�Up�#�{v{�����v��ph��a3wh¯\m%����:8ܻW>=q��K4�Q]6�&:�&�J>a�C�<�$	�	d��0l��:#�K}���o���F=S���t�6�J�C��=���%�uV�b�J31���s��1��q���I3��p��G*�:�:Q�"\wb��p��{��Lg ���R�$?���k34���k�j�?�1o��TC�%�y���l�c�d33��M��z$�{�r#	��@.��[�G u4����S�@�+�{�вI pP3%� 	�7~NOѐ����]�Us�"�܊7.4QH'��\0P^_;�< �|�s�'����噙�&�	
�oF�+�*t5RW��H��r0CouXF��Z�&�	�]�m�IP0�K����2|�[g8T`suf�.Z|�(��}`*�J�ס����ힳ%\���%R�j�����̩�%b�P��4�{�-Is�W6��M��PIV��Um��x^ZRR�����H�
C��*t����Z�(8P��We=W1�JM�<���] Y�@�/��@rN��]dL���[ڸŉ��X�a����o�[�!mW9l-���Z��D���/�[=���'�X�Ag��G�h��n�"*������C�4;l�t��5�}�+6݉a~�W��R��ߝn$����΁h���3*��]��d�{��v� �U�t�3�hNA

��k�n� �����������������^�wR"�ta��QO���ه�eW��H�A��TP9}z��a�[1A_�`P�o�*�$fj瀮��,1�x����9��p�F�1c�lU�@B;+Z�/�	���+a7��e�4�>�g_�᛹%4��c��{�������j�FE����e�h��'��YP5���a,�J�(^�J7�}�~������G���V&�(��f��c57Z~[�I�Oc6�Q΄>9�sY=�9D���#��b���+A���v 7�K��?�}�5��L�D`X�~�w��x~OS�ղ����z��>V1���x�ź�I�ې0؏�P��%w��� `�Zk4��Hrh�A/r��4D�%E$u���6Apb�dl�u�؈yR�xf�y�U�,�Y��E��$�d6?,=b��3K4a ��MK6걢eUY�_a��5� �-@-�R^�>��:fX\�,b˔����/�Q�S�/�]�!7�.E�3�c�Lt��LNܖ�^�[�n֦�ߧ-��Qari)rG�a*��]�.,	����&���f���E�<I^����'�P|���|U����de~|�!
�IR�0�%(U