module ncotodac ( clk, encA, encB, en, mode, sclk, sdata );

endmodule
