��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�i��a
Α1S%� �uj?�L�3��TLei-3^5]E�$��`+����pU�Ei��fj
,*����F��mX���� d���*�[p����=��Ϧ$��y�R��@n������G��_O!a�Yz).}�ʊ��b3���t���FxÖ���o���|*	���b�PQ��ꝳH����X���,ш����H�YT�d��#�~,CAt-�Ż���f4�+�P��*�LH{[ُ1�X�u�<�xZ��o.��h�ʟj�a��mJ䀘�|��} ��Ԭb���עTN���W�W�������AhD���@"�S�J3��I"q%?`��g5�= �M���*f]`ZV��d����H�
n9e;i8��'�eA�4�gw�WP�����i�ټB��A8��!�KHHf 1HX1*�ci��#>�6�;G���G�l�¯�R�����Y��[���X���q�����!;�Y���������/$��M�8t����&�B�K�x�C��8�(YB��癬���:뫄~�L��+g��o	IN� �f�D\�?�$�6�uU���;o�[��،Q'�sI�&�.���fM�Y�j��;"�5����s6�xq�e�'z[��ɘ=�����qu�1���[lS� ���C ���#� �H«C��c�p[���� ��M�U3"�u��FL�g�QN�F8�����G�����Ƕ��J{���7�OƟ��P��re��eKv����ܪc'�C�"���򒾞��tWC�Y����B�'�ڪ��8�_S�>�ӀTu_���Ff[���w}�-,��)�a��Xd�r��Ӈ,�����R�]�_�+ V��[�@�!�-V��*�͎�=q|�X@��2��+�S�9E�|o��9��	���j���]v���fguz�P�.�;8�q�ŝv���bK��%���X�^��%ɚ�Ѝ��|_]��w]�M]��Jl5�(��ɺI2��[�[Ɵb�?�L�0��y�΄@R�dg����K����s(�Z��w�v�QN X���2�<��b��!��m�5}�B��F��/Q�(����HƮhn�7��!D/_�nKA�K��A�FZ������M��+�of=~)�It�N�UN�2��m|W�q����"��843/֡�(���l�FkO��du^��r(?��o9�㠃�9��ɀ�?�7�l�@�>B�;�-Q�Nʷ:�(�{+��@?��z���ϙ��Hz{��R�6��T��T:�?�n<�Z-��Ԕpf�k�������JBێv�oT �-ܑ��=������$��|��;�t�\� ��V���执�}��U�P�lBy�����|���V���H�Yˈ'��LW�� [W!-@+�x$k�_&��@�5\��!�Y)2+�1�����~�MJ�76wb��ʣXYP�A�R����Z��_0�WU�2���;+��[s�����:a *e��O�*����eD%tR٢	�wt\�1,T}!��[P��N50���X� ,\�2���6�.g�.��-K�H��'o�_lC������J5�z.�������޳�=����~�w��	I=����vc�D��V��a�����ٮby�+å'���LR�4 �/��z�S��'nB�x\iU�u�ǖ�G����$=>1��y�8��{�����h���C|Ni�2֭��n�z�k��%�Oژi���Ȱ�]�s�pܝ%1m�D!2�_�Բ� ��y�2���`�8F^�r>k�]�w�a�0ia��U���	̻��ޔ��պ"����b��G<�*v�P�pX�vBnl�&󤌙d=�@er�e����<� r��S9�G
Ɇh<דӐ�|��fSh��1�JJ|'D\�4�V�l���aᄇt��L���gt�c@�F�~Wv�.�q��g�x�Q=(�T�ġ�ϩ@��~� �p{�^KA�݁W|g����Ճ����JX��
��ǒ������V�oW�l[W�G����� �Hr�LM_	�Ce��gwCYx�/`�@��Ю=9q�A�����uE��p=Զ��b�G�rT�(����Yڣ'rl�Q޸%�Ul�>+��M��<N��P�~���P��(�BF�ib��d�Q�?�E�u g�5�����!�~���0F�&S�R�"~�~di� ��W���I��
����[�fxa����Rsu�4-j%���5���%:L�e��c�
��U�N���	Se�����nԀ0*�x�7��Wԅ}�F#BeG�mS��]Q��s0����CƗ%D�?{0�3}����rh����)�������wzɲ`��ʛ��-EA�KI������>��'2�wV�:�\��j��ˬv�&Y�����b�SOA�����j�ی�N�i=�S0��4��sC���N���Ʀh>�`M�̴���������[��Ur*�|1��|�JX���?��(\O����o�/O�ւP	��o,1]�p�)����݄]��X|4N¿����E�cd����ӕU����|�}�h�#��H(ѦZ5,������g�;�r3�ykp"�����X����9��>[d��^rw)�- �k��{$$ n�>6��n	��7{�d��0����h��M�
�$;͔-���3`�V��� M����j�"��o+9�?ݔ��Y�ʂvC�A򴊚���k�I�D���ht%掇x�k��Ӧ�ZʸB���Rv���t&��nN�d����5\U�F�ٰ(	�2aS�������}��foѕ>�E��E�R1Q��S���/�U�!�=x�~e\�|[��]U-G݁��xm?���2v���F7lx>* $�ΌM���*M�e�WG�>L��9 NH�_@�]jE�S�����uȥ�0���[�}w���(�sW���>L�Mx��A�_����W�xAҠ
�kFyxI��,�E��J���7�b�\�h��~�Q���׶Zg�4���%�䉎?�=����@���m6�"u��jI��L����g����2,g��f��z3~���!%�)#4��!�\��e����:O�ZWOPEA>������]_��ο����S�p�Z��Y�y�X��I����;���v��������A�b�;	T;uL�qnf�_�YXv�w-��`%�CbF�!Ur��u���wK�����I"ʪ�<d��4?�y�ǩd��;"#@Ai?�m�͎b��*x �l��?�,��YL�P4bU�-�Ƙ�����i�Xs&�X�����IAI��K���zȍz�@��0P��˒��o�t6��ܘd�Q����f.{��L��d�2E���)�V�7c��u�eG�����(�j������v,e���BYֱU �v�ikj��(��j��
P��=�D�B��Ce��,�1& �}�� �ٴ/a����W�`Fop�>}W�����ф�t�{�P~��z��l�=��s�OV-Z��|� HU�|0�T�c{���x)Z����ҝo���_�7C+.���n�<�-�s�a��� �?�����#T,����0G;�L'װ�t,K��B~�Z��������TBL�7d�I���1��T>��P+��i��.ſ8j�P�%䥔 l�1����	�琨ė�ͮ�����(�zP�������;g��IT�S�����h�:�'�R�6�ua쯙߄B촁���{.|�5�'�n��B�F���yms��z�5C~��}���&,�<xm���5sX�<ܶ|Q��4VN��Q�T��.�u2^�#zQ�\�AS)�5o�������1�;R)��)��|�4QM[r~�Yik�pUJh@�5�oos��G��M�"e�yx�;_Q�ևh��u�8�PQ��<�(uj�my����Y���zJ��>�1
�������ˡ�~��iAF9V�o0V+Ԟ��i��e�qN&*�i�!Q�]�)qa:��9�0�A7����P
�LE�̦K6S=�T0�����o��8eF���ߚ�Ad�:��z�����Y4��;慘K,ӳ�r Ç���73'[m|�r	���8�A�]X����˪�q��')Qm7s�G݀l���Ų������|v���!�3�u0�W���y[�U�?1r�R�;�#l���x1�p�.-��b�Z$Sֶ߮��G4S��a�>��{#E@�0J}������ ���S?jM��6�)���HtC�X����9���l3��������J[�_w�F���ӺQ&�Kb�N69��H��
`����{y���K��QqY/$��1�(����͕X�|�Ӄ�W�j�ץ��o�ݛ���Ǡ�2HƄ�O�f޶�9���;�8�'�>#ںs�|���o{w�=dV���4 ��/W�j���FUY4��˦;����.�>Z��X��մ�q�S"W�\,�v~���.�����D��҉i:P���<��h�.]�6��M�i���1�?�� �-��fc��3�}���A-JE��7�(:���/ǥ���X��D��PW�e�u	�����=�����%F���R��jE췈�������!<��⤴姕|�,��fN&9t�Zò���j���S�cee��^D^T� `��2�u-�Q�����n�D�$�ݏG�����aX����衚$ ~�B�;��ˑ���)�P�\����r��h]�F��䙬݊�6��t��~%�L�� ���x��gKH+8Q�D���B�t����3���"�)a�{Ox����i(G�Y�]c����{!�	�?{����n�%�'0m���%)�B~g2{��B<ZpF�tA{W�^!) dJq�^�L�h!���|L�Ub�o�v��%݆�Xf��5��S�:�0A�S�%x�wA�G�S+�8@��GMm\9���ѓ=@m@�(5Fd�HP��k��o�ƹ��mn�d����ș:?�?ٔ��FUI�34Ləg�뮄x����4c�?z��"ԝ�=ܝW�3���T�A �7��r�48�YB�Ʉؿ�rѬ�~�{�A���>�)���	
�zKM������<�+�L!Z؜��u�$q%�Q�k��9��
���\�gْX�IzH(�[��3�����e#^����������֘k_��Ja/��R��A����������ڳ�;b�G�}�KyΟ��*e��IJ�_�*��;;y�����MV��@-��g��qqӅ������5�FdR�B���E?�{�j�.�@�&U��_�Ѕų�q_Cgag���1�c����	��e�sx/�)G��T���눅2�t�»���Gtp�ɜO�c/���C_|WTN��&�P�Ǖ*��N�<�e��<j�
��@S���gQH�7�^���J��K�k�zP!L0k������µ*�fQ�-��NF�qv�d��]��R9�a��� ݟ 1!�������w���RWrə����I��rfx���\���TŒ�VM��&���M�%)b!������pS�,�N�m��?v�ඤ@��8i����A��ѥ�$�B�;_�#.����D�̺�����b��� ��� ��YP
p�i/�P%d,�>u���x�����4���G�dx���#�'��[!��*W�8!93u���:�3DT:ӡ��m�D�uj����6���z�F�xT_\��A^�Y��Ï���,g��K�t��ڍyA=��������=��*��	����Z	�'4���>�����d�:�\�þ4{A�Ջ�1��r9��Vg��Z�U8*Y�װ`��>jSp�k�2P������b/Us(	В��E�hh�շȘk��`>MJ3����|XV�@�|q��
�>��vS�N�6ts�LWJ ��tsx�c������j1��=�v$�ݢ�S�	�'�) -l"#q�\������@�8�I��3}�w���4.G˲���4��B:kW���z,�&�}�o>���� 4�sR�*���7.
���K~ �[�3�7�Zil�W$���>pG�`:v�1���U<$$1?��37Ґl��Tq> Q�% ���;��1��N�{=E���*0P�U�6��Y@�=��wY����z�:pZ�=A�%**'��5CR[����P[����跄��$c�g�6�h2�� W{0?p���/l�N�"��A�2���,���/$�HLGwi;M&�S�Q�����8�%ƒ�U��	�&�4��ǎNNgE�|<|���Հ<i�P�t� �a#�O9r�.u>����k�(!��>c�_��js3>0u �;�A�x{�m�T�?�]�M�=L{�f�<�(�g-�C���=��f?>�!}�B�� u\O̕�	w�]5�6�jL��4�0�v���U�5��0��ʐԙ�ڭ�㨅l����|T��!�������?�Ue����pt)�~C�̚�]�\��Ҙ3ca5h�K���q�?�Z%�c�3��Vsr�#w�~�F{wh
   �?+�`
b�@s�g��%Er8�
��KJIGn�	�Y9�U쟅`Z˭���ŅVc�a�we��#~��n�Ő5-���c k�$*5I�!N�3�/����?.�?P�?�5�fc�q��Y����`����z�h5�z.j���g^�H|m�����j�6���Z`V�{y��T-[�`�*�SC&Ye�
Rź^t^���8���>�������
։���w�K�}��@$ &lv�⬜�<�����骇o�Y�ڛ}9�@�S�$�G�)*��c���v���OLt��[ �ߣM[�̛�>6�t
S�CE?iRRI�n�B����0��,�BI��(s�
�P����}�,n���`����*�J~�Ld�a~�>�x�u����S�X�T6�*���6�"A!|�_�y�����o�6�!d�Q�I~`�o�Yt��.��_�J�'.���b7.�|��1z]�g���F���>���˃��^~�:���ԏ�&�T�}����o%�fF4�e����4$�=5��J�2MfU�����):���\z��<Y��KLj��+��N�kNl6!��}ªZ��OcEP��^��p*=��\�qg�%fqs��$�  6õAI(�}�P�Ͻk�픖j�<
�.�3u����y�%�뮍c��
�40O���؁�ُQO�欯�E��M1�v#4�ȹ<3iv����`_�e>�)lΡ@a㴒\RNlQ0�s�DMG=����֯@�a�~��w�� �H�� ���&)���U �p�dhW�au(��8�0#��$�{�k�7�/������0d�L4��4��6F0ɜD�Lz�v��
���/��E�;�� �Q:�x�W'qxW�I_�fF�T;��E�;�}_ڣ��C~HY�Mө�B�\?C���}z=��J;N��	��)�s�A����}��CVmC�#iK��1�g�ǹF�>k��>#&#���FQQ[�j���|����4g����~�ݘȥ��Z�k2�(���q{ڝ�5C�_R�S��?O�yH�[���̺s��7��e�ܯz9����YQO9��(�IkKP�.<�[8�>��6I�v|��z��q��C���������U�)ߐ��䆿U��i�I{D��z�S~z�s��9P����UF7��[��Z�3�l�=��o�&�.w秶�u;{��$�	+�ۧ��&��F�b�]ɗ���O�{ ��Q��!�Tô���}�ߠ�dL4�Q��q���98c%x֍�C��p�$�4���B�;,~X�.����"%���P�1y�BXR�>�4�"�^�Q��
`	�i��_�R��.|��G([��#l���k��ƫ��U"� ׿Yă^�B��{�
/�{y��B6	�e�s�gR�pQ�e:}f�ӻh�-��l�\��V�����X�O��n�g>�wJ�˄�
3��5��M-$��xn�6N�����{���U#�N5d��|������2�����x�4�8�`���R�-���4:'`rc8g����C�Qi��ݗcY��HE(�+FޒK쑴�<Y�VU=h^J񂹀.�欄T���97�s^H���e�Y��/l	��w3�p�u�{GKt��\�&���:��0��7~���6�aS&/$�#�=�3>���H��+g.��B�V�ך�H,Nc�n������6�'�o�;P�@�g��"�bz=�ۊɕ\9Ҿ�-��5<}�'�$|��n�!�ǹ;o/�^}����[�|�?��B�cr�=U\����!�f��i�pU	T^V�Z�	Ն�b&�e�����"v9��J�}�5�U�2�^G/��t���k�1��3s�d�o)2�JS�ce���{�ȠZ���y�(��k �۟	΁��J�KY|;�KY�S�;��T�OV�'��}�䊽����6���k� �@?ޖ��0�Od��E�%�? Y��y�I1��������{',߅b�۰EWxX�"L02�-�D���QJB!�4��h].A�ECr�N��!_�1>��
�;8p\Nd�H��V��/<�qUWA�f3����_Y�{��b�g9��`��g�*j�§\�
�
�}��ntYK��x�w<��~kw�O������m�ot��CgN�����3e����l=`]�	׆tj�F�ۢ�X�IW�ퟋ������Q:�o���~�S����w�o��BTU.�uj~F��8�N�*���5�_���>����Y<�'m��M�;��F�],��,�*����8�B��VH /)���(�x��[�mj��2a��Ep��񂔹���2�ƾ�M����!l;��XU�����%_����;���{�c!z�Y�f4p���:H֪���ܱm��+�����[ژ�5�*��_����/��8VM��:A�uKg?2>���"p��1�+w+��/j�V�pH�Y��]��H��"�F��_�B�6۵��U���+�~���6�2 Ё('���67 u���\��]���􍸮FD�L�=6rZ�$-�݇�G��<�H�_@�-B'I%���Q�J���37� k@��!�PR/�$`�7���VJ�i����C���/"?�`[n�W(�*v	�aO�L!"J��,����+S�쿬�(�H�j�K.���-��-I��<\��=�*�q�]�+4��g@?.�.{�@�06�C���@�Բ?�
���jGhF巗Kvոݛ%�}$��&)��gѓCTv7��� ��q��\�ʽU����4���Z1Ǵ7�}�Q7�Rw��������Lֺ��)>�W��?�gb�Ջ<����~,�2��Ț��"_���5�c�*w%	*���E�{2��W�y�NG��F|6Iov�`�!��e"Z4]NUg�3 �X����Ef�A/��p�;϶E�|d2%y*A��~��ͥ�~a�ĮaB�	6�[9��a�6��]�`�i��3�%Onw+�å��ǔ�oK��3�6��_Id9Y?'�k���?��J�9����(2v�x��"ƪ<��&c\�����,.���Z�:���)XW)j��7��(3�� �ۭ�P|v�0�lY��0�Z�_n�о!�F��㫎㻅G�I0���A�a���_�0�Hi`;����>��%`(��ne���Q���x@�Q�It��e�z/�c=�3i����E�>��֭	L��p�μ#��޴{���d%�%һֆЋ�ҫ&@<c�
	Y.�ȁ�y���o��+|ME\ �S��Te�S���5#/r�c''���ݴz�����*��z$t�l�`n"�.�l��~@�L��{rۡ�a��Q7���9?&8�iv�=��H��dw5
�Q��wo���މ�癭P��g+A2���J�o�� a��ac���íWC�O3IN��6�<qHH[d��
Q�.���Z��(����{m� -�Ӓ�8H��m�1�s/��0hfQ��e@����f���	�WN�;�PIf���{u�L8�n�;1�O!qO�����%��#��\ac �aGpg��^�$Ô�7*K������2G0�2lJZ=wɩX��|�a�-X1��ʘ,��&�2�j�`���j�۠A����$AκF-���1�M�i����3��"�4}�\�*^��&�B>4����VPo
�C����<��8n�rӦ��s����}6b&i�
H0皛.���
[�qTT�w�Vϭ�xv��4�
�����Yw��_j_����[Ib��;j�߭w7/�/�%$�:��|��1��x���P7���R�Clu��&D�?�����uvjM�CQ�����~�NZ�'g8��ry�fXR�a��R0ij�d&E��:�I��p�O�-,t'
��C��%����a؎� �l��$�
�v
ZE��TAj�@��x�&�Nq���V0q̂SH�喼��s���e����J���H��曵KxBف�h<�|�����?� Պ��MhA���iF�B��|t>{k?�\O����d���ǧqgy�i�E��S2*OK��z�����@	���CM�a5I�|T%rj/�el&��q��УPu�c��9���ӱڕ���n|�k@!A=Ҫ�L��M��T�ӿ��t�Q.��{�����y�aR典��ƷW��oc%n�@���rߝ%K��I��C�1=�0|*\
B9��7{O1a]/�-6�E�w�N!m����b����������,�<#�gܣeڹ�r�4 [?�V�s�Lro#�X+��=���V'"�t|^ �B ���K�7)V%�	�]������\<lL6��'��Pp.�:Z���w��6]_�NNh@_O�ȘDVJ�ļ�/A���Z��7���K�o�������z��޽MƬ���%�#:/��!u�b5��x��mֆz�Ș��R�$�;�q�O����z��bJ�����Ϗ��Z��AC޽�&�&�0�g����L�N���?���&��=�t0V����8�%71�㯺B���� U��]'�����5�#���H��L��6����p�t��tT�Xb�t�box"F�;/ ~�S�q��e���'~I�μ*�pnX=�Z�>l��n�%��^q��1�O޵����&����g�ݞR��;	�5u�%����A��T�'��{��G�X���o]ͥB�B܉0"�=��w_�4�An��������m}��~�M�����}������q�/.Ǉ�7,�B-�q0�Y��@!�����1y��Rv����M0�U�����#h��h
B����k�jm��:SXo�	���=Q��4*���w9fxk ٷx(�{Q&�z��!e�������H[4	�������Ǳ����A�`���7��T#�m��̉� �~?/Mi��>��o��h#I���MֆB
��8��N(�a��Q<����G�8m����gQL�g�VL&��uzB=��X������lQ�ykH�
�v�N(yr��/	U/)�H��w6�=��V�a�]?���Roν���cf�9�0?�ؼ��S�8�:��p	��>7l��nSԀ<E�Oe1S"��c�-ӟ(��c^ɐ��C�$�vS[_y�&�mB9a
c��[mQ|C�J�,�5_��M
���v[e;I*�7m�1F8JzZ/��ȇ
y����v%�"�.�v�n>h��ϕ楲U؃��g��FK���^��g�]�&׌ �k�	m�/�?�
L��i�=���ݭ�-<Y���|�H2��oCI�(��ܵs�ls�RS�ĕ`B\�3D	��A��g�ĵ~�T�z8&s��؇�w?;%��>�ugqݍŐ<Ϸ�j;�|jBZ�1��E#g���������L%M5����qd�)%!}gŜ�d�o�^��?�ˌ���i�C�W����?�;���V!��]�5Fo*}Aωva޺�8�ɂ����� Nb���+�;��~Ͻa30dU�{�īE2��u~i>�zjv�'����u�j��u��`P"q��DH�6���M<-{TXM�n@ˋ�0t��\�9���z\�*��A��L1�"+Ր�F��B�?m�o	��oD���R�*n(k0X+O(���Hɪշ�+�S1�ib.��� �֐dZ�*�$q��u���G˴n��ܣ�\%��k@�Sq�`��F;B���f�7����e/�:k&/Ӄ�$4�`>*a��GuW��3K�gw��7�co.�/��Ԏ����u׃"V��_���P�b^��(��\��8��o(�����Jo�K;A�}WZ�N�Ul������\U``����I���\��Ϭ�I���^��f������b�=꥿���t��s��l("#CeX{�8p6��A��S�8`�&!*� J'��p ����r��7}+��bp��$��)�*9U`vͼ���g�����r��+iva��z���rgu�q�1�
��ȧ�%z�*��TL��)�S򽇝����>�4�ñN�nۇ�V�9��G����������J�ؾC�l�{(�0[jd��%�ڐ��ٳ���d�����R+���%���h�d �F�x��c�Ͳ�ӧ/�e��r7�@o1�����s��t�H	|&�8c�Cj��)A�=�������������fD傸��<��S�e>t�4�� �"[����Di
^7%X��v�M-73��x�<�����M@.�5�/x̍v)��QYGf����oY?��%+��qx� ʖD�yV�|=!�����zX��S������H�[Ǹ|�+�D�Յ)���%�E�pZ��[��yC�u��i��֍z��բs�^���~cT/_�ԯ7M�ϼ�+!���<�����N��N�#�nAO�ȡ