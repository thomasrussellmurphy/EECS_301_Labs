��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\���V�fnvx��ÍG_;�ȅe�~�>���9�>��Y;�0G���>��N�)��j� �v�{Mtp��aq�q�և���k�S�x�l� �yB�)���{����z߯�2o2�eq�ʛ��'W�v�J?˚D<ǱM�=�pr�˚�ОK��lqi�uŲ�AFF��9|"j����D#ě$�6!��깄�%37�΁�ĺ?�	�pX�F�92E���q��֓<�K Ku�pD��;����DUnŉ" �k���p�v�0T�a��c�:� *PG�|a�?<i��u��6%[d�����~��.w6����uG��Q)*�M_C"�r�7�6d�������ͨ�U�7�1`h�Sy�{Q5}i�B��������<?��}����?ֹؚ/��
�b(8W�����P/>��J��B��K�Ño���j�w|It������C��,���	+"�P\��j��rz9�8,92�C�A�H������ ���Ot�(���V^7��8@[ԛ�_ݘ��]�ڨJ�ꇠ���	��o�.f��q�łL�s)��[e�ͥ������w��3\���0����/S�n�`|T�E�]2/oy��`���(���k��/4) S����9�G)���=yہ<��I���>;�>�������}����8M�m]�{'*;��nO"�"w�/|�QQ���P�Ag�q��O���p�P>�#4��j��N��e���2G��K�.����S����}S�{���o�����y��`k����_P�&�r^^I2��%<LM?���G��o/�~�x�J(��c���G��^��E�P� $c��m�l�Q�k�#�~���b��_�~A{S���B|���e�3�4�R��'�J�Oqa��`�Q��Z��K+"\���=�F5(C���[���������/��"Ok�#�q/���,}�6�nCH"����Q��n�$�wޑ�4��]�@����mRF>�?��Rv6^���t0$>�y���q��V��H���a���g����q%pr�da�3��~ש�]S*��2�r�8�e��
�gA��9Ā��jF%�#��C.@ۤN���aou���V]��`P��Z��
�"�+�? 7[�'O�P�g�?=|�3U��<R����pJ�ey���ԇ=/�Fus:h~yV��G4��W��΍��]4X�V-�+	7+� �gD���k7P#ЛӠd_�'�Z�>�lr�i��6]T��́��f ���r�Ӌ�{��<_)S���C�O�%�e���1�LZ�>���G��ăM3�K��U�=�,� �P.cڋ��/�J,��v�߭�z��l��^���j�������/,��Gw�K�ya�Z�6y����18�c<3�Yi.1�f]g���'���g�RHx�e^h�%e����6A�.���)����v��n	�ܞ��,o�;�%8GĴ�]I��[�Q
l��~�����c��i�s|{/�d0�cl��x}���ywX��x�Α����L��ݠ�c�w[�e���Z�)`=�W%��Q"�H �Iy/M��o� O�	�fު"��<9��C7s��o��C(�g�G��Ӫ�	zG��٣��髦�Ls7G)�so�'.�}8o�d��V�g����v�T���TL
��/��(�bŕx9�X68c����@�46�̰�` �u�8쪨��/ܦ&i"�H1��{�2�]�@~��ට�i6�0��.6!�2Е�Nkk_Y��%��B�R΍Z��᯵Ք�2O�Y�s�U췛��g����$l�eK2v�VZGg�?0�V�!�],�=���NE��
�xo�My5��MV��b����s!Xi+�4�Fw���X�Ϯ_�������h00��~��%�:�����X����
����k�����������V;W>�/�e�ۀ�]�K75�d��H�f����h��L�,�؃Ֆ�ru�dv�<g�V]mՏ�rcӒ�hfs��yU��~B w��l{�A�6D
�%\Y�C i9E��e;S�2��WgZ��d�z �J�c{�j�i}%$'���eE�k�y��8]�'�{�à�����;7���Ǹ�j��V��&5��7FX���0e���/8To�1",�vK�$���GǠ&E�g��oZ����"p�?$����e��h�5�)+�O�c�xB��>�e�wd_����Ј���]�7&K�)h�wZ�k��9{�
B寧�����-�Ǩ���u�K�Gq9�k��S$OE�����p�?�j���yV�����a�VA$7�&QUuo�;+�T�6�N�
ۑ�5�!� ��L�6��V'�z޽*p���㚒fTv����v�LS}�͙|ӵ�8���	��Ƿ��؀.�e� �r2�v ����������%cK���t�qhba-ӕ ��	�Жp���ٷ���eJ���+���N�xkR�y�Z�F�F����)x����%��?�A��g������.�Tvq�9�y�M��u��40#���N���Pb��qC?S���M]��jHO�<�K|j�1=��탙1f���Cz��-�)_ò�Z�:���N3�g}��<�"�Zх���XI�K�/���P� y"g'+Y�RnX�k�V〧�jT�B�[��@=�$(�8Pt����Dx�e���-d_J
�<���cB�ξ���MH���z�x�Nč7{���D=}JQE۠�F{��"�p��x�K�(�U�o�-#��T��Ao>y�t��Yt^��t�?�t*���'�Ii������r����b�'t��|Dg���;�Ĉm������_{K� w�[�S ���x�4 \�Ɓ,�"��@[^����:�gP�)?�/�1a�����W��/�Ï:��gU�6`.����B.�FU#�5T.۴��6Y;ǽ���h��E#��h�d�e��3����s�vZ9�?���%��ã���H�m�Hm#�b'��rnF".q������+v���p��B��w:�Gs0@Q�"�0)�.)���Շ|�lg����K�d��$.$�d�L4q���ᾼĶ��"��g����Ф8|�ϔ�)�n�97��S�:MP@Cc39��o�ˣ�a��)�����ܜ/(��I�l�Q���6��)�-*���[Ig*J[��ț#��(��@�N��pR�Glk��$ԜT�E���ӟ��Н���١k�C(J�w��ɶ�+��&��z���W����X!���}ᑜ�`���&�*/r\��K����;j
ʰ�eZ�����n�_{p+��Q�mM�P׶<lv]��%�A���>�P55�x�����D��ا�r��m�GF��ŋ�ڠQ���@u]WEF��MHt|`i�J�:��Y��ogn��1�k]`�Fud���"���X��b�yt'_���߸n���`�&���X�a�yנ�8�K̕���{���Whh�2V֠v{N�po��o�Z~gb�cEb������!�_�3�76T�Q��J�L�>�0��xͭS�!�Ђс�%�Ayi#��Ψ!*P�C�H�|-B�FC�m����kЎb�����:4�]��j����t���b�Uqn�w{րe��At|�r��8%GF���ލ6�����:U.�$<8��L����@MLx�1E���h7o�I�GT��r֕U��?���;���E���K�f��N��:�3A?E�����k�ivf��H� �,ņ�BE���3��0�_#0�7t�_���k���q/��
,�~dcg!�F�Py���Sa��"�P����m�R�*!H4h�Uv+��wW���q"�A���u�%�N66�wN[��!*g{��!|�Ђ��YZw1G�u�����(�>��T"�0D�dH�3	_/K�^d�F8C�K���"�)�I!�&�0���a�O�/c�a vÂ�Co�F8Y�����PI�x��r�j)#>�	�پ�uqց�w�݆�B���.�}��;09l�]��l[�d��`������G�ױ�E��b����4c��ټ�W�)�#dJ��*��&�+q"i��K�}"����ԟ_�;�<��"��'X��.w�7��^����<�.���q�y�8�t�z|F�B6���T����!�5���Af�/[}�5���ku�����ipť_���s�3�>���Wp#����y���8j^~Ɠ}��K�k�'��N�y�@�=���nf7�Ԯ��f%	��.�7��5 �K��]�����v��������	�����V?J�a�@,g�#��������Q��Oy�ُY���)2�o՜0��TF2����]��Z|7�Հ3�42�p' xȵ[$|	2x��l(zxW��A	Qp'� �I�1:��*������S�5\S3�,�
+�Џ�Xg�q���.8����o���^;�S�9������]SW-��"[lt =�Q�vvh��[X�x�S@����%j��n��h���2D^^���>[���č4�v����p&l���� #_�����k�rFck�G?���� Y�r�5}V�~ 
��:�v��߭���"+�\�!/�tTQ��_�������<+Y*��D�M�w�+^d�/��d������޹�?5��i�A�E/��b���D�_�r{�|���|9Cʭ*�æ�$13���y��O�*�)��%�@k���ϱH��/�a�>j )�dO�T��o�=�^����=cϜ.nH���G���Y�dl����\��]�������޴�[m���-B�R67t�T��DWK���K��:M�����׽�GT�=\��^5泔/d���S��k�	�!S�&�a:��`& A���$`�9�V,']
��}���v-��V�D�����C��b\.$�y�F�Auͷ��k�E����+f&>ҩD����wFC!�B�/pzMA6ǯ�~:��R�{�	����d����5񠉊��U>?���p>�v�7�YoY]��R�ո�z�=�3KթG4$5�����|�6�F%۞���D{ �\�:�hi?pM
	���
F�<}�r�ki00����m ���י��G�m������M�� 	�Y	�OO>˓�mi��|�j�1w�������R��=�K��ʵ�rdBo\K�aՏ݂�Bb�'C�ދ��e]���u�p3�K����sW�1����)�x�,M ���0�G����E��S�"n����J�ҵrֶ���X�� �{Cz�R)̾�p�uD\�IЎ�FWN��ӕ:�KK!���~���+U���ř���@\,1;�eO��D�I�<�e{�sڨ��l��K��f�xh�`�ey�A�m<�B�Eʘ���~5�0{;Lr�K2���j��
�X�s�SC"$�),�� ���UEL�
�]��-���,U	�Ce�:ɛ��n�e����˦
�Î��:v���=�=ީ@���7��g������&G��sJ���^����;s
�m[x�GUc7�*���F�g���J��eU���aNC8T�7<m-��'�B�qh�t�q����r�F�������;G`�~��:������;�G��F�2�e�Y�O�����goB.�\�Y*�y1]����s� o%Y�ݍ�� �inC�A9@Ԋ�v�z������GM%�,4��Ӕ'�
Ƀ�Q}r�4��\���.n��挸>7��f�1_�A��� n ��%�Nl��{�܍� �{��d�8y�0W}�(?���o�5��5�xd�(��ƞ�� Wכ)g�j�yh{��A�>X���jѨ#��	�n�4���	MS�31L�Ux F$`���|+��N�kzAO�m�_������]�}V��(�~�vR��A��2�!|K�>���_3�^| �Mӂ�D)9_Hl���2�%�m�{/��YPP��"���%l��#Y�Q�_�� A`�����-�Z��96|��d%�+$��m�i������jߡ@I�����㠵tx����]���=�\��0��� ���,�R꧂�0��BȀ�7�^�vq�z�B��YB�d�T��ddE�&��@���T��/�4x*����]=��h?�ߎP(R��zoYW4x�j���}iA�t�b�i�M�gRu�����E�u�ܶ�kX��w�wX��
ɻ� ��0%�RV�CA��N8������(7�%hB �!H�n�{��0ũ�81����e��K���p���ѽ4��WY\>�E�a�[���f>}
���_Rځk�R����n��N
X�� yj%�fΞ1�vQ�ދ@r�Ew�}��;�V��K��Vf
�C��)�^ :���m�u�Fu ��x_�ߤ����R��ެ��1�5��+S��"�^s�*�H� ��C1<BנM,_�q�}�q�8v�*ToGK;�Ă�	1Ʃa��$n�J�K�ӈ�������RV���9�K֤Qe'G8PS�����8��+@��l3��i*��Ϟ� "�#�������%RF�J�N*=m�~b�5�&_���7�{(�K�c�;[8��WN�3paC���&�v�}E	��$DCw�6�{��F��@{�ڃز^B���e1�ix�2�as�5��V�� �dEG�CLK�g4%�`�M�hU��=滮�pS�����֎v�C{����Y29j�U8��ɠ�M�nA��ڐ����6���/z-����3����?X$2�� �4���{�5�Hg����(K�5����h�r:b�� ����j�I{2B��Bn�����-R�<R��{'p�è=9�$����B.��o<'<i>����9V{� ���ū��M�Y���G 8]4Ws�k��{���ཇn[��'��],�ѫ���7C�$v��q"��M�K� Q�ha\���
KLV��3�/r;]��7�~_�~O�!�G\aƐ�t'H ��E���[V��>��3C�Y��$
����z]ϯߤC��cN �r��?fq�����ŋ������~Uz�#5��dU�y%9�0�i*�V���6������8��'��&��(x���o3��>G��T瓤'p�u 4,�!�uƜ��ʬ��q!�R�o��Ea[+�s�:�ͨ�v��*��9�O�	��0�}��O7���
�mZ��J�u̎@\~�E������������(�$}ׯ}�8�[#�S�:2�"�l�Dr��0aTj0������¤�V���"���c����|�i��R7�_U� �<�Rߌ�~�eā���Ҫj�(�`��B��H^���3�R0��3]�?��m�<GQ���%_�O��A�jɹ�+��Zj���+��tfE�6	Z�V`��R�K���~��D㮝� `�M�X�P�q�4�U2(�n�����op{����ܦ��)L�� �BN7�]CV� W�{��<plG�B�H3y�^�m���#��ߺ����/�=�]�n�m[������͍���H�v���'5%�[�Le'7+I�ڼ�oyT}�#����&¨A|\�ͧ|x���1vXH,���C^�Ba���(3�(/#�����?ȶp���{�|S �'���~�� X$Q������ID�T�1��?����/j.�w�[�ix�|��T�u~��@�c�t�`H�>&����I~���������6>(����n���7�)X��aE{bc�
K��,8v
$�� �d�d�XI��y�	���g�����g���K۸ǔ�o��-�hǘ/^�َ�YH,M݌jq3T7�ʐ�Ewh`G+)�HSg9��[�<��^��\ Y��{w��ќ��0wI$�ݱ�Y�"����<�\R̈b����Ōk�*Ե�>]/G;{�;���=*ڮ��O��6.���E��򋃁Q�{c�h<�����n���K��d�O��v)�>k\�u���d�f��q� �ףا:��<�L5��D܍P9���.��'�`�z�u{��1��;�fmJ�H0�ט%Z�����}&v���_��'�ctx`�kL�%k�3�\;K��>԰�b��i�7� ��q	�k
W P��� 3ݜ�S^N#��(�T\�Ç�Ź�hR�������q]��m�E�~�S<�zG� �̮������et<Ò�(�^�n�_|�%��:�2=t���!�@c(�J���2y۩M�&}��A�P��h10:�؅4�X�7���;��fG6�I�2��W�1�.P8�mI�s�j�Т�N��.�WI�Bnn�%Wl��n�vX�2z�4p �n�f�[ ���tC���#�}��q廣n��~G7.���E�՘�ͷ6l+���>5۠B.����z�*L�4naG
���LvYz�������A���"g ���Qˮ��\�pOg�����/�_�J�]č4 M���t-�QF��47�,�(�j� �-B���|u�zH��"ی��A)߉�-�Ѻ��̻"�3@@�?�R��;ۉ�oh�_���/N��ijVt ��EUJ�ˢ�J��y����8y�ո��	�r�X�N)�����c�v2�?xpH�����4�o�/�=��W[���6�#���C�d����_���ϯP�1�L�L2*� �5滿�j-�,�ˇ��U���PaṗӁ�*�r@ ���^5Dv,H��@�r�U��1!`_��ٛ��%������S�4� z�#i�։��$�aX�ypN 2���F���r@/���ȳ�n�=�N�:������g��Ͽ�>�+�w���	�%���( U6Z��D�v���CJp�܍W�=��I�H+�Ç�΂��!+(!.�B�3�k��mYZw�㤬l�<����ѓ��-^�H ��dR	�^�u�8:��|b�-E�xln
��B�f:��R�	�_��3]&��#���-w�#����W���F�����2DTR&3E�V�5���(�Dm?�}�H�W���!��"�%�x��7j�~��ș>��� 4p\8��ua�ӯ=�U�BD�<�i(oR�p��7ݺ,��g=�q��i�BnT������+8dw��e&��|d*��!�qn���I�ذ�������4
3��&y��(�L�>!��Zk�����Wc^��d��ިx��^wܪ���i#�r&���T����gT���7��<��	�&�7n�J$� �OP$A�<b� �3�w��)�U���*F�"�N�����E� 6��9Z\����t�Z��������ǃ.� ov�a&|!�?'k�ۯ���+E�$h;&���u�c�Z3U�GX��C~�|r��U>dd �D��j�BׁD;B�^g\��3�a���7��0vs�$\�D����ɚ��Zd^U�
z�A:���-L��	ڷ&����R"$
�~��O����u��d$2B�-�oce8Ux6-w��W���ۻ��o�R���>5�gC-�z"7O/#:���-���'W8�~��xe=�����}h�?i�S�D��cUQ�)2ъ�}�3���\�FZh�<di6U�Ɵm��� ���CʯM��6��O`B�UU��X�4�;��r̇D4߂ ^\��ѻ6������|���o���B�#P3�f-:h��F��A\�Q�B��<�Q6gZ!i�u���O�3�5dc�B��M�[������Hb�j��P*O���(��̱]�:ջ��7p}��+��{�P�g�HV�Agdw������xϟ$�b<K�/��*t�)鮹���+�&0��pr	� �tbo��IH�J���Jq%C�ߠ*���]
��Z��,,�Aei�&���/70_]l��%LZ��7q�϶,N�4[p���;���z3ruG�-9w����go�AP��ŀ�޴{C_�<�KY jİ#\�$+�+:����4W�g������`9��_�0����͏����P�\�/�G|�?J��u/�ne.$���=�����p�s����������"���=�I�$�`��Or���I���F�B�~�o�`�0e�x6�?L���R�Hr�+�O�r�Z7|f���]�-Q�p�K�D����WM]�'�O�}:3w��Nl,a��I�z�h�Z;��̇-�C��;�}����x� ���=@Ot�ё�p�ޅ�g6�
��ԎȢ\Ǐ�g�塿�\��5"g9<� �K��y�Wﮰ��O�A���i߱�p�,��Ht����&B,4���Q�h�TӰ����4a;�E��aj����H2A'�%*�/�P��$�RlSH0=����e�۬{�����^�/����䯈b�g�p���'�i(�09���z��v
!��;:]��-��r���3g^��Y�Ƥ�Kp�p�-���z��KdT+�	����I��Z��@���
v�s��l��H��B�?V9|�R����F��5���<��dE�a`2�NE�ð1���H���?ȗR�]�́�k�
��!����ΙI��^ap2�+��+z?�F^���� 
����.m�~����y����Mfl�s�?`��ԩRզU$/0�lH��^�\�\�U(msi�1�6دr��H+���IBgb���Z$��]�=�-Tj��j�
������Sƣ��X�?;~��`�}92�:�<�[������UN��CB	��u��m����M�D�Sy%}�mXA��#��[SzF�f[N��Ğ!Z�at��S�8�ݼe��c�ma%J�́�o�x�a��|D̯B�F�V��Ke��y�~��T��A�~��%!��Ns�T�7�^�lȨ��a��B�AnNa�P�|��H韚\�����U֏ל��o粅K�b�1�~��FF�h5���&/�
��nڪ�cab�=��t�U��f���,K���|��i���ս�QL.���~����n���bx�d�s_������f}�y��S�7�O��ce1�� ���O�Y�)���pY��$���0�<h����\x;�J`�qo �(�E�������_�O�3� �̝�!
�9����Z�`�/�7)S��%�l�|\�0�zf1/���RX��q��R�BM�W97U�m���.�H���H5�f�YY�_�,V�7}��8\5.l��uE�"��v1s4�ؤ{����;cL���x�Q��^�����<�}�2ͣ��eş')�G�`�0�k��~�T {9�qx�69Zʹ`6��ʨ����m+4��O�)N)�[�]k��\�����e_��R����^T���<t���|��]���A�̡�VC�Y�2z�
ϡ�>�`uMX|��;�~g�����.~�B��'��r�!<KX4���ʅ�[c���݌߸tF��	������?��(
ĭn?�;�^X(keb��oF U]������b������s2�9j�U��OQ��+JE�{���2zl;�S��y�+�BR�5?o.�t�,8T�<~"pymؗ϶jV<>^{� Kn�8n���P�A�{hulpcZx�_��&�yn|�<q�TY�hd}f7ӌD>b~�����6�/&�]�ɭڶ�YQŧ/ ���0ܫ.l�<��ȸ�ףO������WBx1�q�L�P�k��p�"���N�( ;�kч?.��5��W������B����ʡ�G�)��m���4B?��?�p�0$�6	L�铂i1,�5���P���zv�q�����Z�[�XjH��?
���t~��Z�!�uTH47,�&X���#|f���[�v��4L{�m��_8��u@�hcx%�ֈ�=1��S��c�e�/,Ã�%Q Ss�lD�?ɮ5т�T��y���B,�z� �u�u�B�A'�o6�VT��������>e�xG%�1�y��|.d}���g'��K��xE)�ߠ	F��n��^ ��"��>���ś&f�Խ^E=��O0Mr?hj�������Ŭ���Vb�5w�yv[������q7�km�rݒ_�kk>@���6<K8�}�PիB���̊���<�銕;��s�����ytM���������m ���k�!y�	�}�ⵧ�L�+&����d�a6o�8�6hS�����R�c[��
�I�Ŗ�G9/xH
ُ> pu�%Xd!��cNV�������� �+���k�����@hi��;y\�*}pN�49�tgG8MJ�[�o�]5���V�H/�~H���~��+<���N!Y��Zp��_�����a��?r�i�l5%��!�(�=�PEo��<:Ʋ�6WϪ��؃o�Pl�P�ݳp��q�6��o����rj��QΆ�����"�C(	�`��6����~}mz��j�;��8�a���6����6FV��8�3�qg��!*��Tr�/(`��=��gMF%Ѝ1�.'ֆNM]�z�:\�$6I[�:�0$�i=�A����~�>/��{Z�*��݊�w�p3"�Ζ��-�`��|��h��V�i��*���ς��P<ǉ:�Ș�p�"�9�	{��ν�>���ճw)y��=�hu����Ո^Aչi[������4���}��Deˍ@�ic^rsk�+>C���n�U�8���*HCs�� 8�e��<v�X��V�I��P��ʹ~��Gg���u����$� �3���4I�_�@
��;�8
U��?�e�z��%$cU@�2T�𮶅a0�xt���tQN����n�:b�Y�b�JO��z�A�����d�7i��%F�l���EA��z����~�����eqmb�Q6,����I���E��2�I��Yz)1�$�AS�M�OtɯJ�ן%HS�P�oe���ߝ~�>�L1����<v���W�ݛ����+&������)�d�S�7 �b��o&]���<�[Q?!9����R���- �'�hY�w���C��o�������4}.��0����ɭE��R��T���S8y���(Ԡ���Ow������G3�y�P�q�ҕ���=Wp�ȅ����΁9ÏBx��9P�!��u�t����ic6ΐM:�����5�X	S���Uz�r]<�ޤ���%�������t3�����R��������L���L�����P��`[Pz�|���@��	H����eEx�l���`WD��qaʟ��"v-)	����iW�;'���{Z9_ HO��`e���̨D�\�}C8i��9�����R�x:8���:�H��,?���Ak��m���E��߭�~��2>���'��鍍��9�H�cg������\���V7�����K��_d�v���<;�,)J��j`�BtO��*;�o����l���a�8z:�h�j������>ݠ�?�g#�JA�pX�:]��2CR�#zH�,�i�:��DÈ��9��[��f�0�݋�VC�?O�#_�mM~�Wc'�atv�IGѭT\���4=��DU�7"��
 �qG;i���<{�X��#$�fӚjY�[#ޤ��PҖ"���0L�s!^{9���;�]V�z�]��:���t���2�Y�}���V�/3�ˠ�ғ��<&O�&7pP��mt�e�+��ݒ]�䇥��z�`q�ͦp'A�k`B�a��8fYёVPe��V�	S��baf���̘#���KU����m�F:'�Bn_�U���U ,�*9���l
6TÍ�z�:��K�,
&��B��w��x�R2�E�o�%I�W���z�>�Z���v1[�����]�in~��������#ƿG=���U�ȶ�*#�j�,L�;}���x��#Zo��X6��en� �/S�(�uK��Q~VFRk�K�zȎe�����*�%�[�x,Un�i�M�껙P��?9g���@��x!y)��Si�J�;:*6Y=e��� ]�3ɚcs��,�J����?Uz��Ē�^�HV=�g�, 20?��a��GN�A�+m�8��@���� �S�߲�DRR����q9BfͿHy1Ar�J��2�����΢��T�ޑ.�W����\�Q�`r�h��7�7[	�p9�^�}1��+�`�j|D�
K���Bo��)PNZ�Q��q�U�o%/~�UP��ҪUo:}��M$����</7�_��3 =� ia��l���J)�6�,b1`F^Om�ɬ�4.�p����8>�PY����?TNEiPr����kÝ�q�j�����������"�=�(6���{o��v�eur�lu`"�����	� �'��12�J�"_�A"�)��|���w��~`"=}(l)�]ua�Yb�zs� �1�1��7>�(��`�3a�da"�Î��n=�j)\�axA����C��B�ڑ�o�[Y{�ՁX���^����9d����y��$��$���G����ڗ����cW���V�����0�>'��Y�5���/Ֆq�dȮ��JRĿ�}��}(z��N�B`a�'�=��(��i���n<�Q]-k��⓱���*��n�h�3�`�:��~I�L��z�y���ȷ��5�Kh�S���^P"�v�E��������B��o�Ђ�0?[��뢴"'[�	"�!���_q�/��3���~��;����$�Z�g��
�ե��~�aU͹�ɮO+��C�=_N��A�������d�?ur>o�N�RWl(w�|-���fVzPh�	n&&adyf@���	����	=�m��(|NA.T�������u�֎��x@���	�U�{��(����Ԗ�_g��|���E�������0���ۯf����=�I�_��57�J?y3�4a�s���}��'���e��$��4��s��jj�0zI��Rw	��$/�9"?^�
5��PI�ǫ��J���u�}?���ٶ$q�vf�q2����#�G�Pw#��+�a�Xg�`G6)��:�Oϰ�BB�=K�2a�h�p2.��e��k^�0�[�n�׉��y|�ŕYCg(&�������>�9!�50ݏG����J����C�;0�h^�����
�����<�Usؘ=/a��j,��Q�o~�����������/6�������@rf�Xڌ7)>(������3��_��T�P]�A�=��Y����*�L~���:(�.�I�6��_G�w�&xy�ht�5���N"l��cj� $|ʗ���d]T��k ˇ:c8ز��{�r9�Y��`$���#sl~���_|˘�� E0����A������(��|�Q��K�'Qw�=lx����z�?��Դz@|Je��\�l�O<�;v1�D�w�7�����Z�� �b�C�� ��,���_�/�Q����'�X��|��\��TD���NԷL�
r��G�Ky��_��4z���xs,!H=9���)0�(�B��/���ݙ��=�x2У"����Dcߊ�q����"x3D�\��3���͟d֜@��.{\����G�.��=��{�4X��*뽶.��-6�����tbՊ���H�+Q蚺�]5[Jr��}�;+�p�-3�Pί��ѡ��_��	z,R��L�ږ�K�~�q}�;�$�P�R���h�"�O>�2]��w�g�ΓP���%]�s]nO�!��\h���(E��e	��HO!�hj&�r���O#��f���ʭ�o�%����P?Bv ���9����6!w��
46���24�~��Q0������u)�&n
�L��0��"�+�D!����`�҆�Q��U���$uM?q���q�K;�^�tW�i(X��ӟ�e�(aBk	#t,�"?�}p�F4�A�1�Ͽ袻*L:�0?��x�I�w�5�<��{�e�3�X�`T\f��c�#�z=z�.�Fym����k��%����1�*x�Qg�'��|<X}�瞄Q6
h�_���M�u��v��J,RΠ�9α���P���E���`ګ�Z�V1��&�ڸ�J1Ig�B��,� a��>���w����\T�DgW�'�=H�`F�&&F�b��̦Bέ���>��C_�;��� �-mS�.����.%$�U� u��?��5"��������0Ce"���g��!#�����Dx=a�˪���,���]�� �G��zn�c���鰙"S�zM��J��b��I+,�+���1	�=� G	n�L���~�)�.e�NmU��rfa���Y6@ϐc�l(� q����h�H�#���x�Bf '��ٴᑌ�%����	hl�͆&��O_�f�����HRX��B�Xԣ�JOq��7�/P�d��,u�����m����ؽn i��TNlpɠ�ۢșyu���z���$��[�x��l���Rs2ؕα��Ϡ��3�>���NAZ;,.�]�7�G��Y,��܃ {?���N_c���I\�`�ϼo�J�QݶC$� F4&��怉��p�?[����<`��[YY1��r�Z����J�vCO�y�(:�X�3�	�v>^����7�1�W�2�T�/6�����Fc��ʩ<+I�N�oG�}k�֊�˻��⃰��,�IQ%BCr�¼P hX�l$��O�Z�����+^� g�rD��,��	�&@38�_�,?mhM�t��2!�f�R��DT���Wt�l>xE��oH�M\���K������{�C��z]0�f�X��x���04&�k�уe�h�E�z��_?�Y���Y�f���l)	d�XE�[�QSI���|���.���Ƈ���������v.�1��6#�����{�w�s����P8��Z�N �l>��y�� ��O��π>,���^��Ԑ`-n}1�	��#�f��֟��d<����7�Q�-����fD#�����ڠ�ag���쾫V9:!�B� �cd	��&�V�G���0o��䙕X��<korV�B^��JA�g����W�N��_j�� �m!\��� ���"lņC�g�!|�Zp�=�{/nd8���U�da��*�t/�ٔ�Ck?����q{��'�}e�f�X6�:�B�B��&����g���cV�T-�D�Ng�3K6\�u�#�o-A������~�NՌ�S���F1�<7�;����a�ŧ�&�����R��.���}M"kn�.��Ob:.巏����n��F�kW3_���J|j8n�����a��{ �e��s�����P*24��
���흐�O��C����젷+��<�u���������њ^�ۖάo2�;=k�U0�:�$3D��
,�8�z��v����34�~.�O�������g7���B,���}�G�w���~jZ��ޭ�nj���Xw�wD��'��8�4��� B�b�V|[2�G�9O������1qc�(��|4:?k�ѻ3˓���I<}��T��I��	��g]�z٦F)<�j���U�8"){(�(�k��u�V"�Ӹ����۟���6��\Ϛ;�E}e���9bA^ȭ��2�1e78�)�	_	&.�1�RN+��7������������,ҮKhYk�&���1��K��涛�o`'R��\����u������	EF	g�8���p��)�4tQWDgى�/"Z��y�%]t<$����[�u7�K6��i]����s�4�����%��JC�"[�wn�)�;S<��֝%�ye�=�����]h��������A�Ş��$�������k&�l��ZVS� ��%��j���$  �p�F7�ǭn�}�/�)�m�n�F������[���׎-�1�2+��C��'E��Q�\06�d��Q���Jg��T�����7�	r<b�?�Y8У��Q]x&�ڍ��6���xdsw��G����}�LnIwϠ��lL5��v�u�(`#���NM! �"����?%�V�mA��c�|<�_Z4>
�"k!��y��n�x��rɍX<3�jJa�Ϟ�J�<c�͏b� A���R������LP�߯�DA���-}��8�F�J�F"udj�(N�w��*#�a��A׋>���+��"c�����768S�z͞Y ~�u����y�h�-��h>9L�ڃvt,´!J1��"j��r�Ap���i�7�!����Q�Y�:�h-2�E���2�]��d񛯸�Ã2#��+�B����)6S:�t��?��s�q�!V���n�!I��W�	5��b�t4�j��Ď��vsn����BFb@�o�7�m�ox	�U�D4LқQU�2f��>d{N m�p��l�q慳Z�n�ڎ:q7{����ig�e�4�A�װ����Ȃ��Q�� E�ѱ�e��hEV7#]b�Ij'���YN��P�������������[��'�
��B�l����)�Q�{�d<�$9�xG���)ቢ�$C�e�����\s{*���3��/�[4��l����F��|��^��6�mI	l!�LK��.���
����{2��BwG�W�ġ����n�:�"s�z���6ܦ{,@�K�B��<�R��Fؽ�P�ʛ]����W�&��
'��ԃX�{f����2��3��n����|y7\^خ���zD9� �[x=T���v�EJe��K��ɒčd�#� g�\c�9���T�^AIe�@>�iʊ���Q�?M2�p�F�S;s ��ذ�� �^�v�;��`V�{���b
������:T�ǣw+��S���*�x�rv����{�C��rI&�^�3Z��I/�G���8������Bq~�^�Ao�����m�3�X2��\����Jg�b��Il5}��ҷ��y�"6�%�X���43�>��_2e��Gj��J*�R=�V#�����dO�v������.�-2�sq~�⢞� �V�-K�t�N��M���y��|�u�Nvꪭk��CJ8�2�n��F��%ֹ @L��4v7O>���#��X[$9�aOoIC���F��ɂ[�l<`�h�	�>�u��a�T��[�}X41�p�"A�l���v�� �U���c�ER���2hʅ �~�ܭ;Q���,��6�6���M��$2$��\}f0���������&nh�s�sj�Y'�XڥP.��M�VJ��]
�q�����(U
��V;13;�@+���S	�m��3�
V�x+i,��vW7\���V�D��E�==��s�N��~g��!��~�)��q/��._��)�F���fJڍm�^|��f����w�M��(>��pṏn�"�sR+���*�f��1���ͺ�w�1��^�Ƙ(�������Y�< ��L��]=@E$�wU�\�W!�qsyPd�m*W�	����f�x������3-�,�a�ҷmX�#ˌ�_h:s=��_�=�q9�U&R����ޔ�)O�u�T�T<t����#��4��|���4@��
+���h�!8��b�vǍ��x��V��[m`�4���7�笚���_�Nu*�:k�RN�4t�ï�9�
g�ȷȯ�D�"��8�31�d�@��K��K%��j��Ω�����1/T]�)}{�v��z���i��s�;�Y)����hΨ0�KR��h��-��n��~����Lk�y��S3���~T�"O��S�/�ȉ��'��.:��ܑ�//�[&��E�+�6�%0wF�f}։p���(�f8ֆD�u`q�=^�|8d3���)D��<�@F<#���A�j@ʀ�ɠ�t��&�f��*�s�
��P�̏������	®��;�T�^�΅itǭ/T\�u��<
��� }1a������Pÿ8���Ii<�;ih�3�S��TD�G
BW�2|���7�K��}:ml�7��D�������*��S��Aw�
��D#��ٍ��*����9�Ɇ80!�:+ \�5�se��ۥ�!�4�kf�[+nHind���?DW�
/4���K����'u�j?�Λ)ո�~�Xf����̤�K"t��Q
L�x-���_���\��⭜��3Nj����l7�.NI�/M��㊊b�p��g%��CE�؛��*	�N�����O��X��K�0���#M���y�Wk���&�ϲ
8z-�F{Iu�3Q�o�AS:pLn{���N��B�sHﳔ�S��]��%쵛e�^�Xl$�qV�I�������y05���C|R�Gf<	z=kś;x�i���)Է:�M�m�Ts��2T`�1�W����pl��٨,i��hL��}�@i��N6ұj�p)�?����y?��EϮ�PI|Uj�u��j	���p�+��8����Nt|b-���ֹ�R֫7R$]X��f>�E{\Ra8��p1F}�� a�h&v�>%3�G3';s9�,_����vP���l��XV!���˶�G�.���y�&ͪ6�������@��|�y��;�1�4�Z���uݯ����1u��:N0G{I��.F��׎���sB��:N���v�؊]1�a;���v����Ao�^�����"5n�qU!qH
�_���3( Mz��������m�-��g�8&&=�Yu	�ڤg��D��#�k���Љ��T_\XO߭�?��K`/(�2����4��@�^�~AY�w[���I������Ϻ�B*@��
���w�$�ۑeU��W}<H�8�^֢�`� ���<����Zbh�ɔbg�����V��ݔ@���F#��콄s�����
3QL�c)�\��Un;��ŋ��H���+[*ۘ� ex���ˀ�C��i�=�L�`s�+���	���{���|�PD\�_,��#7B9
p��L[����yh,@�m/���ys�E6>pe�O�-&�[%��%E��˿)-�ShOT9U��K�rQ��S�-]~�� ��L�p���$�\�Gcң� {+�Ї
X�0&N(�V�����Q�|�U����Rr�=�Ϩ��s+�Y ���N����L�c�@H
9��HTCOHк��@E��mYx��Ƒ��A�x���e j�ȥ�d33'����})��9����B5��x�`Ɖ��7(���g�g� ,W��w}��~���!�	����<b����A�b����ǓEb�Ry�L˿;q��� �4q/������������ �v��f�T҇�_�a�D��{{�\qОr�?S��6�W"/�jJ�=
H~-s6�q�+I�Ti�{ζS��Wx6xVEl?�OR�V��Tχ�
�1���E��ج�A���)��1{�=�(}��Gʜ}:��=�7���i^�2��֠��J�#�0�ˮ�yJ����#N���KN����ϩΡWk�=A��1�ݖ��S�R
B�U�u 0�#�Ր�'R3���v�'��@���k���\
�i��P����;��N����7��=6p�b��GZ	GQ�BxtpA�!���)P?!��4M��c�Q��|ID_�HI ��,�)2wݘ�#�\I������ֆ\�44W�җ�}���%Px�66�~,�V��v�\���"�ku;�\A@����AQ���;�E�� î|��Oj������q��g:�>��A.�uR�+�e^�Ɨc��J�^��`�^�
�,�-�Y���s$��Pǉ6��+"�kWT�aS�	�ςa����n:�������g=�)vL�j�	X�!!lX��.(�n�QI�G��Ł���Ae�Nߏ<w�s�m����Bȹ��%M�Ʌ�Z�m��0���w��{�Ú�VQca�_H-1P����Cx��������[� �~�9����~�c�r�<��U�9Fd��IՔw��LX.��&l�����R��u8<������q:�O��� �J(��i����#=B���s�ӥ>@��84�B�fo��O2
�%�Q��4�Y/�x7��tK�NT����[u�|� �#���}6�;�G�iJ���.a�,`��I+^�,w=we*x�yj���M�3�7����"�������+�vw�8 �C׳�s7�A�kH�!�7�/zF+�w��k���ip(t51���>��ieeBڄ�)3qt��5�,F�H�'hP�`�j³'r��a��_���<�g����w�)�,O�2x?�f�p���&�eTl����%�!P_WM_9N�]��n� �t�è"��U�Z��mB�Iq�p���R�0�(L�%��9B�QN��D��'������)*��֤(3��{�EJ�.�:����"�#�YG?�_���m��:=�jy�|a'��e�t)HEʊDg:+���K������'��(�����_���X�MB�&�s�`[�&����-����e}�P�j��OŬ�~� �G�X,�<�ՙn��Ø��36�� �ؠ~��4?0}3�$�[N%���OA�=���\\L���_��c�y-����;����K�K����L�[Z�V�H�l��ͼ8��tQ6n}� Cٴ5�15�v���lvϺ#ԩ�lV�;�Lyc��F@�h	���H}�^?(��&����e���|��9B9ޔ�G+�K7�#��^��?"�-Y�m$��O$�g���C���׍EN�bj\wWC��r��E�4-�Z��s�e I;��`��3�wTa��ɦmrz�	�t.}����n^
r2�7�!C�ת��d8�qR�>ٖ#�w2����.�������o�,��a�I�Z�v�C�	"T�<Z!J[D�����3�8�i�ȥ��!��,m��N�Y�R�)u9����h �w�{�Y�P���d|����·,]�K���8�h��q���hŔ�#����[�v�ZԱW1�F�Lr�Tcyx0!
�=G88���ӊ���s(��}�*���5�	-��h���c�]��O�q�db'��`�B�x�S����������V�(:�� ���d�g�ﰌIƀp��G���Y���w<���,4C�6䝁T���n�k#O9�R�?h ����
��Sg���@VII�Q�DCE"��8��1V�:��C=cHFe;F�r�7X�	饝E��8����(����(��O�-����].�0L�Z�Q5��F����N?@�:_}@s� �Y�S�H�p�p/��[D���u��������������<'�h'nk_�T�QU�8r�*:��m�
\�Ed���3�6���Z��S���ԝ]��̻�(�sMbi$��같#x:]�<�fFf<����s�~�Ɓj:/�x�3D��o�nP���,0�C+�PY���g���^����-ʈ%�q��4�5�Xd�2�>Xk��Uh��$V@ҼD�LY��t� �(��0��Ҳ�Q���5}|����l4{��R��J�,pj�<Dx�P
���>�W+$f�%4+�Џ_��Pl� 1O�ʵ�����ГL\���^�}TM�9��q/��K}��A٤�����y�j"���*�U:~�F���]?�i�ǆ���<A��^������H�5Z�
����N�&��g�o��~5�51P:�G����Cd�Y���uQ�{���0~�7v�
�O$�����3*{9&��3܁�*�e��Q]O�R�9��}�y���R$Y�5�@/�(�#
j���S����a;C�ϏX���������6�CG�l.[��b��r��1����K���X��<@
G��f��]�?^9H�|��Z��CZ�b����mz#�����Ó�M�a]�M���N����,�B?N&z�Ը� q�Q���O�K���z�A���X[#'Y��I�:0V��D�zZ��@ݯ�j�fZ�b����7���Qj�A;������0!��ұv�?'�I�(y47�23����E�h�B���"'+����Ijܾ�X��C��3cʎ�m����"\<��Ez�rs�wiR����è/�=B��`�����=!���B�Q��A@e����SI�.�9�
�6���e�]R��x�;��ܷ7����^��4Gά�AU��H���B��ϸ"k�n"B��rR�i��̈�m�*� � /w2E|ύc4��~!��"��d�>:�t���^�ͳ9�Հ�E����Np�l<9��kl�B���e�A3j��Yw��F���	n����e�nK؝���M�8Rh�{���g\m��-��j�őQ��hΜF�s0��&���x�4^���/�źp@o��Z�� �+�@ܺ���((�c����]��Ӎ��3��Y�3x:���҇Nո�i����|���ٍ�)�&������r(�����9���v��F{�zP�kB���\�~���[x?/��*�D.�������f:W����˓����|�������uQ��I��]���R�g~p/��J9�ϫB�_����� f�./�Ek�/I�xb������Dp�������Du���H|`f�o�|����*|�ժX���~�C�zh�Q���'��e��{��jo�$���{��~Su���J�����$��i���At��,���x8��ɧ�.>O��/?�Zo�)�"�-X�-�H<��=����@"��Û""�`^z�;O%�/9e����Ҹ����
$��:"/׷j��=�Ľg��`�J)O�}�I�|l}�w�g��������f��FQ���K;K�i�	�^ߝ�#i&�����b��w5�9<�6����3�|���Om�7���-�}�q���ط*"R��s>�ZA�a<�u5��}�I���׿:*xRyM����[�f��a�V(���iT��ؚ	ßl���"�T:^��z�K�%��?E�8�I��Oi�u�G�U~'��LD��*xR~� ��<9���q��g\���o6��S��M���̲��B?쨛�f�M�z�F�bV,B(1��5��]*�qvl��tde��s����C^���̥�*ǯ`p���9 ����0����Hu�?��N3����O.���Z���&�D���+����=X9$�D�8���#T�R�B��pkOo��G�\l���"�l2�fk��ֈr#0�)��t�I	G�͎�nPC�C�X�Ʌ8n��6*31QS���	�3u������7;DI�i����&d� �鷃���1���n���Y��1空ק=��=���u��B�%/�=κ�n�bz�	������pV�q���U�O
�W����u�A5�"B��q0{՟*�xwQ��k@f����8f��ufc@C�>�R�ثc!Pg���� ���^'��O/e��S%��m���B}��5�.�Χ�Կ�AG�o!5�H�C���'|�h�Z�e����C���\3�CW\|�鯶5]��Ɂ��MC�|��a�5�t�u�`������'��2Hw�}��a��$�S�w1f���-�)�S�R)��PS�>�#�]���@s`��}�Y����J��s�)��3/�Ґ��
9��k�jKϷ�H2��恞7:z_f�`��c�)���^�ܾS��T�m�!{����n���������h9ٮ��9ˍ���9������o�!:D��ԅ��&��i�������rB��CK(݁Ŋ6���R9ʍxXQ|�>����E4!Q0%�z���W�[N� M������f~��!����iq��%��s�2U��u��ꃼ><X�}�ԪO�������KxI���߇juNPۆ�ُ�}�UL�>���H�hI�b�aG����Û����h��rD�+�F@W>Ii@k�,n�������;��?�;�X=cE;�ml���)����"Az$�h�cC�6(ac�9�je�([F0a %J�� �5�O��%���Q�x��g��}�X$˝�ʥ�c�%a���^�M���3�^�sh1y,�x%6[��cZ��U[�ZS�pkѰ�E�4��C���M���\�D!A@&)>�$���3+,� ��el�6��]8��=_���Y���+|�B;�$�!,sbuN�4ȣ_�r�lSJ��%��/v�ќXa���H�L:�;����Kr\�����q1��S̬��� �C<@��:	���qp4�AMݹ��	v����*���dd��7�� Q��VH��u��F#���S\C7'>�i��(����{M1�L�
�3�-Po:p��s�Mw��_�42[�.��Hmv�o-�lS�xM���bw��/�z�_����c��.�:��c����ş�ŘY"	7�g$�F�q-��/ﮘߣX�~[�/0�2,X����MY\��-W�á��t�W����ytI�k��;�8�rF��.�M2.�M���>��Vʝ5��L�Ä����������^ h�+]i���K����b.,%5�N��w(����(�F^�L��D�}�ZVg\,N/kR��b:4���9�(���w�J�]'�m��|�	����cM���j]��NPc���
7�@&^���S����He�%z�o��BF�q���@�Are{���k�����G,��q����R����uOĂP�M���07���ux_8c����\�L��ץ����bha��|��yu�ߥ������IZ��s1�$���%��_A���^�+��w������\���?I�23@#!?�yO9}US��x`p�&��>_0�k����3�Iv��粫 {�v�]���l�����dSFo�����k$�C{�6�bo���I��.J��g��A'����Sp�,�V�@ ���Λ����߫ƭ(�x�nc4,��:��W�����wC��+s
7W$rMt)!�b<I?v�B�Bv��w�x�!�11P	T��' ��tW.,��,vb� L���M܅�D5������+o�$�[�/\גc�>["%��tv�8� �|�}q�@�|˴�`� � �i�d��������E`M�5=�}W{W�҃_v�I���>�zsL�����em���e���_�Yi�F�Z�QS�#����*<~�j��["�f���	�p��N{^�&̀��o-�JH �p��զ�;�SWR��)�JA'W���g8;-�W��u?r����	3�c��B�Ʈj>���x{d��a��g���,��.2�9iۼ�O�ƞ)�Uqt�K�J�<5����NU��n!���z�����-�ۯI�O�Vb�$�Q���N�dr�__�����)m_��1�u�8-��3 �MB*V�V�Y1 8_��~F[�(�tLn�@����b��'��Y�_�u9?����e)��xulhAW���i����C�zR	8��c�s��q�~� ��C`�H�>	��mQ�B3��ԣ4��<�Q������A-��j��潋�1���NS�$��U�����ͤ3�1f3>�7�&�3a]'LՑ6I��<#<�6��b�.���9��	��?���Pi��=7u�7D{*���`n	�.� �-'h
o���*�2$K!��Miv�ϥ�"�:L��OS�lEP0�,ʌn�h��0w[���_�R�����V�ǒV�Xo���b��|[d�0�j�<+�}x�n�>��Z�f�?&}�zG��X/�q��P ��V���^�&�Y�4�����S�2|��N�U5Y2�yr�韴]%<��-�E��3 O4̦��B���zg�������i�=�C��I�Z��T�A{w4
����n�I�x/��d�z�J7���P�}3��@^�̏�MTO�8��U�Q�g�yUE�][��,sG!��ޘ`AU��3�9H]��ڄ�*�9�1��ӿê_�q��xoˌ����G���<\��:�eo�����byC�ɁZ���ڤ��Yr4Ȗ���l�)s2��Ld��T)"|[K�&r
�G��d�<�]�F���	�um�'ژ��n�@�������J̜i�=�6F�`��Jl�����D1C�ay�ϸJA�!�4�����o��t���_�jp,h�
uf:��`4�f4&/��Ȯ�}*X�!�S��G���~�rʊ�6������Ţ
���o/�B۰H�LB_IDj%,�h;�� ��&��	�%�3���+��9���J�^��YY|D�sצ���1c�7�l
I<;9%�<�f�:����lđ�*�O�13ǤU�i���~}�rͪ�:�5?��k%V�BOy�������.��e�h����~�ȫ�u�*�oЖlHu'S�vގi��|����s��T�D%��G�w�5�_m�ӺT�v��ju|ӋR��􃻓 >�T����AV,�[��5��*���{ ��.֬�1="�Q�.�
�=}��W;�,���!b�l��*,��u���QrN��.aę���:o��\��D�r��N�X�����T,���)�4���7>�;w2��3R�#������8t]�Y�7�d/5?rc��rگ�W�p�K��8H�N����h6��h�1 ��$@ie8���*$| �"�d * �g5�̝X����^�k?����%�>�v`2��whN�4-��CX�!��g�C���er�rN�\<���	]{��E$�x����Ç���>���Z�N�uB#�zNEL!]�x_��>Z��E]
� dlŭ4��+�C�R��^��Lm9�ɼ�;0�ʃ�H�/��FԒ&�vI�QRY~����ov��vt���`X�M�V]�_��2M9ZU�u�]���T	��i:�5�A��S
���s�9Sz���Eqj=�߬B<sR��:�'�j��_�`H-;�7-�^��ڗ�m6Ĉ+�ݧ���ɀ�Φ�S=��d�/�Q�����'�	[h&\�ߎ%��X�J�=��>
-�$M���r�*(�N�������)�ߴܶf�H���,n5@�!ߦ�!��IL�n�����}�pǡ�e7tn���7�R���G�Џ����W1��v�+�~��(��>g��,�+�'vҸ_��dM�YFOVn�z��� �[`#���Rs��<.��-�->q	3p�&
�� ��2�A�m�����Sl�V.kI�N��r��?͝�=�6c��B�H�8�%�A�a�!���hu ��MR��6m�s$zY��n|����8�H�_�À��k[\D�z@��b� 8�Tϲ��Z����7eT���/��y�$vi�֪s=�{��0���R1���p�ע_g�$0S��'�OF�����������׺�;��V�g8��L��e���ڔZr�����ha��JF��E��w�8�!����Z7�O@/�b��m�g�3���+��=�h��,� �^�P�gn9�Xb��iLwN�??�ܼ��
p�8M+l�yD<y�y�����ry�'ҭ
]�
�d)�{:�ؽai���a$,x����� g ED��H��X��W{h�%02b��Dl������$YJ����S�LA��ߤ����Q���IEq?x���۳��ܴ����|�,}_O�W�ޣ��֭���oy�6�#9���o�~Ϫz�x���J%s�^c�	/�y`���D��y�ډ#�T�!����u�~�%�"��N�`A�瞭����3�*hE�mlH�1M+��d"8��M�H-C�y��h�۶ī����S���aD��0��� )�6��)\�}?�ųl�d{���\h�$����	9���E�꽝��.#X����:v��(#���2OmKp.k�=dma��yN�ig�e)�c���ແH��T� B)�&�Ln�(�������R���C�p�X<��LɮoҠ�66C�R�w��F8�@Hc��Q�C�?���΄e׉ey�g�b��50d��� -7<���{�KP+��А�	��H������G�����(� �M�Խk����D�o�w<��7�Y�k�G�# ԉ�h�t����S�!�z��*����y���o�����)�*B�;�E?�v=Z)���D,�͈�{$��.�b^EX1���=�Vh2k5$%�iSS#��ÔUX�������2�<lꯌ�-��7�} %�Hꪓ�X�#��]�Ll!�ƨ���4tˠ>��H����/��ss>
�bc�H?/wFF苠�2�;"��2CH;�(�6F�V�1�~��.%|�|x0h�eW�P�[NC>՞�mAH�y�LAf7��fN���qCP5XT��	�bb�vq��0�5Mw�	7ߓ����@�~2��]>1�\~�3�F-^��V�O.��:'w�a"+�v����l��~���*O����.�Z��t��i�؊�ٞ����l��:F ����%�g��:�qKw��S��k��.�箩�ym��j3kP/�'Ϊe&j�XT�/�X݉W��Ui�H����V\�
W�&_��)�
/`@��_OM�+Ē���K.���'29�*b���~�qC�P�t[3]��c�pD��;��ҍ`��������4�m���q��,�	���`���Ia�9�����Z�9[P�5@�I��}
��N+�B�9���_z�1\A:3˅�^��Ղ}(ͼ�仝�O�������w=�V�%��j�G}�uO�(�����.�M1>��B?cRQϢb{(�Bc��ɜ���(���
>'�����7�K� c�����|�,��5�WQ�oz��t��Z��}De捶Ӧ�:fP�'Gg�������1�G�k%$'̷|�&y�1x^Bqo�����l7�����N�cH�`'w��ե.*��8)A�1���]݀��~�:������-xlDC�U(G�(.>̑:e���g�Y4�`AzQ�[o�2�))N������0H�l���'�s�`w��k.0�����CEh��au�6�� 0����y��<{kQ�v�[�P��AUl�^Ϳ��.���H�ʻ^���G�n�iy��|*�͏:�v���~P�ol��|�[r�*fi]��"����b�B c{k鬩��A��'k.i�qF����k�ր��D�KZN���������@��E�#�/�6�|l
��AtC�L�@�?�"��,ӆ�de��"|=/�T��9Un{�L�s/��X�Ih�U�3���9Zؾ���^#JmEJE8���ϟL�8�}u��������V��}Y�[�w�T�nD�璋kc��ɰ�z�>)^ErG���ܶ���!���oSՑ�Ʀ6���1Eoq]q(i����Ó��9���F��� �,""�EQ�z��w�V	V��K7�F�Nix��BP�!� @QjM�N�<�R Hpۑ��EO`|qG.����t�A��q.�y�Q��[c�`c��ɜ^�'��Q-�U:��6�ifᠩ�vv�K߰�f��XC���Od"��o��3A��P�߫��'ϭ�M$LW'���+��)~��T�&p�$kx�g!�"��@B���[��=@�%n���Ō�S)R�@X~�&*k�KC�yN��W�ASoPzح`R��3����)�NHa��@��E\E�bӕ/���B[��3�s9�S_ue��P#�XE�De⾢��x��!�2�|�YIe�u�Ȥ e�����j���K��z#�q��,�2lY�)u�f������ʶ�vH���e����������.��M�s�V,�r��*�=K�|�����Z�Q�AEr4�Ѻ��?i�n�2��d���Hd��<W���L��s4���nˁ�̟�����;���k�ڭ�T��/��ֈN�^��`�� ^�'��������{c|V��C� ��Ô|�% ����d��1Z�?�5�kC�ML�k�����W��L����\	~_vgh}��e�kYѡ����]E��Bbn��isd�xF����If%KT���ƺ:��X�@�"�
a��֣N}��%l,+/"�
ɭM�����>,!�S�� o�Xz�2��{��Z�A0uvi��2"�W;8�R�1���%�ٗ��~$z�;s��+��$#A���fM�W�SR�I�+{8�� �t������h�u\�42
b3=%볎Jƒ�J���\����Լ噞�9d�K)i��D���?3i���G�1��c��b&yg�.�#Y�@����O��w�������&���� �,��q�l�%��D?�D/ gi��U4�M\��$���!�c$�`�e���ُ~<��(��ŜlI��1hb���8盀��M�r�{��n�K7'��溺K�y�X�҆]�Ȳ'�b7�}��BCuMJ�݂��l�����ޢH�>:��
ƞG��/�`���JބU{���7��n�;�̲��u
�JpU{'���I�SR�J��&��H2��5u�[�dX�	O_������S�ZОk��B�0�-EZ-�cI�yk6��|�2��g2r)~6T�n�;��w�
�R�@W��6;�IJo��(��C���<=�R ���vue,�%�g��(<2��̛�x}�o-VI��8N�efw�;��Pl÷�.���9K��0�@��"d�p�gRq4���]$T�!�n� řQ��������W�rYB�w/�q����[-c+F	�Ke:Z��~�B��G;�؆�=���bo'���\yF��Bz@o:�A�W�==���[�dz'QG�h�dz�O*��R��'�|/N�"�3�(���=��H�\.��\z��O�Ue�4~a��l�����qU��B("�A����]���%M�,N. ^:R���i��/Bj��m ���6ly�"�±Ч�ʗt�����}#�2���(�"�j��`�Я�+~�±��tf#m����5=�o�su�4n���Hc��`B#t9�ʂg<�������f|7�������;.`c&��r�jɂ��O,�X����[K\?��{Di;��P�P�wF�=ͫ܂mH��I���|������_$#�0�2�&��ʢ;�S�w���͏�y���4�B{�,�v%�tԡ��,{ (L�r(!L�z���K��u
��lzO�D$`��u��ty�_Da�؝���&��:���O��k%5NQ�/Ր>���0D���GT�(/���j�;s#cq�j�Ъ� Փ������ΚZJ�C-{��gg��Uʯ�:�B>GU��w@L2��;֏\���W,��5�KG+Q|���0�'2�d�f7"dFj
=����.��l�"�j���0�W�k�tĳkBo�"T-��|�_����F���>ٺ��3�ȯ��=O՟݆=yF�<;dӰm��&���W0Wf\�����[!�� 0�����=�ȅHdw����M6�V��D�\��?��+�~N'ړ���C��<���./D��.�Yv��i��u��lt�~�ةŬ�а4�K�$�֥�c����S�{��w?�H�#	���^��Չ�*fK���;�H��r��.h�`ժqщø��Pjߎ���fAN`��]���:��)���5T����"���+#}b��K�����l�|�|(�[��F �a��`I���	-���
���b[SҪ *�<��S~��x�F!���Y� E��9=5���;�l���+�?�7�8KNf�vM�ЗI���9#�Q����# "OFHؑb���Y�@��x���E����2c0�.�;;�}0k��,PN;a	�a�?�\�I�7�&9e���nf~�5��ĕ��U���y���N](��a�c0p>_m��y��/��p�w<���0��3��ӕ��S�E���Q�[���&U3�Y3�f#y̈���؜S���E����_��u��r�j�/Q���"�M~�Y�L[�������\8�Á���p�* v�W�a2�l�q��h�U8\ ��$���u�6-iR�d^�' ��:@Z�����L/�n:4��V��p�Z��K���v�Y����Bq��޻Q4t,���qO�Y>鱩'���e���ͩ�f�i������"�#��fb�|�Rc�/
�f� �5�)�%G$�djj�5	��i4-�P��������b��=̝.�f��
�x�h�m�,fe8B������{[~N�fkӜ(�U��"��P�NiP	���@K����8h[%�[
o��l���1�i�ƞ�;(�Ӳ�o| �H�H�p�STI���.���Yj7dQ�:��¦̯��B��T�+C�}���Dv�mV����w���L.jQ�����G�+ٽj�Yjb"��.G��R/u�5��96��pl����E���c4F���olw�q�����	"@�C�w��Vp'5&D�ב�G4�N(�(�$��f#��S���	�I��X���������m�n�)ۆ���d  ��saY�ȉ_Ƞ�5~-�r�WO3���_�L�x�H�!:9O�R谩m=]�x� ��]4����$����aNtUNcMQ~
�@^��p��)�v�
DΔ���ң/���gwe�� �5�bY� c3�=���M�~����Ǎ
�4@��j%��ܘn)�1qSXuͩ�=�#&8�&%*�as@q
�.��U2�@w�P�0�N��[�fVA�F� �/�M_�Yߺ��|U)�Z^��|���z��r�_�ŮW�M&Mh?��:k*������H����7rV; �j^�{�?J�q����� S��K�a�ߝ�z3���b+�*�eG!��p�8p\ʲ�w�zrw�_L�7�GptD37���E�dN�|q�Az�KG3�.��"P�����ҖT&u��p�ޝ�5�@iA��:ܔ�L�M�)淁�R����7���R�lw11|����)�zC7U���j�|�0�I<S�;4�h�A�m}�jP0�c1����)̃]I��L4����z.�k�_up~0�ˑ�>��hl�wT}Sf�y��Eӻb���Y�Fv�`Gě�)�?9'М���Uq$P���̏�Me��pn�>n���oLI�c�A@�KCϴ/�\"q�`�Ej������V�ɂV�҅�{|n�^^��o�<l`:�_�[ݲ����9v�Zcd�aJ^�#L�:ϒ�H�>�<u�{^"\��b�>l��G3�
̨����
�+}�@~���,u"b$��}��u[`��rr��E��s�ا���9W`�qU�.�k5|)�tfn���$�E����C�W�֕Ʝ$�ɰtCͿ�n�G��4��rV`�C1��x�ٔJ�a�I�y,z>ۨ�&D�~�Uh �M+[0%�Qӂ'}T��jsS)�ࡋ'BW}3��ßt�A��Ucx:�2Y���\p�F�F� ��S5u�&j7�3��vI�,g�8~Gy(��[�Z[�=c���8�i=|�%0*�N���6���s!"<-c��A@}��i1�;cH����hqO��pO�rC��x�j��J�& �LiW���@:���}DVT�ܝ��9Q<pwyQ�ϜO<X=q����D���1�ҩ!�4}P_�����7�~["p��n��ek�9_��k�9+�#�����:�#v�7J�h�p���ʬ	x��'�k�
y���$ Rj���M�mi砪tP�!G[p���U��?RF�2gd�D����%u���D�;��I����pnJ�lQ�+�ͬ;1�Wj��C@��}N�^�F�k�ޘW{(��+X��As%Bl}ߙj��>c��1j�Jt���0$>s^��V��;jEv���Fu_7L��*MM��E]5��u��"U��Ce��ퟔ�5����P3��Ѹ�ٷ�x����Nc���@DG��0�4��)]��LYh�uЃO��ֿ���&r~H}�@~��g��lI�܉�����EÙ:��rSi?���
�{FKD��]5?�O��#f�`5ݙ�~�Z���\�>8j:3��w%<���'_��^@��䨔v�:�����'� �'OX����a�Z}!</Sk��ѥwG�QjEt��c��*T�W&iM����8q��5�8vҰMWذ��F�!���%`/��נń�����g
U������WD�wz@��OK�Ԍɡ0�C.i.@���h`'��YHjq_�Zz9]�^(���_ȵ
��$E������y�͘���-$�S���(z����t�q��)8"1�b�^�A�"LA�o���6~X�@̛ѯFF�G���.�Ɋ��X�T�����K��H�;�lP��')��Yn[��1�J!�Ş��=�%� ;xp���i��^"����?�<<?}���5N���Sn�8�a���6�|��S�R�}&�Oߪ�Y�և ts�?X�y6����U\����v�]d����T�͘�/�9�grxJ!9����kڡ�M�ԯ{ƒ���o�F�.��h�0��<݃�j�1ӺbX��:��Q��Ő�������R��{�w���O�����y���d�,>N��i@��G�v1�	�I�<��HYH���>RcrF��N��ת��f��U����1xH�JJXwc�W ���O6{kC����L�[|��U�145�,S�Pc>8R�?�l�Y�a�#���6T�z�e1Y1���C�1r�%����tE���ۆ��o�c<�<\��K�(��c�y�U�0U���S�aV N(�? �tq�KCP҉��M]�)���fZ�:���T��/EE���:��;/��4|�s�w��Q��I�8c�:HtPǩ&.oa�'Gp	��uϜ���#o��Br*����K���Y��l�� p�ű'�x4<Pe��lj}���wPg�o�y��.����^�f�HaX6��S������sw��8�T A�Ψ��b���9���~q�l�t�X�	n.�f%�\ٶ �Ү:(�ᐋb�(�2��	2L�������ez�^b���y�5s��緿�qW�!���@���e��R������m(��s�-W��F�Ս�ol��k�#��@�rykm�e7>[��&S{��	�c�y�ұ�ל�+@��~HTQT�/�莌Ot��~{� ;i�~7�h��}�>���w95�hūk],jN[Ĝ��ڵ�^�=��,Q��]�x˗j�#2x7�b���A,z3����@"ŧ�Y�
�b"�k	��p�	�؆C ��U;��N�[�IU�}U�HO��ⴀG<�`��N �&��t�#����Ċ��è�C�h&�)�O������������������^�j�R�A,�R���K�!�1�4{���X�Zr�1�Wi�����Fjڊ#�C�{A�
e6$�o�^���)j`O(�8����ޠ���R�J !@V4a.���t��>��nO7��z��??>]�f�Ч�.� �[Ӿ��Ԏx��3d0O�2I�G]����+��G��#k=ϊ����Z��{UI����@	��J}�y�\��"��q�ۚ��w��&ڞ�Xmv)`|�ce�q��\X�o	%9o4}���z?�'p�\��p9�w�\ld6��l�������Zge�����n��;7��W���圜T�����F8��E
�y1p1��'�~Ӟ��Y�`A�43����@�p��VdH�k�wj��GG�������c���r>��rEa+�T���F�u��B��?���_�(ϔh��\�M�f��X�bo�2��(R���X��3�yф� ��M��/��#��6��B���!.����ƛ�0j!j4
��/�ÒAuX�m��ez_���4cJ���[Q���\�� ��-�+0t�ԩ�Z����[l=�����{\��������[��� dH�w%�ǨY�,���6���N��n�9[��(|>�T�YҊ�����q���$גnYv_,\\
��y��D������ߊwfo5L8�䓌���\?(��s���b��
����8J�U�gU�f��ʇմ^J����2쉝o P��愣�'��/�-�s\t��޿�|2ufhkl@���`�6����C?m�"��6"	��D�����b&ZO^���k{��c�����E���'V�G�#$��}/K �+Q�JFA�
?'��!]��Q���"�2��N	�ARAx��>r�8!�E�*�)�AT�j����P��1�#�������fU�2O�٘h���Ԃg���`%('ğ*M���CtL�0������a�]d`�/�M�z���
�E9'��s����β���~n�s�X��9�AU<���n�3m�{��
)����z��?�U�8�I# �\n���6�ɋ0��5���Օ���ٯ�ڏ샳aN���ۖ3OFxC8�����3�X��uY���hYԁ�*X�����UR�������
�!!�@n��*/Kh�������e�DbGMLw�[6,G��W(�b���/FG*ҍc�1x�-O��Ht�<D�U<�(�.��7A�C��-HW�3a54�$H����@@M�T���G��z��T�H�ڬ��1}�ڽ�-�n#���P������f�K��7���5���j��Q���!�!��9���/
��*dn�*A!;�]�YPi]ʍG��1�<7ũ������6�>���y�3��BφӀ�-���^�hqV�܃Q��� ��Kݤ�����;`A�U{Z��;tbI2x�M�+��)ZlP�����}s��H=M����?�EC8(kB{��G"Ƙ���X`J;������ϒ"�j�ޑHJ���H�E��B�`&��5�Ђ��*�
N�L���N���97�����	��(���2}�I��.p�ʙ ���f8h��mu�g�j�d�����z�<���m���[��˾\E3e�P�'��5pɾD��c�j��WS8g2O�"�2w�K�1"�RG"1�}?�>2����9~Ÿ�W��]7v8;���%�rM
)��j��,�1Uaw{I�V�uCq��7A)Ɉ���°x�4�_�up��v)�j��	������Z�_*���J��iD������%��f�J��E�|i�8�h���z��e���xz`�l�z�+��L���fT��R�G����e�V=5�&�+�L���ϰ4���@C�D#Jh�S�;$r�TI��l�B�_aH+���Lf~Y���TV�BX_��X�'�az 4���^e���% ����|���?m&��$��t�o,ٹ������HӜ��}4�#����.�kҋ���ʮ=绡~��n޾�dg��_\S?|y���t�[�M�;�r��nQ��R�wI�Z����M��z�zF��Gd>c$E]l��}G�T萇iq�9I�ޭ�\�G�����Y p����[Z��C<��3�h��qӑQ3�cAM��T���-�b1�y5g�������_�����G�2g�Z���3qC�ʾӟ
�YH�<х�ep�����F|�_�i�C؇R���Y��!��Ƙ���|"����N%D�3�C�r��� �+<�^��lۅ}X~(�L>���4+M�1u��1�ޘa��0c����¼��͜q�'5�"{L�^�A~;
�t��'�ھ����9�}C����ܝr�r����D�Ȃ��nd9�H��[�3��U�R]����j�7zʪ���_ⷻ�.鑞<�C1�G�`�Nf���`I	���@�Z��X]��ý���aȳM� >_��D
:|�+�-%;H�����e|=�qW�
pk/zѺ{7�B�#���B�6��L�<����Z(��g��D+�M���h�C8�=���:�6Lp���9�V�p5J�M��s�/�jn|��_'Z�����r@V�W����}T�O�ab9_���98 3�p����ֺ�����؛���0G�ѳDU�rҧkd�2ԉ"��]�ow\ڟ�b��Y� ��QPM�����#:�~J d�&�
R��u������%�.�(7���T�`�`�;�m��JȤ��/]>���u��W���`�nI�Gיh���?&X�YsA_��!6�?ˬOX�m�΢�3I(��eT�-%x���\߽�.	�9�-$�Y�nLo|�\:6"�ۜ�L��8�
+���!a�}�Y� ������Z�TB�o٠�j�2��*��