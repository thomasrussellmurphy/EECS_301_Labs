��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\���V�fnvx��ÍG_;�ȅe�~�>���9�>��Y;�0G�J	m�_�@���t��$�F�FUk��T	��+��	6i�*��1G'h��];�P�1Z�m*i�&��o�_}b��1��.׊�Dħo;�l��"!Y�1":��k�����B^
 tj
f��_$��,�v7���o�c��_��j<��<YJ	�n��9�-WHsċ.������"h�d��	�����yo�K݌�M�cN�����P�X�5�.WtZ�9����L|���Q����6h�k8ڰ	�Q-u���B��,��G����߷�X�E��C*�h���#��r�_��O%m�`q�*�t|��C~��f���q�����!�S��B���Ђ7e��K��#����{�Ȉx�a��(������#���_���p�>. *�W>A$$�����|S ��ܶ��3>��XZ
kX���ᩳ��'�k`����>8�QjWgJ}i�^f8lc{�Y�+���c��P�W�����[r�an"��6:�������kV?`��]Mo�%2-/ӹ��=Y�R�,m���s/`]�o��1��M�)��ՙ�Y��o��ns����%�R�����u��O;y�|�Ґ�v��Z|�/��H��{uxh+����P.�'I�S��*+�'��)/�� ���&r.Ξ��v��2z�Y=��5����[҈�מ�ܔN��94�����U��5���X�
'���[� g3\����-���W�����ÔS��5�}{��f�v���ڟ۽ vy�[%��?��}�.FN�q�u]��OEvK�;�@��$�#��%���(X��s����YƩ�5R�ř�@�l��+��-{u3��C�|��[wo��M��ɱwg���Q�/��Y�S�?��eUl^�uM����jc��#a[�ևucj���|<�u�L��,����ߢ=;*>uU�rBz�zD�� �d/X+Jyb���HGV`b`*
)�������z���<fX1%��P_"L[v�ӬV�x�6��?�⬯��(�V��1���!��[�ӮО=���#{N7u�����ʉ�J���+X5Q��[0�'k�6�^G<��<�}���m�r��^15�Ih�A%gK��׎Cf����0,��w��Ё���rMC��P�P��$	H�
�nڽ'�YO~Y7ꠠe ���5uh���Z����x��&cR[F��z������0����]���g�!m,F�A��j#�t�ɹxK���:V�E.Y J�q~���+�bc�T1�Q�|�\w+5
�3���������SE]�@�gm�K}R�ɖot3�>�ߗ�v�FVI�J3WkV���bZg�A�\[�e��|�4,#�e��s+�>���T�r����o��w0�=��ܗcё�ǆGe%R�R������Y�?�D�h
�ʆ<��\�X �� Cm�p�r�J�b�p
� �(�nBF�ojPs��:jO:��8�"�
�xRގ	6 V��+F"�^z6^\�:��!��ڌRCx�@"$��(��X5���W�����R�s�w��d���xj�|�aX՘G�2���4��Yҏ�cP��ϙ�o��K@�n�.���o��$ǖq�l��-����q��3��#��;��ˆ���	6��Z����d� �|���5�^� �KDm��+eV�� A\�7Q�$�=Tz��������捚���^m����=G���ͣ�9�;����+�2������Ig,5$?�>������!;�S�f0�W�����7��˱z�{�[o��`�������y&OMqPK�V�7� \��	�i�`րX�̙�|U4N�:�*�܃�8j�d��B��T��5	�X�w�Ӭ*��Y�����}�����v'�smNi�����=Qj��ڿz[!���lW�q:IfJ_}��؏0�%�zS��TH���?{S�J�<���'e�����m1P�M���/V��qV?#K3LJ;6^9щ`�<ֶp`��Eֿ^��\�e�}���
�B��J��H`D�Z��1-:���4h�158��S&��v)HP|,�__�^��ɨ�-���)\�����{.�yi�K�!u�;K�D:x0��N��v��:_0Xl��6�D؏VBn�V�@��H��A��`����PO�P��jީ����u1��y��3����o�4E�ꏒ_�ЦZ3�vT_���8��+[X���D}ˑ���7�W���WY��?�A�����^�5����[�TC�A��ܖ�G�������o�a,��5� UNE's?�L Ŧ۳~�t�^� �7'-Αm'� .(*��M`)m�0�(B���!��	��~��(ʟ�[�Tm?p���� S���Ϟ����TLrN���V[��Y���ca���<�Ҵ)<�v�g��5�����&hz5�o����wß�\�p�����{�b�dFHA#�kjC1�ӶY:ŏⓑ)�;�ЪѦ�d�Rs�\����	�a�`��F���MNX𞵅8��[^1�n����+{=�q�,���w��R��čF�t|�z���_��]���W���!��=_���yqO��_D,2m���Uǩ�9�٦}#-X����	g������=�lR��Y?p�(ihAO�/�N�c��B�5rY��<����:P/�b���N�]sN���G����>�Edxv,
p��.G'mUԂ�B(��u���lB�ɟ�H����F�-��ċʿ+K��81�C�z����ԳK������M��^5 �w�X��UR~ i�b���`R� ��y�s̼��均f��ל� �`^�ī�CB�
%}��b�
n�ڰ�1
r Á)�����S��>4�Q���?�0����d]��-�jI�G�;��O}�l�0�u%�2硍�<U�>���>� �����{���xXd*n,lÐsC|��,�Lۼ�T���f��y_B6�����f$�^�+��Q��r<A$a9�0�[|�Į��~�{�os���	pRhBG�OwYw�ܒ���g-ifN�
N���݄�q�e_�EČ,z�Au�O�"'h���Ty�`�U�����>��ȵ豿=�؈�l���a�l1+pF(�5}�)�/��k��'�/թǸ�Nɳp�!K��ڢ���v4qx{S�	6}����)'��fV}��p�9��e$�=�))����<B�O��ȝq�(ZkXf��x�I�24w� wî���Ȁo�ޠ�$"-�/�c�Cp!�~%�tzb܂L\�O$��)�4�8tH����D���$��0��{r0.W��酕�pY�?8V:ְm�Ƒ9�Le�o���K�>�N.̴~�5����v�aM�K�x��W��.�5~�Z��HY��p*Z)tO��g�!;�Fׯ*a���J�$�\����@Ǘ���&]�`��FK�z�t-%(�B{�@�|���~�9|,N&�IC�~�+}sV?&e1�|�	~��Pg[y�ta�\SyIwX8:*�,���X�1����j���dūaOd�*��M4yzVTڰ�=�.J�뻀?��uKуS.��I.�T��^!�nh�@�L�L9�z�����pI��T9xb��@���G�4���umL 3�Χ\z���ά�Wn�6��M��t���� ��@ͪ!�{$�SΫNcFt����}�Wd"R���{=���b-]�=�`"ۉv���,"��2T_Ɛ��(�)��
����y�����+�3��ަ0��[q{�����jJ����G�ў)L���`YH��w�7�o�a�a�Bt!ІUt�=  ����!fدus#�&��!f�����U-!�?dv����(�_E��<�&d�bP���^�WYF�hՑ�|�A�Ñ��=��??6����yN����Ј�� ��+K˯�98e�j���ȋ}0z��}2�����=Լ^}�:���6�,���)�U��k�ʰa�V`�w𥬆��	/����kσ�[�o�ө�b��w�^^�
�� ��f�D��a��M�������q;��/�	�W��<���<�dK?fڅ.q+�Œ�g�����g��؞�w�/�ރ���'r�N���D�&�nx�n?t�3��l�\��ãr�=2���מeY���[Y�O�<:=���g���7*�; jm�cd\}��b������M	f�,�/�O���;��O4��F��4;d�ZG��gr�G��@���'�Z�M2�ƦV  4���QŅ��+�S|bs5$t�[�N!o0�[���
�Se~��f���`��QP�-|���!�Գ��{��8m*q!�{�G�)�3Q#p���=O"`,�H3 �+��*��3�C���֤�>�z���8����ȷ��)�*�u�j��qq��iv^����H��3K�0DO��5��ȣ ��y��awN��^� �������cM�oR2�3�,�,���^H��I۷��������K�Ϗ3���F��C�:a$�7J%�x���I��<}��'�H ��C�77r`����S���~LHkG�����d7�e�g�V�����]��� ��|��G��X�צ6����J#J�ePn�g���o�q�^	��0�x��Ҧ[�8$�G�sh�N���+�My���*S��d��+��݅=����?�5\�x6\��1[�1.޴�eZ��N�����XZ��D��e�;�����ׯ�7�10 ȰcQS'�3�G�E���(�'X�N=�.�j�����e�z���̈́Oy�@�@/�q0�=7OkD�e𤋮�zn,/%
�o�`sLݎ�a���gE�NAb*PV�(;S�ޑSPcA�	�&j���+�)Q��!UuS7�j�.U��A�1r��9�A��� ���oE�� �`"3�+���_����7�L����d�L�	�4��}fvr����듄�,�k4j����昗�ܑv%`-��oSCa��M�v���a�u�;�}��v��?�w�7^;�Y#F���̔��k��;�-8e����|��:������	��F�*�\�u�􉮿�wFހ�R;;�"Q���F�R���n����p� K������xj��^�r����!�ٹ3��֬�m��ϭQ��hQ�'H���k�x�u#U=��,�S�*qS����dC���,�f�M+z/�T�Y��a����j��+}h�����1�*����_��ŝ)h>�[��5<��~�����W�%>���Nn	d�Ur����i�펻��m���w/=8�)��&5��)!�:��ա71dˑ���>�.f�'��^�'\�i�\��]F٩���$�
����K�R�u[&;72�;���n��/�TG�_I�����PYa��lW���� �+�S�D7P̋8�=��;@�q�����7�Q��������	�=��; <X� (�V7X�	���<�X0��(F6�pzp|�.:-�����sL�aθ͗�m���Z�x�&�������w�&����]I1>��շ�<d
F���^��Ac\R�]tp�9R�
	Y�(Y�.݅w�b�7ev�ƪ�9gm�:��z8P����j<�ΌnG���X�����@ِ�(3')�x��rOę��G��9��N#���b~�"��pI|�(0I׫v0T"$~�敉k����)~A:� ��H��|C*��Њ:'w����\Oa�����cT��N��a�*q{��ORA�ci7�#j����K�݋�!����2̜}@�h�}����^�ag,�$P��,�`͇�b�՗)Wxyj9��pV�8��l?��iӖޢ�)���쐪jS�/���@���R�\��(�aɚ��	p�_�1)�ݲ�f�� .��"��)3�S�9UW�"3��~]�]�d�SJQ�'x�p��ӯ��4c*Ȭ_���woe�s�1|S�r�Y<$pr�6�ð�UDuб�%���7�I��>��o�)�-��9�M�L�h��qp&O���k
���!�%m�֚��gB�=�/f�e$f��Ū�a������S��/u�M��d{:p��EϮ6kW3L�wpN���Z�K��.������\�t��ު�����*�{��)��6��8�6S��u�o
�#�Z������\��l�Oo�@9� j�EL��b��|�5�1Q��oXݣ��s^�~��9-��ɕ	��ƣ�}�7��/i_��t<���ن��qKv��9�v<#�M.0�h���~
���s$�Xh�̿Ὡ^��z7�O�Q#�ǚ��/���S=�x�=����Ǧ�KKڠ�zt���5n٢6�1w|����2}�yO�1�HG�����޸䱹�!��ZH[D�s�Sd��V.ݒ��p�{)�j;,����ԕ�`y�e;�p�2���b=3Ϛ��{T�lH�'؎��K/и\��wfD�Y���/����qA~24�Q8��Bݗ�M-K�d$��ϧ��)��`Du7騰��k:֛�Ǭ��;kP���.zt���E�P���!�m�ܭy��"�I&����p'�m?�1������z�f��ܦw���Z�����^���mbJ��L�}+:'��%���XS^"�v�"(Kc�QAa�(���Aً�����,�Vx������Y����9#�$/�o����f9R`kLћ�k��
$�z�k�G�U2�&��/��!{�؝��{ԧa�`���ET���y�g����j��!?���z�h��E{e<'9ҁ
r(`EB�h��Ө}�����<�FS�{Re�T���г�$,L��|TY�с?N�'.Q�ÃW�H5�}Z�wi�@����F|�uOC��_��oqmA������64�\�\����H��D�m>wܤ/�7L��[��f�a��r��j�L��+�p�8!c�9F)`!�^�?8�cU����!׌5&�L��������W�
�5���cUD7�Va
	xj���>�*g���
c����~�B�S��x��ؕ�3u��~'�����rw���s��[a˾½����ϲ%�T[
�U�����BOu���H�*i�W�*�rsxǰ�Tb���ѵ��Joh��_~�5�-h�!v`�*V�+MZ�c��{�5�Wz2�X|��M)$�Ā&�C#��G��h�±>JN�]��H�M����>:fW��� ���/��vbc^���3]n�Ny֋�*������?;�6������/��Z��`b�B �p��������V�c�@�>��ė"?��&���7$�YW�of��3�gyŌڊ.*@� ��m��u��X1Ƕ��P	��O�B���
g��r�l�y;cM�hz?�����7^��'x�P�����-Ѧ(�*�~�s�q�GS����M��s�q ������Q�&Z�jiu�r-=�>��ʒx���T���iX�߈�_Ϩ�9c5����@�+� ��K�ˑ���z��i���JY��jP�d�㼻O
<-�FHl�B��	$��c`{��?,���UQ킀rO�HI�
���IkWH�dܱ������D�8X���h���� ��:��j�VF�N�x!~�J�0>�a��Tĕ����\�;L��%��탏�̓�II�Tr�]H+^{#UGT���3�N�_2��_O8 �mw��S.<z��6��bxh�o�
Xܷ�4Z�ύ;����?p�~I��a��*/�H.�Rr����g7�#u��vA����b�������~�����d�f��M*Qe4���Q6�׷�*/x��4�B{ᑋ�6��-���_u�@��Ġ��{�m��
K>�TI��Mu�I��P&�fJ���#��V��a�
)f�#J� A�����\����+F���mt����j��g{���{O�]������<B���nQ�`s�P1��Py�~鯓�U��n,��Q�;� n�R�f��cr4ޥ�����Q�'��g������bgZ�5�2���7��QGk�]����$�0f�#��z]&Q���B5�de�=�q�S2���)uL(%��2�Jß/ ��KBA�+�rg ��`�����4(d�ym���E����	�բ���E�
Te�s<ގ��+%j>�{���>����%K���v�S=O��j�t���̠�n�cʦ��ǚi�?�����Ec'��o7ݤ�3~c$��ݞ�?�A��R�sbD^]@Ș�7�W��e���ݚ��b�nP F��7~�M����<z� ��y�;�S ��t�uRs(�X�S���M5�`�©��.�nZ-�O�0�T���r��Ղ�U���}��p6K� ��;�8��,t��!�®_�4(Ӊi4Y�/���,�L�:[ݤ��j���iq�K��!:��g����<¾#�p�6Ssb��5�r��a@�._kVd�V������2ūS��e�n��z0ҵ���X��˂Aul�����<��3��>�)C�-�d�M(�[|���m�!n��z<>W{@��p��0�H�O��PU2h��4q-����I��S�^y�µD0X�ל?�A�H�S*�` 9������vP�1D>F`����SX��x�0NQ�1X��ka3�)(�ɋ��w��pOw��}\BC1�l��.�- h��䦥P�Wb�`�V�	YV��.�	[(��'C}��w��ѼR9��-2�Q��U����O&��Y�oמ-�t���A�eH��S'af�Ud�9:����b����[��Y�;_g@�ԑH�P�,"�#����1z���+ Be���e�w��<+�UJ��|�B�����r����������pN��B�:�hc,�
�ы9:�����~q{�{�3?� ��� ���Z �h'Od;�NFT���Qjbq�u��fH�`��-�p�������L��U�