��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\���V�fnvx��ÍG_;�ȅe�~�>���9�>��Y;�0G��:\���k_��g�V^ԃ��K��9}�}%`��d�lB^jqc��Ű�k�܍llv��ԹP�u�fNgP�;����p��[j�2��9�$�sZ@��AI�olN�K����/YK������ �{a��!�s���Z#�E����r�tu]W�<@C��:$��_��G�N��)�!^��/�:E�)5���ܱ'X@�	�3U�a�3�=�t H�%�)��� ��Ș�K�n�i�d�������5%L�� ��:A֋L��k�5P�����x"u�Gg;&���34��o�(/��R�.c_�n\{2�u�s`�z9(}S0q�V���:�r+u�1�H?ڿ� -����h�h1W��K�	�&)�ѧA�l���3�!R�'�!,!nx��\�+u{�$�d6�x���4�aw�L-d�A�b�me�Q�E�K�1�����HHB��'?V=�F��ܿ��f�#z��N.wq����gņ���&3Ww���f)8�� ��Y0�OY�c�F�=^Z�^�:%�,4@�"A]�1Ϯ�}��=��d���TW���`��q��~���� M��s���t"m�/^6ù7&�\1��)�c�W/�
�=g�zO�]�(�׶ɝwMm���L�^Ӫ�3��j�j��ˆe��@N;�h�����-[S�{٤��5����`���N���J��`/�˞�ʠ��;�0�4�uE��P�2����p�7x{@��o�����8L�3٠���k;���`����υ�;�I�����U�НeTð憈�Q4&�)O$�-�Ka�� �ک��4JUw���,U{�H|݋8�"
��y,4|[��6]R�ƈ�@[f'��&�t<�~w���?�j6O�h��^�0�P�����b�@ڗ�=���@�+�c�E�4͎�ᵸ��~2C,]��C)vp�mJ>D%�|ǂ?�u��A32��n����Ί�;�[��L��5vj����5Z����=<,d��J&�qy�4��j�f��֜'^�^(Ǌ����r�z����#�#�φd[q��	�b8�1-��ᆷD����`�"�>���Ο���q*p�����l���k�'��J *��l-�o��5�9ll�S�S�<6��ϩ	����	�7����NN��촫������O�opl�")�5(�l��Y淥Μzzr��z`��cuotpc)�o�\���m�ؘ;ե�[����Mb�5J�S:$J��hr�=�6C#����M0a
s�0�1��r�0�4�K3�u�gX �y�u�S.O~n�4�n���p�@��F����`l�DM4���/Nz�'"R�xL1˷jkf�+'�ֹޫ��1��Y@U���\���v�.���,:�h���E?n�6
��U�ҕB�u��q0^�9Q�� �p@�D�ُ�I�&��YQ�NCH|����
[s��&OZW*mB�p>�9T���W[d2�ז���Q����e,�~k&�
B���_pT�Yn�`7<=x���/�>�)��rʩ`5ؚ��o�|��?��P�����%0��ĭ�Y긗��(�4%2�#? r��O彤���2���ԉ���_��Ԃ�.��(" �I�_�@�����t|D�SHt-�ˀA5�n�V,򏸅��&+P�J���4����Ȍ���4�Q'k�d���3TE�T��iP��(J�*9�|UI,�d0L���4P����z;K@0J�uNm�&�m]5���%�'YN zw����5y��������Š�%�]�F��,O�<�Z���r1t���&��Wi K��r	��%c>0��pN�bX�S�o��8����Q)�;�E'w}R����5C�AV�� ����>&�r�w�Є��@E��oPf�L�k)��Q�����*��l%&F痻���q����P��}�i^�`y�T�3�	_=����}?���͆��EL�ú��&9_a;s�H,���q���<D$��v��to{�q3,��rx{�����5�L�/�I5@ԓ�	%Q��M��Y���o��H)��ۅU�0{�{�R���K����g�#K(ժڈ�?5?U�Z0�ݔ���m?�M���i�w��0��_pֽgpOA��# ��y��PR]�S�Y�*B�{���P�m2�\w������	��Ё�ќ{��Ԋ��X?Y�*'�w�������
� ��8t��8�37�B���A�\���>hC�\ D$��D���tFT��o,��[eC��{1<{�Hu�AsQ`Z$�.X�"�}tKb��D�7�c��I�\$Y+�߈Z#�M�М���Y>��q��9%HN�3q���m��*��XPr�l��w_\r�/�dRf3�%�&��?}�l%��KP���.F�u$��ֈݫۋo*���=����6T�e�u��:�$�g�Cm��~�!0h��^}��x����tw�\(�Ԇ��po/�f�y��9�����z��&Y���<�>�"�>jQ/A�ڙR�&�WN�K�;�R7���*r�X̎>q
R��@�'��~������+�W?+b�-w�ܐ����M���{�lw��$�aW�|3�G��f5��vge�ybf����v㿥{��cA� �ǋփ��ը�-�!R`2�
��T�Q�F�()��4V�q�p���v���iF��蟰��?����㣦\{|�E��`��1@^ t�����-F2��-L�K���Q�8����apt��Q��д�q�w!	J�_V�5W.|�Y�ZC�ك����/~\���z�bw�B�c��U����3_��|ژ1�/7`����<KB����^�Z�~�����z���Z4H���Mg�K(WCwVk�/cz�3�ځH#���wVss"",G������up9�����~�_-`��K�5uPg@����l�<�S�1H$i72R[mƸ�]�/�P�k��D��SԅL��lH�t8ĹϘpY�糬����Uy��QS�nȒTsJ�Fe;?c�S2�Āyj�����9�T��"e�hBp�V6�w C�G;���*�����>z��=y�@1㰡���kV�A��[�\���h5�ZI'�����u��x��z��'���0u0���O��*tݙC�qpT�ս�19���EJ$�P�㡳�c�#z:�٩�����7M!�3�;���J�XB��Eq0�5�.�XӚ�����1��iC��� -��/��E
aR	����!Z̓�e�3�qLpZ���+�sW�:0�
{	2O�9�[�@��Ũ�HdO�H�"�1��g�L�� .>�X�)'y9(�
�w�7|�a�����b��$œ �%��)w�"/O�M$�ɛh�X��3cS���<�5��t�ٲ����6������z$��wT !���l�a?r�ʾ a��_�s��aPj���7k@<^���6	v�j��@��Pw@L<f�8����^��&g�#����$E|�vJ������7;�
�������U#��l\��=mp�&(MF�F	f��T�8�<�s�(�t�����46�g�0QCC���["�U��ݫ��Z$�;Z�q�����$����JYd�q���l/D�!�\�TO�0�����[�)^/}B������#JD�$����ٜ��很=�f<e����!F��c�A�I����s����&�l}|s�Fis�MN$�'|��uc�&�P�.�u�u�3r1hA1� TPG�1�e����R���;�o�ͦ��X������vgܗ/O��RIg�L�=B��` Pw��&Tv`��Q�-4��`�9�����;b�#�R��U((h�-5­{�G�P�ª&��#��1[P�2�GY��E>����PÎ%��û8a�gJ@����G���f1܎�����f\���(�ېf~���S�6D�h#5	�^C��P5�;Ձ�7�6�k��O�2��&�s�.l�T���|�J��>j:;I�)�a��6��X��^k�����j��1�'?�f�����,E�;��_?�h7�ZR@����0��I�4����Q暳�h$#�7J)��i�Q�ŀ��)wB7���|�,c��b��A/a�KW6�澐!�4!�1������|��v�]�}ݏaW��<�$�V�{�0���F"탊�J�i�[�9�s ��+]�	�d	zC�����S��b��!�5.ܤY�_�e7�s�P�-