��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\���V�fnvx��ÍG_;�ȅe�~�>���9�>��Y;�0G8є]]��1=z� �J�3Mi��	8\��FM��k�sy'��j`�o�CD��&P�:J�Q �/f�7ĐkA�L0\�����\�n�՛�Wb���Fq<��:��� �\��C�#�RN��dGf��)�4ga�&���6b��zgH�y��Deg���Z�ɢ�d��s����n_���2s�Ѻ�wy��&V}t�e��l�q_U܎�_�.��PO�[s�ΚҰ�5ч������[���S���3ݎ� 0���~��8 F?�M���h$'\ԝmE�\�Gz�z���Y[�U��Z�6-�f���,Ch9YN�Uﱤ��!�R�
�14��Lyt#��ie�������S`�\��X6"Z6��3L>�?~q����z��{�Ş	]�k��s C�4�'��)/�N!��H�[Z��� }g<�
K^�Se��o����ca]�+�È�b}R-?:T%�u0C�����0�	w0��*�'s�R�Hß8˜#��ቮ�l�����]�-��s���� ���,Ox����)��4"�|X��HA�x�Xl����MUYƹ�cdd$@SBv�yE���OD2e)�G��<R��;
$�����0�i�D��a�*1�5��~�H>�2%�ٵz����(JJ'��}�7j��Sw
�r�x&X���M&�U�f��=��5^[_MߙI����<	��.�ͽ�-)sQԞ�-J��Gg���?)�	���r��>��6*��sI��s·{*��З��@�Ǜ���[���oL-#[{��7�
޸�{��C!h��դ���۪�EQ;r恆`�k����
�!�s6�EB�۬h�#�8�a��5�n|��2���,̚i��Խ2 Vk�{�f��~�ߙz��Fu���B\H��.�2<O���Q��������
$�{a�J�L��&�CKNs�t����l
�Ov��!��lO�]���w/�ގ��T8C/&����P	�%��"���MJ}E��T����6��1U��Ԯd��������,vnY �qm����H��2�!���~.<ޖ"�)��\"�z����h��-��{~��k"��~�3V���5���5�>�Cw��,�#>��ї�)�
�0+��%U �bY����f�m޸f��-�Ո6�H`J̥�I�&��X(�o�ZMP��Fd��1�z	�FUQ�J���X����n�&:-�n0|/ِ
 �q9g��<3I�)0�z��rw����4��'w�jv�֏�p����^��1\�m&X\�%b�w��K�)�f ;c�>s����DK��M�6������Ӄ��s{�2�O�G��8z�2#�0���vHS(0` r*�H�5G�Z���v�5q�I����=�s#�H�����HKi��m�i���"�.��^Z���Y���#?*CS&z�#�h&miVm��>���@�a��Z�ٳR>-�����s|~�R[����k5<����{�c����e��	��R�\ ��"*L#������Wx΃6ꏷ���Z=
�p ���W�vD\���@S�/�I�/,�?q:`Xb\��)�r%E�ު���gB:lr�tX#[�P	��Ͻ"8Z�Kiz�˘�s���R%[��f������;��cCy]1dF��Fto��v�>�O\����DD���7�ݦᥤrc���W�����c�J{Ӏ�*�<�/��u'r�f�������Td�)I��?h���� p��h��d/��Ll]�j�˸�t  ���lgL�h�g��0��6[�����ʋ 6Y\��h�p�F��%tP���ްe�U�߯	�n d}ʼk�~���{T�g�tj���Yn�>�z��`=�
Sт��+�Y�&�VL�nL]��e@�g�Q�{)Q\�l,m�.ο5��f��������f�՛��y��,���+�m��<6��Txj��2��}8��r�Ik����\������\����X���\34���I��"�re��_݃��
�lY��h~���o�Xz1���#Q6�إ�=:A�p�y�,���ͅ�f���m3m
� �0 ����O���E� XA��ʋh�ff8$��d�8/�a(�(���4`N?�D
�%m*�T{�b"E
���8�q
�Hvt{,�Ck���h��:�9�9�V��Ud������S�~(���՛q-����-ya�M�m����ӯ��<e�c
E,O�V1��F��s.�Tǆ���YR:�����ȟ1Q����w�ˣ`l2���BG^�2�8f<�\�f�+�d"��5��y��3%g��}��a>�����ct�u�hr�������F��:amcމW��-��ȩ��f|�W�˸�NsaL�0̲e=��/��(��aǆ�WkKص��N���|繄���B���I��+6-n��%��mZd��8L�P��(#���Q���Mf&�Z��z>B���D�����4�M�/&MCV��H�?�]�o�d��Tʳ��9�חT�����Q�?e{f�d�ji�3�z$�CM��,�R5d"�
<=�kɣ�����nO��[�Bcr��/�)OX9��n��t������͂r$��Wu$�E��	����]:D�1�@3�A��<Q)P ��msq���s�bR�ћ��N۽����$d�S
�/� K�5#\|��oK�>��i+���ЬHY�����\����br�F-�1��әp���O��"l�mYN>Px���;�:�|:BV����?5�jn���3mR���"������֌U���IE�A��;W�]��z����ї�eE�KӉ��l�����L�[U����%d���Z6�9��-}� �E��2�0�c!'K�o��O�i���1��M��.U�W��7�����y>O����m�$VZ���o����EX�G��(��Ӥ|q���_د�����EV���ę���9�dBuj���Y��J+��C摨�\��`��I�-�Ә��qʒ�h�i�@�4'���[��3�q���+��x%���K����6L��w�!���3u��ᇔ��Y��y/�rql��[��1�F�?��f��4�Ҧ�_6�5���g���je� �
Ʈ�k��&��z��y����/7~���|rh�S�C"�[�ju�4�]�W���jۚû�����~��hi��o�qY[N�4��N����"�p�FJ%�����~g�\����>&��aE�(D�Ş�5j�@�����c�IP�a�i�������*o`���������B��]L=
{�����眕��nN�7�w������[�@��N:�fY�d������4�$�$A;G0g��+���`���W@�Z¦d��F܊��;�(�[�/�.�>h�2]d7��Q�$ ~�c���{���J�|쿎 ��8&��S̀��B`����o4G��v�N���=��yq��L4;˴��t����:X]	aW��7b{�)�P����sb� 3�'�;�Fù���^������,̀X$V9w~t0��G�0(s�94ɑ8,��FU���B0��ܪ�Ӳ&n=މ՞w�D�ǈH�:�~~In��Q�3L�(�E���o�l.0u�MT��NnQE ��xəT�#ǰ��,7a�����Ho���h4�-�8Eϼ<����)�!�%��5q�B�u��N��ޠOX)�'���[Dd���)�?9��+S�֟t�x ?�{%!ԕq��"#Me���;_@ h����,�γN��o~�0V��Rۓ;���yNV6��1DO��k��
-`��c�@2�O��9.|�8.க�\3R��c+��7���ST����?�1��4�Y�ij�ҙ��Uiz?�ϣ}��U�*9�|�L`���VI�#�h=oJý`p���G���8flAӋ�jD4�w;[���d�*�p��j��W�'$�]����D�'[��V�0 �S��|�]sh���D�7/m#Ε�rjQV]n��Z�9\ܲ-)��ʏ���[0.Е����*��S3���B5�U�ʰ�P �u��v��s�%�2�c��7f��q����g|��M����kNV���&�[�s��(�X�e��TK2,#E?
}.3�C
�r|WL����N�ִ[u��C�gk�aUq8�Ҋġ��y+�D��[�&��}�7��Oc""�=zqďx7���<=��X���&���6����tzř�JV�X���v6=	نc���z<G�<k�	ug@�υ�lN@ocF<^��/)fJ�"�|>��O�7J|H-��UȰT�6"Z ���/��k���o�MM�cp	��)r�wRXt��0�X?%�)����~��
�,��9�F�����H����M|7�QJk�լF��1yj���ۿ|p� Q�O�:�{��h�$Iْ���D%�]
�y������
��L�YP��4.���YB�"
�ͨ^�z-�Hm�\|Н���;�OUs1�g��ekG�B�ފ�M}2�S���IDID���]���~f�R����p�������#��xzx���?�b��ʭ�Q��7��N�Ʒ=���[b�����s��eb�k�qDt�Ƚ����r��%O�FH����K(X�o묃)-�HS^~g�s�,�m�#�y�����[;�����Jt�ӽqQX�o�7�4U�p�o۔�|K%�`��/�k|��e<�!5���+��M�с����DBH�u��(��D+cC�����.���I´��W*��7fHCy����~Ӿ�:��\,_@�q(����i�-�5Ǳ�έ���S�nd �޲y2g%��ҩ������$[�?=wwl�蟮��n���8ȭ�f�;xnrT��}�#i��b�5R�y%S��Ð��[�t��C�ڿ��j-��K2;bYdۋR���"���x�7�(|w-��@�5��?C��#w]*�#qTF�`ʊ�~1%�.}�p���\;�K�Cz�J�,H~�T)���S��_r�Đ��XQ9�(r��ٰ� WX��7�P1/���B�i>S$V��ˊ��W7%s���e��{��"��}��(�W5n�{�����t�$Q�	˙GZ1�ι�}H|�ű,���ڑ=���_�j�%w��vO�a���y�IV��lW����_<�<��#�oEF�9�?�׭ �\ P����c|)qw�V�
�:��X����h���bSNM2�����x�l��nRd�̔^�z$^��A\ʁ��(�ճ��2�)��&o��������K�a�/^y"v�{gq��a#�[�[�ꈃ�������@�E�%�:����Cs��Dѣ�>2�^�|�5p��ڊ�۪��Aȹ�)���iHa��2 �>W&r4��#V'B�{�,�)����o.8�G�7
�>�.]3��c�J�q�����/���ʇ9�������;��'�ƭ�n�ɼ�&�X'�}B��):7>���񗋲N6�?pT��T1�On�K�}��v7�=�^�4V�jG)>�6�
�l���.w^��*��4%q�{a��"~:�	�S�&i�;z���(�[������ˈ�:&�C+���Z��l����~�ck} �|��2X�TQa�	G�>��E�l�s��^=�ph=�O�e�,���
,��,C|)+��^`���K�����3UC:␖>�F�a]b Z�,.Jn�[�oD5Г���8��|�;�'����2B�����KTx��	���"4���0֟�UL1����{wT��<My|�n�6_����3�tM@d:�0#�}Y�DԿ�o����JO��� �u)$Ҽ�>�������'�A�;˴�d�a���$H5m�[v�ܱ�N��j����-�O,�!^��ϩ��~��t�J	�Ǯ�UW'_���M���k%2�f�!}��	�ds��M�[�=�c�\msbyMB���Q��ͪl�9�a���6f�<^6V?*�%"ɾ�[��ݟ�Uep�(=RS