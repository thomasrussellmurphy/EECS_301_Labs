��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|n�\&������Y��𗲒�*z|`C������X�:��^�c
J�����'�Z���*��a7ݍ<ZV�aiˇqV g�I���V]7�����1�Ա�o�o�ʓ�=��j�'���#A��4*?R(��-�UcikL�� _��t�G�&�%vT0��5���ⓒ�!aj	�|�Ѩ�����}���('���J}�I��$�_�����eJY<&�b	�zO�}&��y.�<�*&7���|>�O�ao(;_��؍^f�� MƉ�����z�_@pS�(��>W�fk�ݟ�-ŧ���dC��.n-��nAo��b�,���f�dW�է��ol�a�vj Gg輰uXd���}V]n�;,O��T�4�/n��"���.�}>H�y�8E�J0��7���#�-�q6�\+�L�.ӓ�HDh�h�eB֤z?5�ʞq~�\ �������5<����)^p�'wE3a����gI�t���LCx�\*�x�Ϭdr�r�>6y�����vzH32�N^Ѥ�Ͻd�]��!WvrIx`c	���4����KXTm[�j]�VK����$���j8��̔5���	sq��]Y��H�;k箰 %I���W\FӢ��� ��5��5L\��U��!�e�m�s��i/4���@ ���
�g��^tV�	cE�&��V�΁ �o�)���^Јo~���"��8�&4�.5���@�arJ�ͪ�W}ҁwG}5eMH�Rq���բ&S��k��/
�$!�}  	��&Z&m�gۜ�!Bm�.(ND!��t�3�pT��̕Z����*5Wv�
�K�O�^c鍭���\[�y����CծEm7�֡�"�U}���L�Y���IF��B�rMu�[���
,>=�f�J���d��nd���e
�ޡG��v���#<4�<2��|х������>�fAǫ�1�0��N�d�Zdrc�󤥿N��ǂ��0#���xƹ}���x�u��pn�Y3B��?7(�\f?�!�-'FDY8�Vn�7����c�hр�K|�����q�^@�nA�7ja8��́,���(=X�:�&kT/EQ�̠�����3&����!r�4�"�wm�,� \�Ի==aBn��(��?@Cf�H�W��3���RL>�{���r{ɥg�|���>F�<n�"�2M�!�;�����%狞]#W2�ٜF������k�S;3V��N�V��Y����dj��'�]�^��j��۽P�)�N#��q�F�� \_�7��[�\�.�8$�7wf�>���d�gh��� d|9)	~0_�n�%8U��6�#�p`V�"�,��7HF���X��l6W�� P9yn��\{��^4�u��L�}:�{�'�s��UuE��֤�á"<[9�銗�V���U�r>�ζ�,��h9���9MO��T��d�vFytt3V"�`Ai���*4�@45�n�3CG��TY���oՈ�y+��B)kWX�(m�u�Nr�����V��v�����3c���	�R����ܪ�S�~`ō6H>�����J�8b/zr�6x�3㯮��qz��������Z�0���Ѕ�g����T{����Z�"�������~��-��Ө_tC� N���r�5Nġ�̄En/��Dd1s������J�{Q�$�����}�{5l[m����QsD�~_�w��t�}TR�_4��@-B��{I
)P3j%14dk�+k��M���e��d���Mm?_�Eyz 0hUUw�Y��d���Q0�Q���s&���(�Pj7�X�ǀѲK ����U��[��}�/�Ja�2��}qJ�5�����,i��hi�o��Y�-����̗:�c4�|K�g��#��GDS�B��d6��@���tx�=�4���_���J�2O�6?f6���\N0qfc{�`C�OeF��O��Cl���mw��a���#
�iD����-�:<�����ΞWO���NWH�d%:�U�'h`��8�||�6�do�t�v��O�Ɠ�e�T��E�]3�b��bvF[�S��ͼ��7�j��y(V%4xXDވ���թ~���ց�)���
{��}h����A!��Dh�8��Cn�u͵�W��\�^�M�#��ē�ge=Fs�L��QŎԖE߉��9�����PZ���,�m3�1�-0m�3�W}W찵q�.�@T\eH�8��@�9y^��w��Us�-UM;'�Z�fv5U���M'ו6E=�vo:{�j+�e�$��f�B����p]qµ��1ILLB;?{��z���1�C輦��~�/���ؾ<v�;��S�e�/�� ���Ơ<"�z��.E�ph���j�������ue�z:�N�GP�2?k%I�U��Ww������)*����mC��(���KӦק�̶�1�6kΕwퟩ��+�X����j3�I9G��0>��{��s~o6���:yx�Y�k�D򊟗K(淑֕��������¤J��«4�Vi�}�1�� ��U�mm¸Iy<u�$|!j�fR�y�8�vL�q
_4�2	�I6���T_����=���Ln�u�ic{��6(3���Ci��L���j}�s�;ll��nבL2���d���a��O}���;�q.O�1T�s�b���������wx��ƚX�?(
Ȩf��TB+X����Fˮ�rU��z�p�6$�
=�Cx��N���m��C3�E��w����{��vtcE��[>?f�N"X�G�}���@9����)Ĺ�܏1Ll��fi�QTҒ����<�
"|쬙U�%Qo*Z�q~.�<g���k�dե���I"����n�$m:���'d�~��L#Rx�`��u+*�D�`0ۂ�;�-7?�p��A>����X ���S�b4�8`UɋU�� �TI#(G��DG�_���LF��%Aa�4z�McZ���Z7�͵�ډ�����
��; �Y��׊>���1�z��r��
s}�S�_�!�L�|ҒS�^)�7Y>���5f)��S��l�l��� ��3|Y�<�\l3�l��#��H�=_���X�2�^����:ݨˏ�k̶�������ݑ�Ή�_���������
��nL�|Čq�qBD����D���j�~�+�����KC`�]��%��������.�Ԏ����1�35#���F�w��}��v.R�M-�P�J�#��-��z��v?��	Hd#��;)�pN�����,DC-6ݛ�<n��� `�^�	4��>Ӭ���d�x�X<�p��{�� � ���P �A��RۨK5�G���a�n�W�J$\���� զ����S<Q�
����0ܳ�
��h����Q"�з���|��zt��T{�R�ߔ�q1󸎜�!
z���I�̿���G��ǚ)c� �;��XZ?K��\d(�ӹ�RDOS�h_�$�N,�I�m��ԣ���5��FY���e�Z/n����'B�_�e^b��%g����z�h�����T��}��?�j�U̅��j5Ml�<(�6�  8�P\���陗oڳB4��:S�L���m�.��At�:�x�R_-5Y�#P�.����Ή�[鈃���s�>�Op�/<ȍ���w���V%���p[�~P�ޢ�m�R}� ��e���S�bX�$Q���ue�}#�Bc y��yy���X��/�)1 v��,��6N���7�$̯6��� ���C��g/�t:.�� ��G%���n����r�#�,���AG,�f���y��]�~����5;	��z�̧����I?���6!H�����\�ۿ��2η曦o���W�e����ڤew�yq��a툲)
f:��<�.cԕ@���ԉ.�~�-�懆�'E�ϐ��Kc�����B�
�=��Ե֌KpM�)��Nb��Ũ?UȣK�5�m�H8Z�|�F��"�Ў��K�ɪ���T>� <K�Vj�<�o������n�ްN{��tR��.Z������2���x��];��.���7�i]���*��<�l�O����w�{W��=�%G�I�F�34��¿�VD�[`���)5��r�?n=�1����4��_�s:�O9{D2�&^1�"�9˱���;U3V��X[XD[jwp�c-����[��P��K��;��{�%SHV�����i=ƲR�9�Ni6F����@���<�gR%b�3�����t��6��Ԯ��ah�@\\�B�zx����@*�yxp����X;���E?B6���6�_/<�B�������Lh�U7g�pC��Ş07镐�xoD�lCkL 	!���h�}��3��&h>�T�uoy6_M���@0d���_�2K�J��ǰ #�4����]c(�gPDAD�Fv����B��W�P)����<�f�ZM� �df|PQ�sz���>����nt ڷ��j˝��Y���7�������^�VQ#i(Y$Ć�A:3$&���
x��Y��Lߺe��������^��U)��D�3�>������9���gگ�Q_t�?�������Q�B�[��ѫ��j�xwe�V�h��~+�ݽΤd���ʖ_��}�����w�٬N�La~�/l ׵��Օ&�k.�o��}���y�ܨ��.��>��{����s*�Y �n��ȳ]�b]���M��倻��-{�YG<�z�H֍�ߓh�c%���ɏ�Q����u��%�$?M�d�g��{�X$t��p��gQ���mZ�; &�}�8e�=��l�$��8���H������hA^�vb9Y��S���)��i�r�C���f~~�;Z����T�%Qot�ߏ	<�g�4\[VEfdE�[�� �٭���9��)p~a��[�1���g���
�%� 䮣ө=A�Ϳ?��=���u-ō�
#(	���&�OT��l�s�F9��o�����G���l��N+���C}E
�}��͎�D��JN{k�j�n �	k�2��둻��f���0'�q��	@/�M=������cR�oµ:��Nvh}�<9a���
dh$2C&���Qq���X�r��B+J�`{	�][��_��n	t?�7�a��Lw�%s.T���9˻��wX�v�o�`���2"���d��_5��~E�tJ�=H�g��-r�z�%��_����kk��%*���*��Hy�Q�eO,��Cz��:	�>*�P8M�~��}M�%�jO����a����gz&���z����	�n��F�W��>��c�T`�g�:_���������u~\@�Z]������V�ӀߞSo��_�@ �	�Rn.v=?��ӚI���H�d(iI����$ H����`.�$�Rt�$S�� �8�ٹ�c�sG���0Z��*�r��&��}NE4�d�@�v(��m8���]����X#{zW��r���[���L��1�h<b<�
*]˫7�:���6���ux�0��C�#+'谼�c��"ؼ�$	�=6��Ȥ���ވJ��JZ�;!$�&�*څw�o�ͥ�X��)��\�ZK	K�5 �g��=�c�옻�=C<Y��N�����}
 �?��@,a��nM���j�ʣ��JB%���<�s�h����f8�])R�`g�♫��b�[bc� ���g,�Z�Q�Į�����ӆ�:�*Ԧ�+���! �+�@&�{����O�Մ�oo��g������ a�����n^r�~_��h�$ǡr�n��	eG��*"1>{i8:`��I��N'lM�K�/�w�P��%���5�&�n{j�ji�%G��<��M,���n�QG �`�����Yd�	�x�6�S{&�=ϧ�0d�Ĩ����G�..��t�Gnì��2Ds�Nk�ٸ�O�r�J˞�|��}���I"f�5#q��hX% �.	5]��z�@V.(1x����L���.jH2�K��Wf}��_M�$�m�������t�F{	/#�m���ww���p��E�����O�Vʱ�Zb�#�r��H��<0#���ӳ "���*���1
�=,յ�'(�m�����^���V�,�O����|������(L�\y��º#V�(W5�X�uq�a�Fi�,�����,4�K~��)�������S����R�p������H��W.WC�����)Q>�{˅ț5`@��`�P�2N�쒗�������H�=J�aY���K�FК��i͊ �>�o$�%Q�ϗ a��C�CJUnD��9�X	�f��	"UvEA�(�D�ѡG�k��o- 1�I���H����JY��O>;�V������s��U.�:�P��[�!�Rd�>� �Ou��7��`KJv�����NP3!Je�Vd�w�-����s�l�u�C�@BL�X+�Fݤ��V�t��U=egߝ���)�g�.�;��t��Y��<>d�/�_3��"��GL 1��M9��t�(����>'�L΂"��k��UNbY���⪴�� d����L=�fTc|��?ٹ���	�0���3E�r����G�#r��`���k���;�¿����q7�G����t�~���4I��7�i�g��*�Q�B�[��|�\�m��O���~���G}}���$�����0,�(��[&�<}C���U6��s�bn,��<��R��! �̭���~ gݝ�e��XAy�'��P�/+8#��~3Hi�Y��-�"J���G��wp�qc�A͆������G8Vc��:�]�}q�(�7�413�O����>)�җ�R�2�sm������)B:Ԥ��hA��l�*�� ��?����nK��1_,����&��l5X3վÚ:KC*�mba����5��%T!�:�Ƹ4 ��\h|X;is��I?J��(@0ۗ&4w���;�t{�B�����F�.�<v-���|�PB/�:����;�����"�W!Rbc�� tl��G�r&��+p�0i�W��Ү�8����Y1eS+���5f�C Vi5V�"Ar-)��_���P��9W(V"��E>'�_������b�1�TF���}ӡ�h�"녻V�&/���ﾼ,�FЍ/��C΀�phdH���٬�n��U�πz\_V:A ��!�E0Ӥ�������(�p���}�������~[ã�.���
n�������J��7"�� T��K�v�LT�+�x}�!	�h�ny��,�8ϩ#+��W�|k8�A��'�hm��AM��K-x���Dk��:�8MG�o��&��Us���Iؓ �(zXu?Luj��&�$����CV��ԣ�m9�bl��w��!��\p�;�������k|{1��x��"�Q��.�8$�['���4�)rKY���;� �,���,��Ú#Rs�����_�߃�#�%A��Y�!��펝ݤF�� Bg@��X��6<z t��#KO2��k���3���N!hE����g�5D-c�o�G����6U�+�8`���΋�Q��J���8M��9OJ�P 1A�S��0c�#���\w�8���wl�m�&{-�N��Cus�F��v�t��f�OD�B�K��πG��C�'�E3�2�=�"(xW�Œ�o5�:�b�����!�X"����<=C0OkG���)A�vu����dJΠ5I���l��Ju�X.�����ͤ�S�'�15
�"�[c��u�[�X`�<v��(�.M�|!�����8�z����?�w9"�F��� S<ǻC���B��[
9E�?���W��c/^^}��O�p���y+Q����v���v
ҩ�w&m�A�l�u����|58d�wr���r,�5tk��qo;���M��F��$��췺 ��Wvf��#J?��fb�b��<�
��S��[��٪m�|\"2�䭵�@o-S�nS�{
c˩����O3�F;���bΟ�/���'� 50韨�FQtM�(SL1�r��PL�As=�IUK�>wkM����Ǒ�x#��x� \Q͂Ȍz�M�Mᷘc�m�x�-��sd���2��Ȣy�w��er,�aO�@�6�j�á���@�b�T_�
�}���CMaΆ�޻��4�w���4͞>@��X�-�,�Z�Z��&?@r5�*]��	��@,��܇���3و���ښ��#Í4�Xk)����\h�W����� NOB]�=�dE2?�v�2MžT#W����Bj��]7��N懰�sv()؞�?���?�g�z��v�or=���Sn�1z�$7N���ZI���ꙉ�����̯�v�1Z1��w�/����0'��^J���sΧ3:�ق� �֠���Q��U�<"h���u��$�b(fi��[%����<�mLZ��U�2s
H��������Y`>$	��w�ߴ�3Gy���d	T�L �7�r�0�O�r�I3L��*�:���Q�z�8؅�Y�Yc��ܶ����:<�?
1N��-lFr���ھ+���Y��KU��&�
\i�dl۬��.cF��u�J��ͺ{���΃T��䏂p�[��A}�I�[�p`ĳJ��n�==8�Q�$�Ɣ�yA$���"�4���u��ɼ��� R�P�؍�Ii�Gtw�Iz=w��$3�����.��h��征�������R���ڛǆ��Q�)�6�QR�Fi�rV�,*^8k�rԨ�ab��z���؅'��ZI�o�8��0�Kŝ�.�_&;?x2�Z� �{p�T�N��%��VE�>�O��B�a�9>���E���66�oǁ�L'?�F�i��+�U��iY<�yn�H#��M;��c'>7�u�|q�j�t64c�ç�<�?f�7���֯ræ"�Y��fm��<���.;���
prW��9e`:#��P�M�ElD�Nְ�a�a� ���Ϗ�dIt���};�M,=hdxܓTΠ��R���>9����-N�0�Mܓf&濾|�\r^�:�J��~U���)��������H�4������;���	@!cx�	nh&g��ԕ�<H�h���f��A��z �����k�R���D]z����X��`m� %�J��F"�R�`֍�tmVTWs_�1r_k�CS=�l���  ��,�!���N�
��Y�P��Xz�	S~��yKj�ğrH�(��ɻ>os��V��r<>�fl`u䳹3R	'��>�^�N������A#m.ua���&�YM4I�|;��C��KRM���\Q����]C� �TFD��
Cџ2W���kՓ�o�-W�$�剼��Q%J����&��2#�.+��������ٱ����OI��ޱbB�-����y:�?=�
_��'\r(�G�w�f��
���̶(�a���{�`�׆	[�3��@�q�B͖;���w6�/�߮a����M��jXސB�&de8�⌄�%J+`�gm?����Nv��%z\/	���JC�T=	��m�\�( :N�i�F5r��t*C��])6����נ���Hգ��ף|��5}1k�NT��g�e�]yjڲo�� 6���z���ET	��Nt�<@��W���>�"J�cR4�^X� �
�V�-�+��S������ñi�>�Q��\!HN�(�?
�W{�cD(v:�S�����Z#lmNP�1hb99Q8�y�.œd�z�S_GKg������@��\iݕŸ�sg"�[��ي����A3	~��z�IE"
�r��:��HbY���r���@�	88���tI�ӪK@$~3ٞf6{a7�dHD����yoZ�ơ���>cB.������%h�e���h�i��;o�a,�7�bQXXp�W����H��9ރ�6�QU�g+ծ9{�/�<�`��[nӋ�1Q���ԃY�6 �%E��[m�
qӷrw�{������ͪ�Y����q	m�����x;�v�}h1y�ÖT�'C��̚�1�._���}��_&	q&�k��i�s�@�.:m��|�S��'9W�G����[��@�v� �P5+G� ʯ2u��&���mOhRP �f4���L�;��`�-���VK[��g�W;c��h�I��S
Κ��:���uE^]��I"&�(��I��Z�³�+�f��� �����C�P�R�A���\c��i��k�ꏊ�U"4�H^i X��>�jR/q�õ���DO�8��e3G@��"l%����5�Df�%�)�>;H}�	KQ7T�~�7���q�����?��M���{��U	dQ��A��w��H�l��~��'�,�����)ì�O� ����jH�k(=9�m�Ϡ���%~H�tc��Mت���u�uN�����ch눊�K�F1��P���]\P��/� b�L�q��8��+��a;W�{$�Iѧ"u���e�/���;�F{e����8}g�<"�Ե�U@p��.�PZyѮ��a��~���q�[��]��b��1�=+͞&�pǂ��˄k��V,��Ֆ�v���Ym���cq~Gb9h<���_�#����9�S�QǁV̎Po���(���q�2�0��O��n�Э's03/)z��sǧ�`�#98wT� `����μhS����*��3@;O7�L��,"��J�g�EN?�u�QEc��&�JFXG`;J�ŅE�h{��vc�͖5Yd�n�Վ2I8�������f>^=���o�|�Iy�p��w:�KCX��{e�>(�����X?[����3�A�ұe���9���{���B,N�T�ģCe��Ѭ��0��"���Z1�KS�d��,-� ��,Nv�ĵ��g�
C���)�s���Y�-�R�^��T�\��7<������3�'�b��%'��7a��S6U�S�|"���X\T�M��X�����|?��-(w��'�}	rz5�\�<v~N��P�.�m�s�Uh(:��@W'�D�;駓d�<��d��;�%p$YiNe�G��vbd����Ld7����#�0���ә�������g�]5reN�@4��U�e.{b��ёJ��>�zd/ޑ.�:b(EƷ,2?�;��=\"1�d5,�Z�kB2vW�M�H6,T0�MنI(��ck7g�`���I��d�Σ��B��6�X���z0k��V�n��pC�|S��(��,4�OϿ	(�P�� �7�8'�l�(U�	s�6z�k���=,���� Jgh<,�a���NS��@zM��Yz,d�.�<�vw��'��h!���Fx�-8��� yɦ��KTx����H�v"�3G�#��d���d�QS�V"v}��]P�*ő.�ϰpB�p��6K�x�t?���O���Ï�E#���z����3�����e��3`�?�}�ϧv��鯞�T��Qo��	څ{;E:dӔ7��:Ic39T���O����Z�R��t��	b1`5�.B&��(tS�^0��W{�C���B�)�:��V�����L�yGs�p�T>+������s�r�������5�~�;I��8FQ��;��V)��J�"�Y0�4���Er��:�x���7R����'5*��S��o�L�7a^.P�)@GƘ%� �~���5�-4F���L�[��T�n���-[&^Lk��� d��8�C��~����7O0�c�B,�!YM��������>��������-߸�M2�@��}N���>���i���(C�[ �[����d:��^��}��	a1�J�YB;�,��VC��Kk@.�xͫ?=��"{�l\{W6��q�Y�nG)*I�׎��!I𶑴�ځ}Z}魙 7H��9�=�Q�6�SAT��?0����h��oe��;MeM���J��7>o�F��C����Y;�'�t����F,�lyI�p���cBz2<3b!B�|.�Ii�+�.nYs��
�Ȏ�m�%*g�2��r��U���"��tL�� C���]Z���ʐVGi���<J�����m��	�hh� m�3k���+��pu�]�D�c_y� &46����r�)!r���?�P��p%�>6����X�� �y�80�$�^�����g?ZU	�Po��g!�'��,) ��AUXP2���dI.����D�F ���`�R:�dq)�e�r"?Pc8Y9��]J����}�~����W���?��������K����73���f�'N11��ϵ��KB�,�+O?��?4��+}ϋnD6N�2�7wn:�N����IM��_���8����'���ͻ��T&a��
� �d�0a�S<\i�/���ن4�q�J�T;�@��>6��6u����"�ֽ��*_�R��j�t������_��:�^v`-�f�i,W�|�K��r�$�t-AL�YP��"z��.R�Rm6W���,U��)V�\���"YOs�U�����[��raW�FC��M��³�G�K��r�hB�	=Y�؊��OpE� ʓ�[�5\�V!�b�T+ZG�Kp��m;6�##�o�f��92�]�"̙�HpG�p��k��e��*u�^]��Q�|4�[�&����w�u�x��1z/��*�W�F���`���T$��U������7��߁x'e�����w, y��e�;�{؉��>���7���*�m;rݽ*��0����Խ�����_�`W�����z���M"�-$la-�"��cNԋ2�-ϟ�IӋJ���K�-w^R��s��0l�B�A�d�؄�Gp� [�Ż���|}]D��D�ؤtN�)��%,G��}����q�5nU��FjK��Ͷ�JxYZTD��I��@����d���٪�B,���k�~[s���B��+2���8���G��o	�%R�޾^qMƞ����a��Cb�����F�0�IC�k�>�%����k��PkW��3A��)a�݂y�I��<1��J��3Wf�C�3�U�I�m��h���`w�Ru���8O� 1QO.$�~3�+.u
�L
P�6=5����V���]+�i�h^��}t����k��F*@�6�m�=���<���"?��h�5�����S�G�_�GH�%?	�G�e["4�;Q��C��;T��a�BYϢ��yN\�7ISa���b*�`��ri|M�'�WWF��".�<��{�X�v�P�E����4���	��gt� ŭF%�/"�Z˖q�:�����H�d�����2doӪv �0�*�fB�z��s;2��QH�����z�Q�&���S�u�>z��ތ��/.6��z�XI,�i;Q��j>8$��l>���w?(r_��+�}�UM���,��"ub�����O�#�>�h���m�Y��xxs$k�� ���R��"f�MQ�Y����jmyrB�<�F	(��%�S��M+i�s�@�|~*��eA��oII�M�W�5���e��\��䛩�M�����vvh�u��B¿"�*;cJ{t�j�<��=��ڐ�����H��ͬ�fr�@_���6��W�kEԘW�ʐ>5g˕�����Sǒ��h�7��9��
�ٿ+镘Þ��"I�Aa��h\D F�m�D` �r��� �Q�i`��HeX���5����M�� �7^����U8����T�� p_���vç�sT�%��ZB�,o�M��,D���i!�����cl�uY� �̮d��y���A�I}�@y�,��j�#�`����J��,y�23��]�E Q�ϔ��V)�H_�!Obs	 �}cd��BRj�݉���@N��s�x�W[%����F��8W������?8�+u�r�iR�^G7Uv�st��>/��Y���~+���@��S2�1k ềb]^&�9̶�[���IYH���_���VALB+�H�� c�
�Yt�drs
}m�ŧ�U�N�H�r��V��=�L.��H]Ќ��5�r�9+<4�Tmt��s�ax%�mB�U#�K�U���$�����Kw��ѭY��c#b�a�-Z
�p���l��6X��?�r�Efꩨ,�t�T��#ZoW�Ɔ�'��U�.��0[��c.���2����4�u��+VS���:�8%*
[��*����=4ކ��d���2>z���W�ڹ�+Lh�`E'�J`j;�m�jh�1|�i���P�AِO��x���r�>oֱ��0UJ�G����r�_�s��2l^��2�_�j�岒�������`�cb��g��˦��[� �$c�M��(8�*�w�b���!�
 ��ur)�+"2���AP�˝�j�oB�����H��~)M[idN@!T(P�����AS	�n�U=i�o�,l��pĲ� �|=�U*�_�ͦ��'�\�R';h"�F<�Pu����RV����ۘ�sX�W𥁇��� �^��@�|���"�fj}6x���w��DN­������\�%�*���6��K���Ҏp}s��<��YG#^������%��[�/�����(ҬRA5����sLg�

�o�ͪ]d�֒PDR4���C�6��Ṟ�'����eM�����E�9>�]��;.�@�(�{�{t�t��N��gqJ*6�Up�R;0�z��d �F�޻�Aj&>t_2��չ�1��D+ݑ#j�>�O¦7]`Ѱ�:��h�v1ˇ�}cN)�D0���I1�ahǊ��9
+I�Ԇ�'�/A�=@N2��Ur��`�<M�ՇG�ǅ���?Ǳ|�7E��+X~�	��FCX�%��1�FAX�~@O�fK⩑��R���ڞ��ª*N��(>
��G�~,%�5�~',��~G���
��,�]���Q����e�#kh5��W��xG��B ����A��W.\�G�Hރ@��yZ���A��5��oG5A�EO�;Č�-��:�s���b(1��q��PF��D�V�N�IGa�W��Q��[��@��Wz�e\��;�6�ʍO?�$���D�\Z(���I�Y�����@x�&���|�����ON�� ������/��o�&)Gd������֫.��̜��KJ�T����l]7��;qvFc���� ���1��C?�^���@��`�C��