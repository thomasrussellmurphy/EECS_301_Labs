��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|�&���ڴzk^�2�z�eY��W=�=�<8�|S�D*��i]�g�Z�fpC�d�?�~���3b[/�'�hdΖ����n�^G�%�m��\'s��e=cVH!0�hCJ���|1zp��b�wl���kjs�A,_�eo%5D���]���8�$5za�i�""5��W;%bV�lwP��H������˅���W)�{ۻ(�B���M6�.��Ɗ�aN�Q�I���K?BȨ)���H��na�NM��{J ~��< �iLZ8�m�܄�sc�	hD7u���3�� 49섳�����:����t��K#�.�-wω���Y8]ݸw;kT_�)��|���9㥖����g������QU�kE*]�>���VL<��2B��PQ�Kl����e����oŁ^�vI�Wm�ZkQ��7ԝ��:<V���g�NpI�M���,v������}����9μ��+7�wZC�u�)�x���%�b�yX�cwߩ��F��׈2�dy�AȄ�Gu�-�r�C��)��ɡ�?V�ߔ&����fn����N��������O�y�.[_��~Z���h��]>e%�Ϟ�H�TM�arto�t�%��J�d�w�"�R��~t��{05E���-~!�;��25;m*Kxf�Y��
d��;�U#,`ݾ�Xخ�@�<����q�ܻ(}�H �H&#�NR����'z�b����ڱ���s&�H�Z���O�Á��;�܎�*�=�����Z�+x�\�]�'e���A�pg�P"l�����e2�H�%��y�q~��y��ST��� r�|6${�`�p+	s���1(H�Z?��3�#߽a� 0�ǲZ����{(������{�ÂRº��'��u)jY��,=����m9��"�<�Ԭz�:@�<oM�3�(��7�#����\��j�����,KÆ7��/��n�!(�6��'s�� ?���G�,��k�B��9'
Jz�����l]���4��������M�c�,�ٽ 2*��Ce���O���<K�#���E��O͆P���v���d�0��qzU�Q�fz�dL���S�dìdv��֒�J�q�]�:S%��2�i��7-�w���Y!9����F'���������l�cϘ��ӭR1e	��ܓ���L�0!�1�q� e1l���x�I�(��4����R�J?�+,f�A�'ڥxs�?���nI�-~�H�M5T��ߜ���foW޺�%9���{�Z�Ad�,-�UU�n�6
7� ��x���� ;��T�c0�-~pp�ýN8��ۋ�t��4G�nY���5g�_��![b��Ξ +���f��Smv{�=6$6��F���c�dP̅�@����l(�����Db3���+e�d ͥ�C�I�y��i��-��d5���	��ߦ���≇�8�};��s3�Ϯ��b>�.�P�T�q돧��82�����{[���sSS������]�����~��[�	�W�<p%�T�%\����c��V�;꬘H�[p-�Ͻg�L����:d�_h�(H��?��B�heC� qH���*&V�f4�;b ����PK�(�%q|�Vf�rd@��1ز�V%�u�2��8���Z� =�����(�I����A�O��'�3�CA}��^z�/j'8��;�B'�i7/��W!�s����� �D��K��Q�S��u�2��K��NGgi�8#��Rq�*�>����^��#k�4��~��Z���l�C�^���j\��Z�D�k7Rg;�h^H��)�` H�b��L��!�m��Y"|r����LV��]��
����I���ݞ5%ѧ#����w0��]�7�Ax�l�N����G�]8j��l4��;F���ޘ�ϡ_�_/>�2�N/v+-n��h����]�1��a^�{Ѿ~�ɦS,j"�;�<�J�i�zv�t��n���ߧA����w�7RIP�z�xtƒ�Ѵ�M�*Po�M���V�vQ\�A�)�jj4�Y\���-���Cb�/�(ȫA��^In��$y�%�o𱽊����#�P���,54��\�=	ع�v�Ñ�Al��)z�]�Y�+$kP�K�5;�l�h���4��VݴX�\.�Z�co����)|�=3����y(�&e~<(������lƩ�`r�!��F�4�X��%����F85g ��d��zK�����<	x=߇tSyw���X��L�X�q�VW৊�0�`���B�D�>C�k�[���y�J;u�4	��So:���q-�-��k�(n�0�*Sb��"s�҇ ��U�\b�����F��v����'4�-�����M����$� =+٧���8;@
7���(���Mرm�G�.#�_y��H���x.s�> Z)CGW�}�7G[��6-����7oӕ��Q��ܛ'��qIަ� ����Q1��M�Xзz2�[���co�;(+�� �'�"�2���`2uu~���	���r�f�hC�<$�u��/�|53�`���75�N� ��edd�� j{��BB���N����ۼ�^T��������S%¯b�VB�����#�@�צ�L}s.�L�z������D@3������%���=��B�0�/&��/`��̅������w�~�p��x�����)���ݚL3��8�yt���s�[�%�<Z���0Z(z �9���}T��ba��΢�u����a�r���&��f0<��hNH��%d��0�����]��^J��R!c>�c��Fh�^��&�O69�ch%��k��y��	L�{vR?1��C�M�������f����
.o�p|D W��u��an�`I�\��h3'4�7�*~�[��)��~@-���ͥ 9XF����:S����Տ�,�q�	�(�߮@:2��qڍ���C$2I��"�o����'���g��b}<�;M�����mg �7�J�0t���3�>��R2F�ήF��[̱�����S��=})h�:�ܠ46��)��.P1ƅ��.W�@qi�sn�2U���,�dC��d�d |ܷ犦�&~�>����<r:�����	��$d�����
^;ò��	��ꩦiqG�\&�j؄eC^��wj�4��RtsVL��Ø~�">Xfa�,���v��MM,O�-�3�u�@� ��a
CxX�;<�(o����_���S��ҋ�������|)5�E7�KYHw!F+z�
K�ΘX�Ubc���{�fBNO��ي�f�+kgXt��.��l�����C:�_�Tx DY�=e��lr�}�=����������� �!��ބ�+����θ�An����r����5]\~�90��&�=��M�W�
/��I����B�� V�����i���/5��ӹZ����'���ag xv�Ø��D��>�f�կ������v]%�T/�Fy^��Z��e4ߤf�1���;�7���G�xN̯oK��[m9l���S�x�33N`Q�RE�QER�T�c��Ҕ5v܋�0�#o�,A�B��~9V�ʍ��������%�M1C�c/���ﱍ�lY-����jWTRȥ��k����?=�F�"4�2/0zp��S$T�6���]f��R�~��@R��_�kK2*��W�
�>�K�h�e�SVG[�n�6/L�A�afE��� �nGkw5l���(c��r[�����=eY�j��k�I!Z����o��㯬�����Z�J�_W٥���m�$L���-O8G��OWY�⿰u��%8�\]'7�>@7i��J����F-ؼ��;�a#]���Kӣ��,]�&�0$Y�v����a���'g�EX�a/쐆�y���-8�;T�S�*i����u�X�Y?�T:BE���ΰ�6ּ3����JB��d4k�g����<w���M�M8�����-m�	�i���ֵ�����ԐK>���v*��.DUds�[����>+�P]��]n<�n�f���beE֓�	�oyf�j��r��v�M��\�S���a$�����I�܊�� Ps�嗢2»�����E\��c^���2\���	^� ��)+d��Q|��^j���d����<�{� >F[|���Ӆ��]��@�y�4���R���	q����{�����>�\���z���w�ǈ�Thq��@�������K'��#�]��M��$鿡a՚g-1�)�R�f�T���0��=R3{��h��*�q
��/;%<�_��t�wٺ���/a��:��]�}ٕ��y�!�tE�@�Oqx[���;�ˈ��td�sJi�b��1��� N��n�C��d^�P��6����R�5kt��.2{
`��'�5H�[Z���YH�O��N��ʬ���PeP��`BH�	�����8'��<�l���F��!c;����CJ��z��� �}pLg8�t!Ӹui�n��0Jl	����$���?�7�-w�gQ�g/_��ח��c��g2�E����̗�'��5ݥ��j �����پ�r��6
��8Σ)Å��?V��jM�5H���ӟ����j�N�����y�.M�Q'HJ"K�p)*���
�!�n��)l2�=�M|p�F���./���1�rzQ,��2]�~u���Z7���m5;�= �c5��λW��TZ��2O�J�J���9A,%*O'7�~�K<T��tv�q�u$�Z{�w�R�W� i��1i��v0��,d��Ǿ�@X��4����x�0H5l��5��*�0���پ��������!D��`<]��gSѨZ�4YSݝh��W���9u�3��q��ܭ�;� 
&�\����i���(��=�K����t���@3 S��Z�(׉��zSB�׿c�,������V�;�}ڼ��+��p/��78�S��qC�o;O�*��@Ak��XR����ג�W�������W�(��k��؋H��������e*�s�
8q��?��m�,!D����ل ׯ%��޸�:R�G#u�~3�͍�/Q 4�<�Yʍ2s�9L~xH��8���*��	��Iu�;z���i2q�d��Q�#��c�w��+��Qv{�.��E%��W��^�m�~���N�d����H���Ac�H}
g�%G�L��l��5���	���v�ϋ'[�pOX{.����fh�T��)��Ӵ�E���#�-��	���L.[$��0�B�?�(��� bE��6�U@�QΎ�S�
�
�g����9���U�-+K����!��5K�����y��]��8o����8����-8�rQ�뙶Aj�E{f���{�.�i(h�)�6�� X˫J�7���SMC��0wG��my�2��T/���v>�T�Kx�z�ZF̂�kEJ���"�8�1Ͷn�>�]\I��85�<�������M�X�9�Z��]1�O;z��
�2�}���N�z1���-�0����!��Sv�t2̍���.��K�E�ԃH��%��r�e�"����;��6����o�@��;rE����(B�g�;��&A/��Zv>�p�c�o:��{�oD�l�*�MN�:��1��c��ɭC$�D���[)�����<DNQOFn�<�`�H��d�nK��)��A]�#=��T\�g$��r��(�@��y�ߗL+�hW����ևWT�,�6�o��6f�D8�N��%�Π�n|]��ƨMIW�#�P�t�O�sq'�H�1�!y.�����������h�*�g�u�>K����^��C��ˌ�{�P}j��m ��6�Hw�2L0��F}�P/�;���*(d��"�^ѣB<A�f2��x��$�ey�6z�-�<ţ��߿�v&ņxh#A����6�����7�!��Z���Ka��0�T#�dsG/��AZi$�R�_��չ�Y��G.�I@��x��p�����T%�:~��VzEH�:%ɘ�%�$��>��i�l�f�Re������:n��7����l��槨�>X�.3#��@�8���p/)Tf���c�G�ѳF�̵�b-D^�PoNxt���_(�Rw�3LKN:��w�&j��¬dM��1	"�0��^z?Mq�k7,�12Dl!���8�۠�'�����=Tyv�r���z/BO@8�Ga���(Ԃ�
�E�V��2�~�Q��{�A���ы��dO�@