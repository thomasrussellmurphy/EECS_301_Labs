��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\���V�fnvx��ÍG_;�ȅe�~�>���9�>��Y;�0GP�5����ȳ����#�{���$D��P�&ˢt��#�����+�p `b�^En���!�+��xs+�m)�6���c�޹�e�+4����,P��V咪�B1=x��f <	����K�&G\yOkZ�4E�;�;\�����Ҹ����2����V\9i�*�$�������7!�br��	,�'Eϯ�q¾�OP��>���U��n��g�F��G�[�QI��]��t����5G�nwtDDn{K���Gn��sHѯ�d���6��\.M+k�y��x�E�h؊���rS�r�D:D6x�s��w�����J��a�U��̀�yeQ�����0=��о`�ƕUTȟ��U���J(����l��D)_�˾�,H�J�ޔ�Q��U�.&�L��ҿ��ȃ(�B�-�WJ\�X6��ߓQ`!�?G�ަ�}��g��\qo��E7�uc\M��i؈>6��q�b^N�Ƚ|q�`i��l����x8E>�ဍ�r��Ũ�f��g/�4�!��Փ�ڑ���P�H�=H��m��bQP.ˮ5�)�h�n?M�~bfI갩�$��S\MQ��<�5�a�l����F��6�NzH����X)����-oP�1���"��m� �t$b��YF,B8,ջ��TUVV=-w�Q�FUK�<���r�{�M�]*��T�����g�p��O?��Pq���]Hĝ�e�>��[4�Y�K#�hiG^�������- j������哟$�9�J`�mst࡮~e:%�7�N���˅���epK��F�3U���7C���3U�vvl�<��j���6K��n��IT��idli4ؔ����jJ��z7�y7 ����/�����\��02��N$]BR�*-��pT��P9Tt[�vB����1�8���#(.�/v�87^!ȼ�����y[2���ŧ�%p������E�{�5�ͳ��|\5{�<(�f&�y�`�'cT[6`o {�g���쯫�*C�3	'�՗���5O �1{Z�e���5
���{3j��pJ;�1���})�HS�m���[�}6�)QM_&���G� �u�K�b���|{2�rr>�e AQ��&.\�]�����h�ߞ�rBk�*����}"A�H���`o���!�%��9�����oYō�����v�z�!���d��:԰��څt��!��d�0${ �O/�b}.F5'�cg"��ғZ��XK���s�W$�������{?�z�9S��z�0X`jf�BA(F:=vųV�_g��ƺ1��sR�H�%�Emw�
V�mJAu�Il�<� ��iIzkm�T@ZM���Ҷ���wD�s0���.���Q��3u���ǜ�H�^k;zY���0 �DH�\@�C">f�o�$���JfAyαHu�%�1j��7�@e�Q.���g{\{R�Nl0�-V8Zj��/U
̱IZ�X!X���r͙i�'XH����gp.Bbe\_��7�h$ Ĥ�Ã�
� O���E�L�؁�����[�b6�n�f��mB����u��|�>N	�+q7��"�m�M� סS���#q��m�{8��� ����S9]E�Q�f���Qg΅�{��u�Wˇ��h�Ns�RKB��2�a�!�0��k��.��z�&�M�Z3�;�{
�; q����1�t8!�����V��+[�1�֧MjA>��Ҩz)������Y�<�߾8��
=�<OY8*��A�s��s����@<�Ė	6�̞ x4�k-z�X���$0��({2�>Z�8���aO��So^e�n���]{��l�!	�N�:�ʳ�\dq��($S�A���fe��Ue^������A�.�AI�Q�r�����2�ȷ~�~���n����Y�{�jD��\�'�ڒq~��;:N��@Mj�c�KP*��,��:�Ȇ0�Dڼl�9�4���v���25Rde��	DW�J]"tF�V�t��K�@C`��&��\IC�f��9��klf]�:b��.��u��}�,(�w�rݗe3Q7���n�n	ɣg�;��mIRE��$�^�@Y� D�ve������C������K�}��c$�L0�kSq
�i�a䏎��B�|���΋i��R�h���v����/�{R��f��X?��L-H�'�% ��P7P��R'��W! ���~���xu;�.b���L��^��7)�k��g� K��In�K�R��)xY,>�F�DHE�N��q5�3#��(���jϘ�'�	�ƒ����
��y��ӱ���e�B�5̋T���|��j�R
b�u��gq�����A0�N�*��Z_e�P�R���"�6���ć�|��o�Ѧ���%�t����Qw�ߤ�+��_��wq�I����X7�BkP%�=B�
$|�k��#��&P�ɡ?��}�'�,<��GiԊ��݆�ֳU[���6�"Ȳ��?n:0<k >��1> ��ߢG>pV�J���^�h��������b6dc�Q���%������1�٠�JH��X~@ϋ��&�j5�Z���bC��#E"�`WqI���Ct�eg�.�D%};=No���Q�c�p�2l�Df<���ޒ��RM�Zmr�B$�Oˊ����soqw�:`��e"�#��4�)i�����4
����A�iT�p������I~���lGJ�W.mܫ���uU��5#ն�X1�F�=�3�������+§D��"�F$�(\V��%�a�שh`p�n�f#ǲ|iM�Z^6^�M�%�ǜ��}^�e��&0>Z�� Y�Ѹ����T-�sћ�s�$�}�O���9B�ף��\)�5V���o }_ˁ)5�� /MLyE�eۛ��e�[v���Э�g;&����[�o�ߞ����|My47;�7����a��utBRD�q�)C4��HuO0 B�&P���ҏA�ܻ&<V+"�z�5͋�Mq��*��GZ�lݩ�"��7�B�r̓4��y0����a����=��ő�o�T�����q�@Kq�m�a>��/`Tmtft:�ںd�T������'E���<P5���-'6�jA�G���mJyͅz����&O]�$�0�b����p;Qg.����$��Ēcw:�k@{�#��7�p���F�Q
m��L��F'b����j�0�����՛V����y�>��w�<�j�XTu�F��9���qTⰴ;0H�Rt^e�sZ���a�cAc�!����T��E�vU�?��v^���y��k�l'��ᶉp��%��D.t����f�K�6ܢ��L7���}�En%��b��wN�/9��]�c��X'd��S�	_�I�d�S��eo��􁼘b�g*<$Ep?ձ�ta�=3A����#4��la'�K3��X\c�)j���J�ꟹ0R���0 ��$��d9u��p��h���׌{G��έ4�~�˩��]^֛@�n�{����� �,����	�!�:�0p!P���������q��[T�XN'��@�z�yO������z$ohu��t��H�v��p�;�Hsi}��5-7�g`�@C����ў�H���і�.h1e�䚩v+�?&��ۖgA�RI[��T���ӝ�-;����2ҷ;9H8�X�n0���qԲ�&h���(n��'/��0pnBSQ����cE�\�������`=G}�Z&�ܙ=W"����0JrϋQL����`( �@��م�J�y78���bc=Ԟn�"ˇQ�f��O��Lcǰn�)����cPFz���Q�%�U?���X
�gx�e���i J�3�y�>�1ȍ���������N�K�_��L��@��;$5��DbQ@f�4���#��&S҃��hn��ܒ"×Vc�c�&[���9^v��)1�ɦ�z���Q�l�ew.��;��Zl�������c�n�۷=�.�[��`X�9�1}ۀt�f�ʲ�[8�4��@;�`��vt�#��6~�:��'�H;T5�jaِ�§t�C��%ax yK1�'��P��
�5�xlĹ�sv�9J3y
CA�{b���r�Dr����bp��IV}�"ee<ެ��� >��y7����������� �<� ��d}���2���_ۛ��\N��۷��3�*�ȎF�xYi}�T�E��Ψ%�(eߙH�+��B�k#��N�4�gB��;/�ĕY^A�b8��B�3}a��E�?J'
�`�S*蔶CJ��mM���'8x�xf�zRZG�����r����2���k� �W���QUD�^�(��	B�!(��K&��T㲡�!��dH�"؎'}D&�8��#��L��~|�1�\�3�6�<����&�P�1|���T��K�ͭo%9����9����dK;�*�N6J�;|=��q(�i�V'(,�8� �D���l�<��S 
wgp��o��ύ@	���.�����R�s�D'�����ÊQ.~���4Y<,8�Y��N$� ,���+�"G��>)��z����Z��'�UQ��Z��)��\�o�T��4��܉�����,Xaa��}��{"��'z�\��o��(�B?&�"�WqP�!�N�
3�hyV��������H�T �]��">*X�D������C�t�.��CɛJ���XZ+dr'e�f;BQv��R��"Ӷc��<*l'�x`�-����B��1b��W|R�e�,��w̋�T�Z��T7C&�?��v�h��aì�xV��vo} ڛ�s���|�xv՜�>�h_a��K�-�J�QJ��Էbb_KA�i�!�I�~�ס�.M6�%�dC�4H�E���'$���)8�a#}pZ'G&qT��V���f��)Ao����`"=<3�����-����C�*AJ��E�E�տ�L�W�.�ܓ�A�q� �uR���,��e����+�?��.��U� NX�%G0��yjv�t�h��y�F������$d{���GX�L��|c!;{H<V�:��uf�\����D|N�AI�/Z/�*��/N��H�&��(T�l�KΌ2�c�&�(Ġ7yrS� �~X�������*�<he�f;p�Fn���P�s~w��G}1�'n�#�pX ��N���p�]���b|�i�U�J����3&��7^7�fޓ�f)Ӿ��z�n+p4��y�Ā��S��V�G���U��s.���hX�L�p��w��Ž)�.t⨱I��w��hX���d�̐��.m��"��,`y��]�y#g�-R�,U<aQ$D/��,���L�s�����P�(�ǜ�s�-aCק�ȕar��O��&�7�/���.�^h"�""FVP���.� x�UsZư���;H ��T���:]��ͳ{��RXՃбY~������
��K��9uX��ȠŮW�!z;]a��66�8j$�/cj�"�5z���3�0��������\� K�զ��co4�n!�S$uձXfor��F�������t�����G�@ᐫ������Z����˥�BH�&�A�&����G7��̤(o��}_ڳ�wz�yj�?�@o,�L[�����-�yD��9�ӭ�h'\�Z�Lni�?:Y`�H���֭�
�0�i�eёuY����vZiȅ�vC;�7x�:��LC"
a&��,��g[r
���V
�G�d�$�3L�����4/����Hc��.�D���i�;�YJ��P�Gq�W��t�ʧ;���9��D�`3�u*�,M��}�&u^����BŸ�o�C�!
�:�m��3��yk�t�O��ܺ�K��v)�,���`��Ο�գ!�L ���r�n�e�߮T�DW��e�I���g��[cï0�IV�^C},�	�������U*�N��]�昿��g�� �������Q��7�'���Ad�57�bG�x�''���$�����:ݧ�r��0b�k������	�fe]��kB�]���{�H�_�i�Y���~'ʦ��@��+�\�]S�(�ia���;�I�4]3�t]�jp���[L����B2��@o�痟�½��&�S�F��hY�G!��P�=7���R���1=D��!X؂��1y�F���2ޤ@�Ru�)G=,gȮ�,�O�={�Hǃ�#���h�tby�v�Ь.p@�g���I�{`Sk ����n��Z�3���g��t�^�e|?
�]�p�!�E�>���Z �8�����L[&E��ߵ�^�`��s���? �L���G�e�U�^��<�&�.�Mߙ�V�M����R97�#C�E��)�}4����$��N��u�rn=_��6%lq���R�w�h�R�=����_��k��������;�l=��{I�PX��>a�H�t.z��72.[��_��pH�cӸ��$vռ�h�U���xK�6�1 ���}:��Ta�������b����h}g��:�R}�ފ<�9����P�v?��8�V��A����ã�w}��N�{%k_��DIa
�"ϯ�Jc�����4LH��=1q�O������50#�2��^��mڏ��"� ��p�6Ss���D�7hzP�d�'-W*�h���^&�ۺ�)�c ��{��'ߓ�u�*��5�:a�y����Xnh�h�s���`�J$�dx+A-��.�t�㼰�X���t@���%[��¡�O�J���P�x�b�[3:�%����$��x<�0�R�\�3���X��L�e������0�'FEd+���k�3��nɥ�>F������b��I
���#\��K�\�x�~����(��)�]�W��tE��8]��~�Q���0��ʚ�x㚞�mjڈ��Y���cƄ��ɸ�>��>_��H�Ё�q�Nǝ:@@t�顏��������T�׆�Y�,^.�%��"���?�P����3'����?�4~[�.����Fb����Gi�v�'Lͤ���~h[�*����P2DG��v@*�Z]B�	����Hp%��=7�� /k ���U���r��RD$%LAԇ�`j��ۋ���3&�z ��F&Q�1��O��R��).y�Ϭ��.qf8zj���������l����Ҩ�'���r7�=�u�8��_�gM���j��q&Uc����L��v��G�"��Z[Š�3�Ÿ��w�J5�Ҡ�*Mw���(X��N%�
ۯ1�_��~oK�s�o�2�2�]�_-q� 2���$�x\8:���$*�N��I��
_z����I�{c�i���1�[W�ȸ� ty�G��������\i�`����IH��./�『kҘǢ����Yb�ɳ>H"����K-.	��{4�/'��eGQD٣���o�( hv� ׫�;w���䌑�dg1Ϙ��@�b}�/Xİ14�%����2�ȸ/4jW:���(����������e�X�_�7�5����M0Z�qc�in��yZHR�MG�@5zP��/{�WVɮu����U!�B/;�3@�s�S���E���d�H�MA;�R��
GP1^����"^Z��dDݡT����WKa*L��3SM�N�n=m�քWω�iWYf�~��N�r(ۋȄAfׂG��^x=g���+��[�G��#��H9K�^��Ӧ}]���n���&y̋��@��h�`H
΢o��֟@������%Xu���5MR��C���z�,��T�(رb~��� e��5�A=.��F�֡\��A�G��������'ҳ�/�S�/�B
�>|���,R��$�nA����E��t�S����`<�N
j�bE ��������k`�	��݇�Y�B���ܬ�+�]J�G�Yrf��y� ������J�zw%��V�����ASh�v�4�Pi{�Y�<8D�[��I���rȱ�V8.\��2��/4)����k��&0؜�(߶y#P.����B�>��ݐ���}aԶ���\���-��:J�d�o�2�Fx�� q����~�O[�'��� �s'�-�C�h[kDH(��O�l�5�Mp�uV�!k��5c�X۠3�I۟��:+���%/ٟ�c���0�?�5�Q�M���B��/�e��/%E,��vE������͌�3�l�Q�صv�"��l�<�Ǽh�x��uc��5KҖ\�����jM�wL�}-i�r�	���`���7�\I畀��D���c�Z��8N	�[��$�ϩX����C+�O��-��q���2Voij��z�|U uݣ�{`Ug�ɱ=C
	�Rd|?A,�3d9xG���g2��t���؃\]����s����QC�7��bD=�1�?{u�E�Lտ]�G7��lnJ�{�(��S>LQ�H͔�x{���^���8��H����rp(3{&�K�2��jko�����t/�@�y�o�A��q3͒z����Q���[FB1/������ǩ���+�H뱆mM��1�:.	���)�I1��L=q�r�D9������ɂ�����u%n��oJ��I��?�"��TC�6�"旡$�uE��"=�7�<�����~@���=�F��1v�H�#�������&�b��ՁÐr�?>��K#��P���5K�!�����Yh}Ӟɒ�ca�3k?_7�v�jX56Ɋ��؉��k��ʖ9�FT\�s�E�� 5��*�Qp�?#$�A�[bDD��ժc��I]9�����>#��.�?k�|m5e����G��������M򹷛�i�V�Ce���.GՒт��a���
s	�yq~a����-@�uN���6�o{��*:�D��nOAm�muɵ%+�>7��悡gv;��� 7����>�V��13����k��[��'���E}�#)�[0-1�r�M\Úwa��\�?��p#BF��HJ��R6���GAjC��I�6N��p��Yd�h�='�����4a�!����ti�A��x���I����	���g������Ccv)洯��|��U�:K�]�����`2mU$��%�����Yz"�O���K��r�v_\I�� �ݿ^<��[��'�)('�v��)�BJ%2���.���Q�\�䋴�wf=D�^��6T�ơ'`�Mb<�O%��]A�90�k���vF&�`W��u��l�rFc�09m�}Xf�p�#\a��w�d�}���y�D{�SR��w2�5�Ǳ�E����nk�r��H��� ]�W��cۡc_��:���A�$i�#�u�G�r��8.�7��)~H�"Li;�����$��`*쥲��|,�XߘU��A��~�q�*3[��GQ��Ўr~�ru��/i�����'����`����E�5�WJ�EgJ9�0ZOf�F��!-����#v;65Z��wf)�>� m�`Y�8F'��!�`Ϻ���C�I��Q��6ٌ�[��y������"�C���={���x�	����^�����4�p��ž��d]�1��*������5�N�)�"��E(�)h�peDrOj�CL��K�JFP���`�_�� �YD�3�Ȍl���fܗ�|$�{�ֲ��U��t���P9a@����� t�%������[�Y�0��4��I�:����+��c�I�Y��t.�ze�4[S�ξ��ƱBVp25&�^_��P�<�wg\�"��
��A���s���z�iQ������:)co�*��2��:;2��EP��M�Bą>�ڳ:�hSnjE8WOOn�"�3|*ϥ�\��[�����+�a3��?U4�t)d�)f��b���=l}��L�_ό�d�h�d���!�'�3���RP�W��o�����n��2���w�,�X�Ԣ��ı|$�ׅ���6b���_c�=ἄ�L���ɍl'�}�TVMEe@>{�֋��,x�,qW�����KQu�I�lچT,��m���ۛ�%p�t��_��g��Y�ە��#UoO�r���$�4�A�(N���iFF8e�;> ˘�>��>����'8�i�Jk_���3�z]�*�7��H�&�e_�o�m�.e̢: u��s�oꕜ/	��Q��� �v���&z1P7Q3�lE#�Ä�A����L���7��Z�u��UX����E����D�뎥�]��j\7^����U�D㭄�T���i�keNB�|�5SDL��"��q��V�f7�ͺ�J��O���mQr���V�G����@^s���va�O9���?�!���C�1�A�{�²yHF��e��!���'�����T���b�u�Z΃o/DZ+�a�YM��.��x0��iL�;���l����C.]�.�y�dE�Ң8lWЂ��U����Nl=�jÇ���3<g��{�Å`-ЮF��`��+�s{��5���B�ڧw�o��χQ+uA��])g,$X�M'�
ae͏�=����b$��J� ن�O�")_=���7���H�U��b�k�h��ۄ�pa����9�9�)�K���%0l5��|Ac V��i�R@vjz��D�j��;ۺ
E$�����;Tk~4^�B���f��%�{�T9�KEo�Gv97H��ňG	*|ԯ�$�;�������%<+fN)���;mkt�Q.���J���C>{ā4��8/�)Ph��ˀ[��c�;/�����RF ��/t,�p���ܢ�E��	]��߀��/,��ϫ\Z"��@co�<d}�363[FZ��d�6e�ړŗ�yR���Z�p,ɗ�I�q}�\�LS��V`�f+�11"O@�Br�!
�_]�w�S�j���M/�����E���x�xö�]y ���A`i)�Vp�1ދ�T�Pޯg��\�:"��֛��N7��<���=Ȣg���!v�0ԝq��B7���,��X�7��Y )�)�;)��$��+�E�,8��T!��
;i�E����8���4:L��jcK�����#�JM����C)����s����L]� ��(nQC֢�b̈j�jB@�WM�����I�!���,�������G�Bc~߉��%�L�f��=cl��ƋOC�a'k;�Qy~L��]
S����:2��j�z�5�zw����xS�l�e�����D91�"���:$�3 U�k	JY���}�j�2*��]��:_t�i�`�%KX����2��x~�m,�Q�E7�.|�� �haA�ֶ4����f�ʒ�D������\�R	Xܯ�-;tyY��^��=�i3�'#B��)~ZKw�X� ^�M'��c���߬ ���	t�?j����Dޮ�Nw�N��A&�in^�c�J�ҧ��)�KT��L����툜��),��}��Ȉ��O�1����֠%t�������"�'����i�z>����f�.������ҧ�T�<e.�t;���nc�J�d��bYa��!��^[Hc1�nD�Ov��	i�t����(]���y�y^�e*�oZ����⋰ȉq��L<�w1���b�T8��B�P����vM�#|E���3��Qu|��n���X�6zQ�QxQSᚦ�<|J.���f=�����׺<�9����叹4�$�~�o���c&Oi��ZkH���/b� iB��*�A7pcX@�<l�K.e.�m����'A\)-�d;:ae�������6�|�	]����C�d=�|P�˗�N�x��	B����a�Y��K�5wE������M���&��j��
�e�jWX��d�� F�M$aq���f��������R�Y��8�R{�� z1�g%�!���LN��W!��XD{�+É1�䢾��@;��S}���o�0�?JX��O�$�g�W��Ѣ(`+%��p@�ѵ��$H8G����oC�s��u�S�2��G2��|S<X��|�|�b��߁�
�qST|�5�ƅ����Or�B������;�	�N���J4KѤ��;� �M�E��yB�������t���qHV� �܂����MRg�z��{`��N|Ӎ+��f�DE���W�*KŽ�ރ��*��n�0����^e]1��z1��\8�?����pl{hb�wo��6��'�����}S-݀H�͢��ڝZ���v�r�;%��{��Z<=8���B�αm�\�Oݘ�Z5񬚿�z�i.�����PR�����ܼ;���>)]㉞���?�`v�o�&�'x�w�. ���fg��+(!h#��gS�f�Rɬ��C�(�f�&����p��'Nb�N��?�>Ӄ�H�IM:'�#س�eߙ`9�M�;���'i�!��}ma|Z+�$�����UI�� �p9���<0��A���N��k�:@}�9����i�| bL4�J�֝sؿ㩳�G��@����C�o�A�^V�u�)�尬,Lv���2�Yj C^4����҅��D�9y�'�;RZ�J�!䬥��Eh"	3Fv1]!�'WyAټ1�@� j\n�V�$� ��@X�nu�d���8⪌߈`\'h�p���	��(ۨ�Y+6P<�Ac�yz��*�K���:,��07�j�B~(9���ƍ�/")!ډ%J�4���?��Z4I�Q��&R���4��r[�Q�)/NGp�z��4�\� ��PȄ�a��d�~�Av�Z�d)�n̐}�<d�?�q�\�	�P,mC�ffW��(��j
!u=�	���
���1���`�L�c5v]��3\�R91���, ��gQX#�s��<:���`z����:�t5P(j�(Ξ�x>�g �m|_�]��/`�$a�V{2z'�OG���&}�ɽ�e(�^@�m�:�aw�*��"���	&��ڮĨ��Vz:���
p�.�`�)u�ĿV;��R�~�P��	�/í�� A[���0+D�f�e��+�Q�3�J��o��Jmv�+U�>���Ĕ��1��P�"�?�%)&&D�t�=���
L�ܲL�����~k�J����������3{F�8`�1�܎��xc�k��@4��ɡ2B�'1e�(�zbV47�'B�0}ǰ]��/M�*%c�b�4�W\U�὜�P��F�߯����v��bN�Q��wgu�	�$#N��.��������E�i��>~�GD&��?�&N>�`��f!�Xl��lz�eǢQ�<LU�ܛ�W2w�F����q��0p/>�mh��k��y$��FGx��V�6�����ۈĉ����߮�	zmr�u�'�B�*���'1��j�~&}�{˨�R���XGY��1{n�'ZW��6������A�`H�Lr4.d<��"�/v ŧ�������k��!_u\.ƭ���Cn�d~�8X�D�Ҿį*O���s�nE���(~m�f�×<`:*��LR�?$K���(̨����k��;`�K$&Wx�)آ�����n>h:�N�h���e�^���
Zˏ-�i2�aN��BT��e����/X+���/���l������Y.:�b7��?[q=���O����I,ų��_��$I��qr��3���CE�-��5��&�i�^�N��߃�K^bn��R
�'"��IU���H�����p�;�!�R�U�������ݔv��-���� ����o�uz� ��5Evho��֗dYtۤ�xG���oCQ��6.�:+�4e��)���.�|Q�Ԑ.)~�-R����q]\N{$-`?4�E��4c+���j��j���+�2oc3)��]�+YB����l��M�S�]��쭜ȁ��l#O��{3-�V���
^�,��8��p�K��D�}�`Ae���tuY�84+Ԣל�E�M�C6d't����E�Ե�"\���F�I[��ˍ���1Nj��4�Հ��Ut�Ȣc��F���0��QSBn�v��^+_��>���	�O�T�K���Rtw��ͅg^�����U��.��!��(�������;��z]]~�d8��n�Y�K��Zq���`[L�so?�&�8���:��B1@��֡߂�R����C����NNp���������8�]���0����k�4:ϬY�����B-&˂5D�Xi�8�h��譝��b , �'Jz玱tv���A&������οTŀ�������lV-oE��h�C�6`���j�	���*s`���	1�J6�ߎCr��e�.w��%���'�9O������O�
�ڀ�M Qߙ�&�
�0����Mz�+��0L_m��#hU�:�9*�;lakv��(�+ːWHM����3��ˑG���[l���tp��9��Tm8���f���̫���J�CZN�хS�m�񾦌�Q��hO0dЧO��(�l+9o�������'��K[�{�������|OL����5fܠV����[�$^�m������Q|Js!��Cq�VHZ�6�j7��6Q�AaI=wU>������b%�~����PI<0�fN^���M����L�Z_j���_q�ԟ���"���
��o����h�r����R)`;� �����b�ѡ68�����;�JS$[{R���D6�M������Ԣ�6\m���p��2���m3��S.��Ǝ
��3���8�8�t	�̳`�"����	~�լ�8��!eM�WA#�ʇ����~���G!ӝM��|<��c=�_N.u�H̃����Tx��B�g4�>���@'w=x���߹+>K�	)|HjF�Z�M�Z����rʕZ�J�>�py8\��p4���j�wq���.�'�(�N�Wk�1\y����� )ƈ,�ΠU�OU�x�┍���{�Z��i��g�����l�]!X,?`�7"��HA2�>oK�/�V������>w�=����q�m$���ʕ���Sm�h���kl�����	4j�:���u�L�.\$e���J���n�U��T�(��C���L�`�U�	���D��^�¼Q5�l�0�*2gL{=|(��/-��oѐ�Z��FOӺ�ݲF�吚�o��]�#�� ��~Q+L�R����S�~���*;zZh&�ݧ<ƀ���4�e���%ۨ��ۧ���I3Us��M~=Uq;���\8\B��� ��겝����S��H&=H���v�D��N��	�T�{� Kl�q���܏?Օ����Ub�l-��sT��@;%�$���W�j�-��;R���Z��E9��#9�gNHd�C��}�Ue��y{cyðF�O�a6�%�������E����v��h��%�7���.4[\V�|�W��ȭ('37�Ʊ�Z������v�9�M����^,kn����P$P�{�K���C��Dyv�?ѣ��޴�
���|*L~�>������R�#4�Q�O�XXkH ��@KQD>[AX�ӻ7�NL^b�;z�oM2���o�t��4?�����f	��HK�.?s��5����YՄ
�=��a�����4ښ�doP]���$���e����'6��$�#��rfϴ�j]^�?�&����A��T�y(TECڒ���ʓ!�s������o}R�׀��4mmT�p�A�y�͇ �t�[c��o}W(S�;���:������u�����H�|eߵS�KԺ�"8�i`��s ��R��y+�����R�;M@lj���9%|B�H1�\�f���Ӣ�8���F�s�����2'���z�԰=��*^ZD�Ⱥ�
�ln(�`�$�~���Ɨu�@����c�!����0D�*�o$J�����.l��F%�h�Kjt�o[�B�&!��Ta�I�Z�I@���<�pQ��%j��h�I�c�1'Y~B�`.>ݻ>�y!���Q�}%��I���2�S~�f�o�O&�|��j�b~V�;+E��D�U���FXF3RӬ�b!������Ot�L�v��,�&��d�n�<��[ lU�<�(9W7ɧ��F?9����s2Ck��j�[
��Q��jz�Ф��x�zbm��t��d��$o�3���1}@��6T弛�Å��t���+�`ߞ�{Y$B��J.�dRBo&�:©�jy�?���/a8���m`�٣�{�V�����j���Ѭ�+���=�}�slL�n~�����/	^��.��S�^3ݍɨ�d�����ocf����BػX;|+��>� A��l�ǟ���&��jN��A�,b"����#���zq��W�\s�U�RWsI[�j\�&�F�p�
��Hӱ��2±�pc+���.0���L��\yU��*�W���	�0�D�����?V�A%|<h�B�.�lY�~�M�1�`0sƽM迌��8(h�0�]_���hJ':`����P���������>0�MԆ��m�I�y!hd~��Y�b�a@�!��)2u��]"8����O��S4�ܜ�āT�1��܃F#C��K��M�4Р���_d�q���e�I�-�'�$s7��
4�����e(ڢ���qm��+������N(bNeS>���3d7.�w��Ew��%'�P��tX�i~S�͗����W�Ad=k�ˊ�������Q�)�L1b�g-���Fem46��o���lԝ����/�FN�!��=#��b������,s[�;������.�8bI�����|q��?C�����QN�oM���^B<j秳<�kk��>�9�3��!R����Ƈih;��\���&�m�̋���"3@�5l�x��S�V�z��R��Mi�B�2��N5���am��^�,��E��Pz�aM����A�vr�|�r����Ɨ����y&���L�WZ��5�L����h� �����en/픏��֛,�u��l������0�
�3�KqZjB��p��<��JE��d��;�0wQ6���q5S7׹G��t��/PU^4(�h����}�߫����>�
�ճc���yՠ� �L�91%S��^��cw�L���$(SV>@�
G�l&����7P��~���Mc@�6�	Xb�W��"ڬ���`�ƠCP_��U�"3� kG��e	r�	$��)A��Z,=�{�64�yK?k6��9/���e�L��Cz���;;9L���0?=lSs���1�	�n�c2�2i�[:r���ےi\0E+W������q��gHq!��)�$s=G h��i���l��+\�@�x�vJ��������7Rq-'�VbJ��p	�:l*G<��g8�UR�s�=�,�sQ��q_��u~_�R_0�3���Z�՚rp>�+F���*KW8.�X�aJ�,�U�D
sN7��Z^8��Z�eӗ��Y��a�|����k�n03�FxS�R��C:1�HJ���N��,Q%;���iȓ��?-����ب��CGhR�\��oa8�HW��_Q�D���Ȋ���?w��AV^��K�/}v��0GwҮ�Ƽ�����,�=�P2��_�V�g����aPd�^�3�@���gv�,�е�z�=�Z�Ha��j !�q�nM�9�vw�C��sP�#��@M�-�R�Xe(��C��q��#ޮ�D�fL`I�t�a��K�"�x3�t5�)P�X���-�s^��2ȁ�}4�G^A���M�˶�-�Mp$�3����KY ��{�i�܅���.�n�v.��k�4�er:w�`��q$G�OF�;��p�s�67R� X��2���Iļ{��b4��W�ڔs�ٌ��y[�n=A?�r�A4J���ؙ�,k������o��Z�ʜ\pW�8�Wj�83o�!�s�>l���s|�t�ʎG&��� �������d?:�6�>ah2Y3���_djp��o6�U�b#���-�{'=u����C��%���,*�/�%	�t����iLH��G>����i�t���������ϱ^Ov��/ǧ�Ƶ���H7p�v�߻@�ħT���|�_�������Ƀܙ.*��xI0��g��|����)H�_��,�<��_����� yÊ�t+w���� �5�X���y&y��i��͋͞2��t�1ԯ����D��7 ,8$��w��w��m�ݬA���bM��tEA���V�v��[�P�+�(|*�l�$���>��MU�TQ����������d+L{<�01q��Sz<<��hʙ[�,
t� ݠv�S@���s�HK��s��3O�����ia7�����I�е�O��5+v4TCg�p�5��''����hM�o*��;�ɞR;�㛤�)'���G����.z >h'/8�����iKYu�2@�����6	Tez�'6%R Ѕ1t}�ƁbR[�%Y��M攓��#��P������D\6�k�����_�De�T�j�D�����u���#o�=	���#?��5Ozm��f�,���ޅ�:U!ma�@V'�۴��a�S�?5�PE�G�����-�B2�e����}
���f ���������
�}�0=�_��S������:j�օ9A����ͫqJ�h;�[]Ot���[��R.��8��%�������"�2�qa_