��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\���V�fnvx��ÍG_;�ȅe�~�>���9�>��Y;�0G+��X�LP�n�O_�I�	B#Z<��dٌ4>����(�ʰ�j���j^����x0�r�,��]She��w�ຳ�&�/��B���\U�0"�b@C��@Eܬ��Z-[x�"5Ʃ��"�rgƯ7�Ѝ]H�k%���)�������Rr��ˌ ��!^���V{��r�$���=/���j�]���>��W�.����5Q�tl�LF{5�ć��\��0c�3����t>2�8�
�:��(�ю�%��
n�_�|��/d�I�7~�]�^�@����Sު`��0,٨ΐv���k�Ct���Vn37^|���P~�}�p{[�׵�J�zX8C�s���ڮd}�����$ %�"��-�|��;f�ٱp�;�dmA9���fwG�r�nl �����q!�.�E��HT �,��I\�@i��I�m~up���_�;;|[����Q<���t��_#S5�5>�O�M}1\2�R��'�J������6�f�#�r6e�OŇ��K]ڬ��T�o�'+?����I��b�!��=1��χ,A���V�L�,��R'�3#N�%K�w.%��,.R�R5R��v�"6��86[��?[�y���gpŻP;�ШnF�.��� �]D�d�+��K��0��al��A���U���dI���H���]��J���(D��J�NҦ��T�Q��̷���� c��Z�*3˥�L��:�%^���X�j��V��"�03������MX��ê9�F�7��{
>-�$!��#��s � �GtX�b��IY&��e����L7�����j�,9��u}�o�<Y��L�����)�$�M�z��I�}*F�V��9
�AXA�M��b5뱓��*ws�� �nj�np���w[iБ���M���aZOz��vÔߜu�	��Q+dv+��Ɩ5����螩���F���4��JW(Gn������X�Ԋ�X���#:Ђ��6�1�������d_���κ��sEk�"_#4�aS�ٛ�~���p�ُl!3}�4�'u��Q1g�n���_3���C4��EU�*	Dg`s�������^��`	�0W��Co|s�2ު��#��7R��U�{P�����"[]���XN�~�±��<�=� ���w:'�O\�Z� 1�)o����^c#��n��Y>�Vo�%�I�Tc���i~�F��~ƾh���k�L���Ķ� �e�]����c��uP��A�J����ْ*}�L\�e`�ii4o�?h`����!kSw)",�a�P�/�����x�d#o�:�Tsyp2�T\�`�����xq�x?���&^|^ʆ>�%�a��wf������2�(���ZNvaT~����<���&Nl:��Tgחo"n�5�S���Mq_�Ϣ1F�a�m��t���ia�"T�$|���)X��Lv\@�P,�^�xT Nb�T.("8|o��̓�2"cvP��P�&��.�FN��}@>�3YN�~��nhWn�f`,�A����� �t/��:��M�<�|�:��Nj��|��Y��30F�ը[�wA�~5"�5u��j<u0R�TY{N%c	�RZ�R �$P�	�,�v�*������տ�'��ᇥ(����C$�`�0f�M٫q�����%<�%hBROK��5�T]�0��p�m���ŉ�y*�(�1����+�H$����=~mg-���T��N#Em/� �G}����=�M�	%:�A��A�!����flИ�<ޘ�KV�.�j�����ѡ� Qs�.P �2���2���~���&�]���Q�70�hy"��d��º/�i��w%|�Lv��!��z�)�{ӖNQ�Y,��{�@���_�%ö,D�`���w/+0�c�����)�*�ۯk�Q�u14,�I� zrx1�ό���Z,���{��ۋ.�O�( ��n
3#I9���� ��+�Z���yD/�9;ǁ
��+�ǿ�N�sDH�gD%�?�m�a�o���	�.�Aw�C͚]�:��@S0�"��{�L��m\X���ơ��'h���iP�����p{�[f�D�Y��oF*=��оPa�� �f6SJX���1�Y�*]g��=rQ��16�\A�	PDS����1=�?�h�s����X�1Uc����1�j�Vw�c�ތwc�UU�i�**��}����-=?[;��d]`���i�i(�I�쉺���f�'��`������[�1�$t<&k�F�^�C�YE��2�\0�$[�+����V ߎ�ķf�J��P�-��]�����ٽ�)"ث��B`�r��L������p'�բ�Ȳ��L�(�'���pt[���o�����5� ��>f5��^C?S/wW,Kk�۬z�+�T���X�L��4�����o]�M��-V��%�E�ԫK�:�t��sXl�[3=TQL�����R�S3C�|l�_EH6���`1l�o�m0�����S�W�����Q:^�C��֑��'�!*ql(��6�[�%����~��߷���h_�;�Deg�7`L�=nWg`�p��e�yğ�rSѵ�ٌ���
�Ǆ���'b�U�/�Ab��F�ŵv��_c8&Z}����qsȫ#
N�.�<lT:Ҧ�&g�
w�bi��7�����g��$5�ei�x[�X�����MCp�͙��JUIn�FN�<�e���}ʖ5��#k�W��p���첅�+��vȈ�cf�A�oO;A�4ΐ�-�Kj1LU>֖���O�TT�5�WD�
]�b�֢*���/�Hls2��Q�Dڱzf�g&,�dO�����:��X'g��uD���څM��&��a���v��6�'e��C���wї���3谳���VH���ޗ#�i*@��C���������,ᛀ+؈�ܲ�]��{�a�)���I��#dd��E��}f$,/ �W
�K�`��a���� �8�T��r��Z���$:<.R������@+��'���֚�gH~�&�r��U�	/�������Yr�;����l�N�\E2�<�N�����}�_wg��DG:�K��:�L��/��NV��`�>|�h�'Ɉoͣ�峜4n����My�[5d���w�c���^Z������[#@���A]*>���l�o}l����2���y�#t����?��1Rє��z�1_�M��1>F�ܹ�,���7�����gg��W1���A"��)5�xF���]Gn�ki#�l�Uz#6��ds_����lDv;�=��w$��N���R��4f��{�Uy(�;���(���"�z����S���{�r��?�,\LO���*ҧ*�j(��!��g��+�V�sxto�&�L����/�|�g�󋂿�uK�N���i�V�|#+���.�3P|q������Hi�B��.0ޒ���sÓ�{D-����R7�d'�c��
==�!�7�X�ٚ�o��\;>��c�i��%�;}>�)������p��@G?7?���-X��f����Q�N��bٱmR~�¥f8 E�����2"
���R%�q���3h��q�G��=]gb�sА��i����l�$�o�ٱ�3�^�J�qT�6��gtơ�m�?)�.�����ި���ߖ��a�@�돵�'�h�0��HO%�"c�LY}��Q���O���fWO�蠠�좰��)+��Ȍ�is��V�����Y�Y�O�@�h'����8��h��;��D���(-�g�s/�h	tT� �-�	����������AJ�sNU��3x�Z`��
�jߘ������E�S��ng�U�����s[j��?So\�%��"����*������ ������&�>�4x�H�.(q�zxR�\BV�n/�G�X
��O�� 7q�X
g"p��B�\ݶf��XY �Ӱ+{��y�H�dx����<&�cM�i�f�7��m�\KF��,ǎd�0Q;�vk��)�15Ps��ٕ����G��Ff�L<B}\����%�m��c�?�1�-��C޳6�qZ6�X��S(Y��8��@��)�}鯕V���� =�]���=޺9�]&�Fر��F�b�/�ߣ�%1���}8���&���<��i	������4�B;W�:��B~u15��}��\�|ۂ��T���+�	 Z\?��!��+��W o��;7!�6�i�<��vdyI���_�z�S#F����c�f�ڜ3K�y��_�عhǍ�C�Z��9��v���!���ƶ(�H�*�b�L��:����w(�XXZ����]7 ��q�\�m)d/�^6�S{����s"4�4�sbTE��6���j�X�"�a�k`�_�M�Lʸ�j Ki �;+T�n�N�x���_Lz���tDw�� �*�aL8��7o�"P�s��0PF���ʴf�B��q0}���#���(�3G2��S��(�Ҁ �%߄�qH�, a�7�F\�R���Ҕ�Jj��*�������Yp���x�S��?`v_��kA	@�S"Ƃ�5&#3kH���Y�b*��,�]QB�i�B�:���i~��B߂·�l�p&>����`ȶ�ɢqN�61����"����Q�^�~��o/��M9�G��~>���ϖ�Igm�y�9@�}Ԫ�Q��n-��Z�bTP\���Sň�dَ�۴��O@`�]%&ծ��4RQK�2���<1/��[e�3#��
�����@��yK���l�����=}��;q�3R_��d��ؙc�����jK�:�i����q*�E\<nS��%ʽ�;0'�D�o1�U�}���vÔ��q1LI33#0�k`����V�~YW�v�����2��*��"_���ՑC*_ZUGg��bH����E=a�沒F�qw�A�!��y�}C0�X*R�d7�,��7.{�����}����?�8fF���
}E�KNtڏPyp���g�l���#F1N�N�>���Q/TZշjw�S�%p�&N����
��XO^dK"4}�
�"1��&?�e��4��wj��#A�~��C��a�C֖E`zX�y��>���j;s��"W�7�#Om�t[vu��m$ˍ~��j���DWJ�B�A=�9_:�j�����j���`9�5V3�D{ϐ)�/�dn�X:�,d�s��MI�����dY~M��-�G���వ� e�QIX\�`G�nI3�á����9j>@�q�8����\[�#,pV�