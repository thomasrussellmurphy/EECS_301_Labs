��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>%��}w�K�.�TfxJT��1!�J]>�Pv]�5C��7�T��	�M��X��<��T��PK�)�0�Q��*H�J����04.<5_�x����'��̧��b�^`���D�����%��1��m��a�t�[�ֶ�|�MDnՍ�f���`k�P��Q�8���"L��c�A�]�r��d��ƕpիS��뗤h\��x���l���F���ƗK�a��0��ڟ�ƴ�r�K�a�ϣ�ᭀG�CQ�7����|��~ S!����tDL��)���C�Wu*;0��6�����2�@u¬�4�B{-"F�k���{̴	�Z%���#��}��
�k��7Noa��?h�tz|.��"ĝ»zB%q_�JP��!R���>�1��F������@kn��]ޗ:�^���{Ya��b��	%2�e�lw\��@��8�����L���K����\��+�^f?-��3G.���:�H6G�����ָFb�s�x$���Yt�+y�Z�Aq�p/WZ¥/�(j��RU�rJ>~�ִ����L�AK$��b�"ؔΪ�f���L:�jÃ[5l�\���v&B�ȡ�T�2��Hb&�tf��F����o��yDS&LE���B0�4M%����F"tR'�(r�#����o�B�� �� �* ��G�{��f,�������'W�ޓ�a�I^g<�ƾ����p�Q�
k�q�ĝ=-+}pD���	J0�a�4�~V%7#�j�����_7A���j��h�Z�"G�򮭔���f�,4��}A� �'�����r�ܱ�9��E �v g�C�q1gn��&.�i�9�!�~�h-�qE���7��n �A��E�C$+G�G�H)5F�����r"q8põ�;�^H��\V��ּB��4��]×��a}�M�S��Z�R��b�Z
�Z��|�.��mZ�1/1�������*P34F�9��s&x��3�$|Г�e��Y]�$v��@�L&|�����i��i��#-.�lV��	�{&qF�B�?(M4y��>�ڣ�R��&��)��Oa�#�n���9�α�`=wjje0��P��`<��01�3kc6��צ�;Xg�%ؐ�(CC��������0à��Z�HH�䛇RaE�+�p�5���Rj�VHy!o�Hzӑn�~�j~���QYbr�)����P�,���T���M��|A�2�iU(%O>�Nl@ȿ�kD}�j�zz�}@ow7�̈�mM�����<������P_AZm�dR�(
ZSmr�	Qo�|eg�S�ci�ARU-�b����P����O���֕B��gy�%�<וuHF?��˕g�2HnlL9�f��+����}gY5w���P�|���ɞ6y�%�v��'� �9R|���=��aNr�� ��a�����E��жܯ��v�6|"B�=5� ���j {�5nFY�[�S�Cu����Vb� WSy�ޭ�V�\�T��:vo�3��r �tv�kTcׂ�J����~�uG�M������@�Qe8/Y��؃",3�?̠��9mY����I_b�`��ޚ�_�g�;��߈��̑z���u)�`"UC��
Pi�R�u3v����n�c��W����4�`�a��~���n�o�w�=r<��T����2)2�r�AQ��-A�f����s�e����5{�?�xG��U,Fể�v����u�ư
�����<e�k����4ZW=���z���옿|�0=�kU˓�|U�Q��~M��>�E{S?�l���y�	�8a�M=��r�<��{ӈJ�%-?������ ��e�kkٺ\�>��Ʊ����?�Xxzsg��ܽdN��߷ގP�kv���.n���&�/�Q�F%ܰm5�W��U��[��<�����������N�
n����둥i�����.�����G�v��X�=�8#�E����`���WD�l�\�}B4�߿)��B��#	Pp���A���0I;���0���P/$���Z�����������7�=K���N��GA������Ϡ:�����m�#N�,6���/����Z�Y�-��"79�����nu�Mg�a}�-��u��X��f��v����r���6��,JZ�8�ud/k������.���}��<g̳:�b�rU�v�i��ׂ���`�٢�H��eM�Ӓ���u _�A�|]'�3��Ů�����{�>?��6����1��������ȅ�����k&�X��6	��'�	p���s���V��cX��,�����Ο��c��.�!�bI*ո6h�z�nkɃ�}7
���03i�B�2;�X�M	�;k�FY`7��q>z���2s>���}�@h�)B_B�t�1!]#_���#���7��݃Y���5a6zMl�b8D���E-o˲+'4p���ᩛ������9T�҃�n��%p�u؇Ðo��M��z���b��/��儆c�P�u[B�)s�Z�}ok���ɷ��s @��Y��
�` V�|כ75��R��
V=y4�1��W�#oD�T�$:V����H�d�ᶁc�p$� TW2��L"ߛ4��t��I3n<�d�.re�g�hw����(ֶi���|F��k�B�JtI�6v<o�h1�2�.i�c[�ɰRq��?����W��^#o�7k6AiX0}K1p�>{��ʡݩ�� �\2��76e���porS;r���+狷����&)17i�:p��!b,=�%�k�*���[s!�3nH�r�tQI��NH]Y]�� foU�tf���if��Q�|��~�s/�Z����dnK(�=<����l���k�e�B�/�f
]!u�,�X��������V��� ��TA@��5�j>{DdY��g¤�3�x]v7���a}�mQ�%�(�N��~�֊��G?5�_���i�3iɋ��f�L�,Uȫh�x�ϳS�����$%9�p?�S�
�UN��][�7�|��X�p�Nt�m͎bS�&� �P�� K�X'4.]I�"��b��,�\҄�v;�al�8�]�"���c�K}�m�p�6���a�7OXw�S"�����Q�L�]ñyN��A��%t]6�T�W:�]���!P>F�w������!j��Fȅ�PUl�Y�P�I����S����bG~"����iKF?ka͔p{F�5�U���c�@���y�&[���*��q�e���H���dp��o�>_tx8^9�س㆔D�Az�T3�R��Co]jL?��Ո���g$6�������/K�	�����ќSՋdR���>���C���c���b�*lv��b������,���R�*#h#��BG�,�mE
L���c��غ:�����q���LWK�ҏ��G��zQy#ޑ��|̛�~Ocȍz�����(ܧ�6�4P���Z�YЬ�a�'!�h��p�^��`$(��$�bޡU~2�l��X{�+Lȳ����푲�p��;�q53��+�NV\c�����>��w�qgB���t������4�܆����H��%�����C�
�/��� �w�ޮz�i�	�C;�E]8�
Hg��c�G�_�99Y@ǖ}�����ǉ�J�j�yRg���2'���H-喖�.�^mH4�ʕ~��"�h�v�{nB���u���'J���!��p��D��/��S)g�JIEX&T#c;�<مRI*Pў0=��jAo��|�t:��u��0f�yD���<��1�A�PO��ē�y���*��+`+He��H_�iFA&�5S��aܔ�:0� ����4JV3���v���}���CxE�A�ں��ǒߖ&��:�����A���7�|�8��,b�

~�Š��⏞�S�d�[��A"�@�|����t��RI�vnnt�f�5���%Mn+��ѥw�S�x_���E�����+��0f�U���s
�@�^������R�P�C�ڻZG�.e>��Yp7��a@�'�+J}U��-5⬑����Ao/:Ҹ9
Z_=og;�b�<4��}+�C���$p��0���m��Ig���A��aq񤧑O��a<L6nb�����uP�7�`�};F>"㸨�h����H�y��P�Iϭ	)�;�Wȍ+ ���kü�6�b��"᪴}(T\�s�cO�fYu��X-ob�Թ}HNu�!�8��L#F�]AtU��G��| �ϵ�^[p+� �)�O�����L	�l����}j�35d��")}9.�P ���������QX�78nn�;�����3�aC�	C��?��B��n�X<��E�8�p�$ًW;�Km��o������[4A��\��>�y$9}Kd<2K��y��z7�*�����2�\QY�:B�
@6����$ŧ�z1#�<ҏ��7(,�={�
@/�+��/n��0�!R�>:�B����K� %V�5�S�P"��4n���ܡ'��%�	�RX9vB��2,&]��	� |7��vj���aS`Q�G/��$͒�E)�ߑ�II���i��Zu� ��*a���iV�'Y�e��Cj���aZqw,s�J|�^��	It]v�aʿ��@!��c�)30nXJm���Y�������뷮�l�$v�K��E����ڬ;]�U�$�p���X�}Z�IQ�$*�E���%�4<�&��b/\��G�m�s�����l�Z�F&��<M�gAqy���,��?O!�����s�����4җ�&Mt���,V^�5J5!Ūs��(���u���A�[Ș�K5�#�g�+ih/�%��7g��F�6$F�I�ڋ��<����r�������Wkpn�TF�U
m/lXDA�U4�  �%/�n��g��Gz� w6C�.��`$�Ú�6q�YUDa�q*�(��P��O�-����{MN�뎄��ȼ;Q<�e�����|�}�ʜ��I]r��"<VW3[Y5�vK0���  #e���ȳ��,�t�ex�ܿ�$ٰ��W3�Wn���tK���Z`�i�!����)��@ u��+��8�7L��Kc�v�ݢ֨:�/i^8�h��8XA��_6f�ZHD1��g{����M�� �Nl	[?��0�a�D�@P�����1�G���벦��pٻQx75a�)�(�jh�zoa7M��0�r7���_�R?&T����"��/L�>����ئ���Lj�
k��k���ز��l��� _����ť��?2��AR��f���@h���#Q��=����3��#H>Xv%sC����E������ԇ�ӻ{�P��EDց&��Dm�H��Qa�F���G1�h�yl�Z��h�6��xy�%kt^u7�f,s�fEy��n��Z�Q�Ds���]LmSa[]GuZ���U�TZX�cR����D�����?��	U��l@_Z�pϝ���~�hǈ���"���3�i�����>�$�-c��<�������,�?��P��W�s�Em�v�d�<���Z	�w���i�%�ٮ�����å��h��5棚�����֢+��͂�x����>UŹq�.Vow�^��y��������L[�ԝ�ED{f�H�z�#s�O݆�$eV���*I���1�u,ρ]��nr��Y&�S�c�Ŧx��-�I'��H�:�C���G}�8j�c��X�Ov�˗�`yyy��x�0h	6��觇�q�+$a���@�W�I�}v��v�e�hV-�/�(Q믑 �ɞ'���� �;:�e ޝ!��p�vj��1�ƀ�����l���"�^��&3Z� Aa�,ԡ�$ˍ��,���q}��^����d��6�a�H�hO���D��I�k{���]��0H�N�yƷ�A�YV�Y�����7��S��J����6&R���c���FιV�������o-��4�������(e�{=�c
�\�N�@���_���ç��]�|��|"��6�)_�K1���S}UwFj�[2��hK�_I$`{C5�l���^�bc�J�9t�T(a+�{�u�8��~�?��(�qZ��5%�+X�W2zm����ï�|��`SE,����*`�lO��V��)YH~�r�!I�.�pig��I[�e|�Q�sl.�I\�U�4��	'��ư\;�f��[*.�!�jq��t��e�V�1���K��n��w���O�:��b�9L���Z���ax v5���*m���y�B�����*���%rC0���N1���N6���o��b��(z�RLh��i�R�ee�|����� y;��2{Ϥ�����	ƫ�9q�?m%r8p�i.רJ� i@�Q
�t�k���e>>���*�^��2xe�j�<�UU�������2}XU#3�i����ʟqk�@'����O�mk��.����B��!aԔ���>��:�������;��#����;��DԊG���>�U���
���H^�������٨�Y)I@T��@�\�b��b#�\9_l�l�BU9��F�cuUKG�`�*^1)�e��� ��� {��Q �P�#�,W�ƖG U%�Lh�-e��������ɘ�P$�O?%�������1����+$jԴ=���+�3t����o�j�m*m���`']�-����+��{��N�i.�����`��i��e땕���qƢ����*��캙�Z�=��JȂ����ehJ�H��)_�X�L$�֯�&��@bu^%>�D���@?�,�r|��$q��4���!򏷆dUfN�h�3Z����͜� �)�1Gv���|�+Y*�©�����9Oɫ��G�"�҆�qT���b6@_	䶿M܌�,�x�<�{(Ќ��D�����eV��£J:'I��B�Kp�Tq�7��9�K�
�F?�=�\h�`�(e�������FVxԭ{�w�������/UR��"NH[����J����- @΢��	T������zڽ�ǩ��'drYB�*H�'nu�T)��6�$[�%��Pn/
��.�Ԕ���H�0������N�vs�1M�"��/���V ,�����}�ʆ�o�4N��#Os�2�i�׋�����x.����W��#	c�͇�[�Q�RGĻ��Нp��#�)ω+h��C�i���myvvL۫0s��cZ\bJ��C7�5) ٶ�rF���w"���B�4��V������jH~*d$��:o�E�{ZHDAۿd�nT��~�&E�?�������+O�po����I��rO�恲B;��r��q�] ��F��I���<�����ɪ�:�m=�˥ev[,cχIB1��֨�?������fp��]0V�p� A�t�2���6\�,|�M@�k,@�)�e�⧝=9Nk'q��/팥I���R ����(�����0X�{�v���i�"z���4o!���f�r��lk��4@�y��;x�u�E~ I�AGKJX��b䫋f���Xk�$kx2�t� ڧ:A�����]��z�l��ġ��+����2� �x����<gM��5f��iw��qkJ���F ��į��n����H/J��f[KR�6]0�B�3���}"��O����wa?�u�(~H���t��b.��	�|2�s���"�,��չa~q��UE$�����	�u^�i��0�{6�T]�&P~���C;pn`��d�2|��1�j�7�	������<�/����J���E��QȐ�ϊ�����f���
:X��I�����}eXw��=[�@���(�u�.D_�<�>�l�8
�
�iFUT0��?���䍗P��!�P�\4��?7Qß��>~�\�M]�ʩ�^[������T�����A\��2��tL�m`� �R�0�	r��LO���C������&��]�P5=�O��ɫ��paV�|�H�n�8��{a���������I�a i92�������#����Q�|�u<�+E�
ǽ�I�Mk-g,��oj�vU��ܷm!O>��3m�����.e�]o�Fv��o�1�����I_,���;�B
#�0��۶4)}��s5h<�nw���c��U6?Ȕ �s$�!F \rd�������>)�t(��������ƹpK�D�>��R_���d������p$�Y��$��;7n�kɹS[�Y�Ij�1�ؗK��}
��~f�q���R��y8�� Q����� �9>�bd�F�l�<TY��~}�@6�����eCy�(jɽ��|4<r��SrO:��i�'���6\�ê7�sھ��m�w(�e�~�z��@DVe̡�?b�R����=�L��x�"�K��=�K���~�
�� ��YT�L�$�v�h�5څ���el#�N��&><��H4�`�>�"��Jt
�|B�^6�֔JZ���˵�X�Msi:���F{�a_v�v��
����j�|�:]azK�)���#��֒B}|����J|�P�5ei�O���oaz<�� ���_��z��	�ն6���z���2�V�ڭ{���}��̫������@�Ui�K<q�N�gZAA��N�s���"с�Չm7h��)�h��m��Td��=$��L!4�f�~�.*J�����,����e�o������x�d�������RV��l5c��G��1%UU�X��9ƺf�PR��V:�Jr�iBc��Sb���9ǩ�N?���^|�q�k���A*�w4���9#���u���!
�����q:��ɟŃt͡ʰi*�5�}H�7e�=��{��6�$�� ����y���b4��.m�j�P�~N����i(ݎ0�s��R�סM>�K)�o��v��&�T
3=65!Vڡr�������9�_���d�Y�����w�_��iz���I⭕�� �u�\�\�np���m�!	��/�g$%#��%,)��ˉ$�?ڈ_®z�W�}?1�9��l�" ��o(P�(xs��p�X|��VQ���]H����$1���(�9��:wy��-�J�����}�� �`vصM߻cnM�=��җ�@3|���Z�.���A��Vl(���J�B�4�p�']��NwX$7�
crT��7K�;���nnPq����LP7�8�t�M�tkL~H���_@n�{�	n哭J)�W2�9���	ȣ�l$�/�ʖ=ؘ�����O&gƞ��	�w��4R�d�n��!0�	6t������r�蜾	�,�qYe	h;�a�����XS����D,V���`�R@���\��EGW��3�"��4>|\+_�GȰ�]�/�����wQ��y�s�2p�,}=��" ���&�#���$��c��ͤ?h,�!C�}u;��(4\��uh�8�HGx�[�~�h~`>�Ӵ.� ׬��f]mH�z��` �(ϙ:�.����$� �H�� ������i��V��Iq�\���6� ���F���M�_���ȁ�o���*?�%4�廊�<o) ̵m#���$��Fd�J��/�k����:���
$�jͳ7`m�����&p (.Jg6�)j��G����j7���oUv�cl��x�Y��	6T�&�{�ߊ���X�``Eu�6�{\1.o����ʴ�,%�;C���R��ܶ%&u�Y�A�XzwH��~�r��o�{쐽�b��6h֩a4�9�@��'+�;��y��S)8m�R�k���12�����m	R��WA0�S ��`��<'~6�Z6���c�l|	���U�P/'Ȇ���;��8���i�ڋ���-C�(E�8$O������+�6B��xl#Dq>yV��$(1�|�l�q¶��jR3]8���� ū7�M*�?k(H�~��EI@��.�� ]ڎ����
�d>+�7s��t��Z�4�ĻH�xN�ɅP����}I�`�e��Q��繑q\/Q�e��c��P�ţ����]�HĮ���	��[h��Y��g���L�J��q���B�	M�PL�C�q�M�R"���K�o�d�[����f9K'V��L�e�5�_;-kS����k�;�YMRh3p�΋�!�A�b�G��`�P��V��ĥT��c�7n��3z(���%.��Q���������w��l����a�i,�ԑ�1mbʈ�3�w<6D	^��'H�(y�!m�K5pK��UiTCo/{�8x;�)��x����RY�Q��69��ʑ:��|��AlS�7�P��J-�e�):v���C�a/s�I��YR-���8ͷ�_�w"�B���C��������_���!���Zޛ��u���Ŗ���ߔ�P�̀qT���Ks�/R��g�;�/f+�Zx�b��9v#DIu��^K>���<���Czt�t�4q���h�6�Y%v����f�'���"'��+M��A��g�A'pB�۹�>�e�1���]h.�3�&j�c.��Y��p��XT�(`n=���g��\�pC0T�@x^Aa�J���u[�ꐁ�V3�I� �i�Gq��Tm=7�:�Z���rx�w���H�J.f_"j���ʴA��	��H��e���#6s3�뤜������!��-�k�B���T}��Ԣ7�%��z�'tީƻ�=(N�87�4̆滲�~���:����3��+<i��q�C/�4��0��?�g��}��w�%�π�GeM�xB���nQ��'�)�#m`�E1W k�f��ޮ�g+i�V�"�Z��2�-��F1*���%�^�]e�T�|���eM��g!��ѳ�Y��+O��r~�{�v�r��ׯ!�æɍ��5at���db�e��qu	����{�e���۽T7+���o�Vo�c*'�*��%�,T��'�Eɬl��89�$&~���Wq���M�&!b�q��$�m���!�����W��${Aݹ��ƼĆ�3�����D�B"F݅b�e��Q�m�4G>w�D�)�n�?�`���υ�k���5!�v,��������b�\"�"o����Kat	�|)ٮ�L�K=�k���'٧+�H��ͨe\���a<��K4���_��L�Z��dSӭ�	[�g��6[�3�\MQ5e$�v �����f��&��<��0�<���v 1�`�z o�8%��7��y~���>6��!]1&�p�%a�!�H% )E�T��=7!�x*�SF�5`��Ɇ�� -�u�@��@��e6~�o�D��3�����"������"�1+�x!�a���q|k�7ːst�=����Px#u0�e"�x��vˌ ��gf1��o�/�O��E��6@
������XǯF������.}��L�0{wV�D���z<O9��߶��NH�6ƬE J�-
mP���JsA�Q��T�dܵ