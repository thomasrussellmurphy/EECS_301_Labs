��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�i��a
Α1S%� �uj?�L�3��TLei-3^5]E�$���i3ϐ�''$�(ع+޼$���V'��?��J�?���.N�#�W.��c�~����il"�e�{Ā.j��N�(<��� �c�x-�\�u�Zqh��˞	6��4J�-^�.�e/��
�j�ΰ?lտxܑ��Өd���@8�{�ɮ���{6a�Ciw���h;���r8�3i�)����*���|���0��6�G&4ݔ�*�9a/YN�h�^��O�4Z/��׆��K�+�r;�����*��H�|5z P=9'���4��I��X�JR���%�x��25@,�CR�_��_ �v�j�gAF-Պ�8'��9.0�S}���J$����3����\�������A?��Hފ���Ϻ<����~^��a����������p�D���D6�L?��B8B
�����y�n8&�
ܙ��ϒ��������C}�Q�-��.��_7"b�f�S�f�8j������@]L�=��Tӂv�=��N$�՜���apF<�w�G(�S���k)����/m ����T������t��wŢ!�(����M� a,�t�j��o�E���_%͈Wr��g���U(���@���?b:����p%��#��

Y����l�2����97Q���p�p�����&��Z�į��`;3��諯�Zij����\�K�C����d�pA�1; ER�"j�������@8I�ƣ��wYm�Hl-���V��&�-�n<��Š���U ��/4ϳ���#"t��ﰜ���q��zŒl���M`�����C������o6�����L*DH@C��9S�Rn�9Q�ʀ�yt�D�A	�Gзn��u2E���+�4�IN�����@�<A]�5�T��*�E��G+pz��f��1ʋ ���hM��~��\=�ܧ�3Ly�ZkN�-F�L�c��G�� ��[��ۇ�S ��:Y[���fϢ��}�c<�5���������4�f�������A� �?X��K6S�`��Gڔ��%/�,?L\��5;<��ȏG�� ��N�۝ �l&��K �t��<��
�1��	�x��P}�_�$}U槚sP��ܱ�Dv	kgc����vf����V�\��p}��Y�y�������H��X6�u�ѺR>�[���d����͆1o�/A[�T��fF������$��A��K��P�IK�e�e��첷c$�A� =��ԳxS��h֚����0�F#b-��ϐ�$f�7�Հ�Xny�|�C������Om���ၢ���̜;!�H�L�N<�}.�vO�������Li8��(B��KG���O��r!kr�kt���֭���z[l��M����RC��~sE�Y��B�����Њ��|I/R�Wn�Ԡ5�uv_���r!Sv�Grn�L��lkq^���!
���'�)[�Wk �H%��#���%4G�2����8!o.�jP�r���Y1����p$�VCSȃ����6��/0`N �$o<D�K�,u��n���Ɇ�ޠ��9w]�E2�E���b�1[���.����P4:�v� �S|�����u|��D���q�3��oeWK|x�3��E��Z,[X2r���͘^��J�Sc����ǲ���
���R+{J:��rvii5m�"_���J��k��8� ?���y��H����J���'N�bU���� ����jR�H�<"��A(;�V�2�ůd(�-/3S�n��	'5(~^��֖��ٝ��4��CNw�Ơ���v��Fb�lF�^,`H����A�7lK��sh������a�z��<�(Kʆ�����⛎&��"�j�,��2�d�gK����G���@��8��BTB����|;�j$`���?l@*-�ő�R�����7�˳.!�]d��!�9���d�v#��ƌ�ۥ�������j.zU͜#ů�V�J��/v�e�"̾=a�HМ������h���j�{��᪼B����t�XbV�|���Aû-�}�jûY���bK}�$H����խc3B�y�	K#�uB,smp�˞t��+R�^�CG��=�Y�h�3�	�;d?���{��y��xZF؈0��}kZ�A�����_�o�7���� BCDlVY���'��;��%��YT�9pqQ�ޝi���]�.��ۑ�gT�cn�?�J�,��ѝ�Jט��q �dߘX�s��!Vw����g�` z2r���⭷Ʋ�{T�,�%nP�j���+`�+Gbצ���RCG�5�4T���z?���<�Z��25�AN7a:�8��OT:O*>�n�g�����ަ���3A/�<6�s����T�� q���,p�:�5�h���ۛ8�����Ն�n�����pʛ� *�RT���Ex��P�(kv���$Pu4� ��)�b���%��4]\�Ըv܄�h+�<Z���߫������8.�ޝ��f޴䚍��v�;1G6=I�	�us��W�'Ii-=RMEv�D
=�Ǽ��]+\���1o�)����o�j~jZ�{#��K���2A��"ᯤ��2�w�7͹T���6)�cz0���S���2w��n`3�{)��xm��{��h�����ғFB�Z_����]��e��P�C55�T���� ���{k�U�Nd8�8XTx�u�+�Z���z�k�u߉�%��:�K`��r��9�検���~�*]�Wv���������#x���N��ã��p�𓬂��g���q���������A�6��=�v�m��L��Rh��.� ���9+JsWl�jn��t�&�l�쾋�}��ϐ�
�o�P�p;��T?<�e�/�`��0�r��S(��.���X�vMD��?8��񫗩k���gqI���g�b��)=��VHᓓ��@��z%mF�1�����;���k��R��d�
��/\��)�v��Z�Zk>~	�0@�m��l�a������h&z{�)��J�$ ��F0��f�$�P�ʿ�l���k����,<�q^����In�sAօ��l�f��j�-�,	�gEA���>b����9�y����TI��S�B0^u�R*�-���r��׮�v�N�Á�-�w� ј�J/}0zQRI��b���2l�p@]���Z�aSЗYɤ��q�
Z�����0�������l�A�{x�۬��1�9��(��t�9���R���Vd�����7!�d����-V�
QaR�+!��Jl���K� *��Y?�9/s�g���.�W5�[/b�wo-it�9gf�O
��A-�򊚗������F�ܶ]����[n��^ٞ�J���3#[���.p�N5/X�%��r"YZ����9�'�e,`J�]v�#�o}��c� /�1�6��裩�w�!�N��e��%|�z�5N}O~��>�2˃+П��o'�N�#�e���M�6���H�ShS��RL����L*!b�Ɩ*>.-Nb$_�*�O��!3�G���w��9�"m|i�������CoZ�Zv\lS�������w���������8$ٕ����~��J�a�����E2�W�/b� ��ھ)@�����#���}��BL_S�֦�l�ѥm���,��6EfG-=��qI2�wĸ.�
T𵇌C�=\I3�D�+�uqJa�^�&�=&����C/�\;�?�>2S�<9G�+B��Ω]�2n"mk��l���!�I)�'�_�1)�gn5��l렙�o+t�����>y%�6w�4���ߚ�k��c��������%b� ���D�/~��--H�6�޿��{�)�~4S�AA�=�ԃӨX׾����s-_ mr��Е��kxs-��1�U�����#��Ѳ��I�.E�4��|��D��u��r=m��0�x�+FF�����x��6��Dۃ�s-R�����>�I:�ѽ�$�M�ܛs�4��r�E½1�������O�����v9�38+$�oOo<]�x�,��ɫ�b�BM�g1�y>wW~-^��}j�h�,+.�r�iDΊ�
Z[��p֌�IE��Z�F|�į�e�o,)'�=f���2�B��k~I[�G��N
R��v�/�������Y1{�<���%�K��*	��9�;�@���B�g���p��L�|@���or�~�WX������(�b���!�X��V�"[�e!�J9���%k.�����:�ߊ�[���G�X,���E�H�%��=xZ�a�S�-��6i�8G�j2�Aқ��v���=�W��96��更�dt�����g�ʍ=�♄@6*2�;�N�C!�s�Ӝ*���*��
6��*�br^շ�g0�O�9���Z��&�h&�c±+t��"FX�$�Sj().z�\;�
�r��*�\yό�W���Aծ�A�aC�_x�X�ׇ�~7\�Ve^��gݱ:�m�΁�0i�"Rѕ��Q	~e4��7~^�m��+Vl������>����P�A�� �W���Lqaf\PTg)�g����]E-QY���q��]9��zq���9N��m7���{O`&�c�L����EG/z}^/-�f=G�PC[�����z��С�m���I�%����d��S`��\/��>����:���jj�G�w�A�E�(���ɋ�/��2_?�6C�1�|x�ҷ��������l���M��s�c�90���p�[�W ���v�ڐa�;�Q�����{2ҫ��G�2��yN/�d�j�j�ֱ8����6`!v��zBш�h����K̍�|!���b���
�q.8@��Ũ�OA�+����k�D�$�4� �.���4�hڂ�{g��4ն�Ĺ�N�Q�Y��N�P�}�Z�vO�Z x������b=W.�xĲo����bs�6}.�v݃��l����z�Š�#`P��^�ĕ4�S"X�y�q�K��q�Vi���P�<g��^��z��EF^%�-�/o���Z���F_��c�6F�=����,���v��{7BL������&��C7d ;M7	��&c{�����ѝ����X-=�Ш((���؞�9��/x"���,kII�o�RWU9l,��7�T��le}��x#
*i0D$=�G�K���%����#*b�xQ�fD�)�D��$�g�"���K�졺6��ǊU�:�p��n���7���
������E�s����6z�kӞ2�F�pu�4�D�߾��B<AJC����Zܟ��tO�5P���WϾ0�wmd�z�]�4:�;�X��||&\���e�U��"��MҌH%p�ֹP�ȩu�\��ȃ�`�IlPa��f�֐����!JA:�����n��-��y��1��A�TY��F~O�+9�
�a-a�������T�rAƅ��,g��a%�MH
�\X:�}p�@��y��#ޞ���E�.�|���ˊ�!42��b� �8mc�=d-f�cZ�k5
g�|@�fk��Fot�W��O�.��}Z�~�S��w�ף��p�����|Rҥ��,C�U<S~��~��Ո
U��hR�zYН��=���y�E���X5�af���v�4�D�%��6ofQ`ȵ�z�dB�&�T.��*\�t\�/�*�]y�2�a�D�PBXkeQ��;�����p0�f�+H�rE ��g�d��{x���Q]��7K�X���-�3�u�/�����&�����L�Uȴ[Y�2&Dg]6hH������Z9�t[})^"���F�P"8�U�3XC���������L���Sdajh�!#�8��	"�������6�g�d�Ml��ڶ��}��c�^⏻�s�UT;(�4~�Z�����y��2����!C�MY^�6��=W��Ć�����;�d�O�ꪘ��FO���s3y�x����"$�^SW�k�<��㺆���Z)��d!��K{|RX�/T��[%�c6��q~hQ������$�b�d��9yR����@.��?:�}J�/��p�6� �?>e}�!_x퉞�T����ADX���uO��:y�NJZVS��q�*�����<��q��8�K�/S�)B_�Ɠy�n�ϔ����4a��u�n�H��)i̽�+��m>�Dv��aUж4�W��k3��¤��:O�lf��^E�}�2IPE��������A]���.{�R��jq�	T N�+1�ev��F ,�k�.�n�ph����b��@�N�W'�1+ <`��#�w*��j��y$U㱰��T��}�.��X=U*�8�|b|����6}��b~�
�
��A�v �ܽ�$�=0�C�'��IAu�f<y@D:��"m�gO��K�3����,�)~��	���𧇘hȇ^V���6�Գ��$�E$�q�+��_�����ֵ̜V�
����d�
�rJX
㕃�n3�T���r���g�x��#��{p���I����2fV����e�W;�q�ֱ2�x��>��B��p��(��UjR�=^�ܭ��p��H���tW�|�TE���9�^�����r /���C1t,�V�� E��bvWPu��{����_���������i�Z[H�+���DSՌ����`\7K�q�!ҥ�{܃�����#�3�T=�e^6�:�t��X<%��^Ԩ�P�r�����ΑD7���V1jn.x�Z�^�	�O_�L%�Td���((�m���熬�3�����G�a���+y�M¬���U=&\�V����/
�ܛg3'ǋ�G�ԏ)�IK�|�Lg�{M�G�DD��Զ���l;E�~G�F�)�S9�+`G�RSTQ�7f�*,��#�<��G��B+���{B�E�0n;��&�9�� �,\�t�9ܚt�7y���6�$�� ����_�O�0 ��^dt����e�{�5~�$�W���"�e�W�0%cv~Mm�j��1w|�=j3bt�b,�AE��	o�6��z<�,%�\����#�����(A���<�{�����g�|�}�/���2�*�L��_d-,�M�*�	���6K��э =go2������<lw+
�CZo/{�%D�B�|��xdyn��TS?���l��y�ƛƹVʦ]����<d>>���s�Y��G�X�[����wNK���I4P�.�9E⠕�iQ��6���DH��tC|UP�$���ڦw�+�~+���ѦZ�.>�LK#�,h��6��~2�Dvi!���?R��U4$�E����'� X�A�S�����̺���OF�!�JC�Z+�չ�X<Tg�0gz����U�g�	��kc��<�?�ΜU���EÙ�O�!��C��/|��F�?,�z!Օi��=0=�")d��кVHMN��r��f��z�0ƞ���)H��e���2���E�'�0���3q�|Z1�.d1@�.Nf���ഞZ�8X-����K#�.���Y�1��O��?�֦���DW:�Tzsv��c���}6>z���.�=�`e�����⼈ަ�RV� �����������������^ߟq�W�����3��ku.��4o�cL`���c4#k5	�<� k�;�zC�+9l��ZFP P�3�~O��Tco���B39Y�#�u���~QL�!�R������(�2���w��5M�}7� ����g��U�͜$�P�܎��%H2O���*V���9j��qk�#�~kb@?��n#8�x�Z�Vc��J�o�-����knwY-��$���[�En��ɨ�\�������������>K->�:.�����/�AP�L"$Tl��<�:��A�r�2R�ó����-�fq
i�cE����)��)��Pw���B_4��������NS��fU[1���r1��f���x�}MWs9��MT��d��ạ�"i!��_d��I3/?��aJ-���e�m.�z�����#�g�oVDE��!gx��Cx��j?�>�Nv����=��yk4�m��̘�x�H/1H%olm���=�lz�>��/v�I��#��}�G�I&j�gg�]3QHT��[���<c��31Wm�P�$b�M������Cu��&�a�O��Ȇ���7�vR��ö- 2��Sݜ  ��A��6H�˂�YB���>[�<liE@��3�B���ڲ$o.��vh��v'����p�	u�>*]Qt _r`���Z��ED��d�;D��X܆�JPWC�M�$���[6D�.kjK�լ ��ht77f��D�y�$�l���K�ʣhګ��W��跺�Ԑƍvi04'瓟O%����g�KU9��K�D��W�\oo������,�@̻&ű?���f�a�J�	� ��,-O�=�^-���Ž�F�I��Y/r��2����[�S�`�kʑ��U��RD%���B������V�C���Z���T�3dd��(���ſ���u<�I��W��t�`����
���9�+����ePӬ����fS�.���Oi����)�=�>k�PsciBU~1�! W~5�2�6�S�ƺ�N�8G^|��]L���~^ϟ�vAt�A]s[x��(�Sp��{4]�T���4:�|�k/� ��	�p&�(d�d$~ZŎ�������#;{,�$:��7Ev��W9�]t����(�<�G&9�3&��*;�T��.��=6��f�	��ryG�_�������Z����~�C�4�v&T���6-��d�"wa#(�߰7�-�:�d�$���Q�c�;:qt�\��&����U�4�Y#{W�iT��<�Qd�X2�K8��rt�eXkØ~�wp�����,�k������s��� e(_GDv�%+z'w�Đ:��|�O��H�7Yf.<!�����q
���U&�ոwqX���|��S>�����g�uxj�h]#ˢf`l0]���B��R�1UP'e��Mlx�o�O� <��prd,gg��C>,�d�{���SޠFG����yR��D)�d��K �vج�8� �@�V�Ԃ��r�hPo���{��tY�Y��f׵�jT�_��S��Q)�]����$q�a�+N�|.�|�?�[f�G�
�n��"u��W|t�����Iwu!��L'5ݥ�m)��m��BC�3�|�������; O@��ע���7�"֦�zC�� c����O%�A�L¸Xi;���<I�W���RZ ^�q�F+gҥgU>Z2B׀���1��հ�d���DGYXLܠ�����a�ky.
߬�W�c� ����T��?Tk9[+���8��׉koL�du
1�2��嗩5�u��w!�:�T0���/�	�d�98��Y�Lծ�T)df�/\��lt�|�y���a�G<��A�&��D�a����6���2��p�@���q���h�*�f=��W�\R�&�
�d�`L�R3.�$+7�q��/�e�DT���Ț�X���"�#Z�!5d>����V�ԠH<�ͯ3����e�:o}��L3���(�2z&���Z������ob
�M�w����qlH�8�#�
��8tݷm�)/�>u/�	�4s���'UN�p� �82�ዃ�g��p�eP�ǐ�o�m��>���;Æ����g��=MxR�i�w
����t�	�7f��q<J�|��%�d�	�F��fg�ā��䢭n��2�ҹ�vDa#�?ɹ&4�	W̎3Q�S'�(egGT�,��~���Dc���Xɘ��QP��9^p.g��2F�"�������J;*%�S�����܏����&{���h���qD1k�)7CЊ�АlP��K��-�7�0���U3�ގ�9G�05�	�CԺT0���[{N-�b��q��"P�NB�T6/�CY�d;��&{��zGq�r��[�R�VU�X��T@�sh���G�H�?Ϫ@h�'LrQ�/�ns!,E�	x��:��J	���ZAl!0�����[�\�h*3��(	�ם��V�H]���`�)z���x3�*�hc�!7�[-\��v�A6���m�-I�-�l!���-T���pV�#:b�J[�����q�MO��U�x�X9����� {�;� :燬�9���t���ĺ�G���]��<�fK���n�������F�-%��h#c1�-2����
�����Y��_bd$vAu\���	d��` Z4�{nl���|�xҒ&%}7����	G�A�:v$��u�U驍��j힮S���ubZ�5[��K+rnh���nn��	Ul������������J|c����/�v�ߌ'��M�N�is�5�����:O�W)@C��A�&�|�7�)`�wg��W������;eǡO?�h}��5Ԧ�����R_���g��QF};/���Rݑ��Ŀ�r�iP[�N�Hܴ�T�����$���BF� n�V���Q*��
�rI���)�A]Y��P8��^��	������%����kc)����+)����K��IG�IPJ��a�RW���p� >g]]�4j���(7Q��c��g�7���؜��00��:��Č�`:pH�W����Nm����ު!��x� ��nGL��aq>��Çb�l�"F/kUH"b+/�-�K�i"^�Is�,��>��E�:����'�9ܼU���K��s���ʛ!I �����n�?>��$�0�9=����h�#�ǋ�_�-{�ѐ:K ��hx���>���W̞6s��Oh	�;Z2t�I���	?�w
v��aք��?��x%z6=	&m	!MX�-�ѤiS Q�Ŧy�\��L��Q�9�B9�ȑ�z�/CLf��)�o`Ө�)�y|�gF�쿩vA����?[��k��6G(�^4�;uF-=������i/E�Y,u�:�)%ze����jG�*-����i�f0<�8�����E���U������g��AT�k?{A\5k�s��1�����wf���Ǌ��W�{��Q=�pG~�_�A"�u�r �4.z��./�@Y ���F@�Ǎ��F��󩪭�c��5*�9�T#��
g�æ�~�m������a�|�o-���?qw���	��o����(Y��z�k��T�KY	*+�PW���	:�N�A=z(Y_�BLO����X�襪ģ�PtR�C�lR�a���/��z=ζ��h�%�ef���L�)JX �xZې"cp�1٨?����H���b��c�Xq��9sS�PⱮ�n�h��$�;���mGűz��/	���Ż^��O���6�z��!h���,���I:s�������c5xۣM����TGx0)Ac�%���T���i�ȦP���;w��P��"$l�5����ؖ�63�U3�=n3^i(��P�𣶱�\<7͍ui�d�0:��P���B8��r�϶�n��a�t�͸�<F��߿jԡS'�<~ZO7U�~�	v��JeC��T
Db�c�� �?PT+TtCAr����g��x�]GE,�Ts���?�D�n�ԇ}��%o����h+��ځo|1z	F��꾔	�m;��Cg(
����3�"�FST7^>�4��5�ZA�R��O�5��Ԛ��xsa��e�mG���S6J[��O�#�\^Es�W�)I.�C��F=!��)1�Z<�$�Pke����v���&0�U��V��Ya^��2��ٌM�?C�j�S1)��=Y�#�(�_�~�X�Ğ���n���a��O�z(<t}�k�Tv{���]O�g[�
p���v��jS���x�IT��}n����D|�d�4��y:,B�TY�p�^�����;�,�J�?���K��D�%j��AU,\�!�����C�*bV���n�b��үq�z��f�řT�
ҝ���9��n�iV��{bY����=��;�h��@@�4�S�Pqny0�۱1�GbI��R����#, �xiA����/J�ӗ�[7����߈kܷ�ڢߜG��%.�O�+���� aH�WoOB��j��8U�Z߿l�ʽ8�.؂�%�2�-n�����u�#pZ<��5y���#�\�)�f#��0S�u��H��T͚]�&Y��+yYp��jRaW3�3�@!�j�v�t ���3��kEŃ6ݼ�H��F���U�N�`�JL��ak�	n�N���2:�/r]z������Zbr�CA�w냳�"J�I�H]�z!1����s�,��(�g�e*���:zt�7��I�L8}����(jP�v
̢`�ٽTJO�B�^�^���9.[z3RR>fM=�$E�/� ��
QOP�[��?[�z����Z�~�5�_���!*8�P�7��)��*��) ��k����iS���whb��pL�P����0Y�f�0�/����	��k"���5!\�0W�������NҼyL:�8�M2�E��@�\��Ő��3������6g
X����ƣwƋ8�6y���B6J�2��u(Y�;iG
��������%f��o��q�\�M�Wbb%���7��$��s�>>�M��>�*4���XU4t�1��������;_�#MM&�|kN�����G�):ɰc��
��R]ժ^�x�t燶���E��?�t,y@Yd9
��u�R����$�����5'j�b�X��e�[�L��&�ς�FM.t�|��I�ɲ6�%�*7N"LU�$.�?�̶�ş ���O�v�oq�Jؾ7�Pq�*J�d뫷(LHmF��n�b񒢮�R$��Y3JW2��
*�j|��� �W��c-]���1��670"%��Ԥ�����f�%-�y�� Qԓ[|z�i"J���\:}�-(��Οx���]�O)��9����IݪyA�.�,�u�v������'��2��ku ��fF%���P$l4{���>�S=�&7&��{c�`ίWN%Py�m�̹�]����(�e+?eNx)j}P^}N3� O��L�͵Y�<
����-�i�k��J2��alH�i>T3H�3v!dN������{�l�^1�� ���(t�+�w�+�f��;N��>ȟ�K�w�e��)�օ��V'b��(��n�����"��Ӱ�ǐ�6��q@Z=;M�S�>mrŻD#��*�:L_T��\��l-� /g��mی�d�v�=�%��Na�{Ko�������L2a��_��)��w�9�/=�����h*T��`�7t%��аXW1h��(r[�� Z��v���ҒB��M�3��7J*�%�Ar8��:����iy�K4H�y|<��l}&P�zo�R�!j�����۾�W��@�C��+r�:����P���e=��,��!�u1�g�[�1�I���p�v��cV�׌%��e���u!c�7ze���Y�,|�k�֟Ci�/s]�5��)�3�z0D%��G���@�Ux�M4^[��V Ӫ�#II�k��0G]r�i�}��ts��ss:��-�G���]�5��t�� h���Ħ\KF�A��O���)��3GaZ��mւ��{?m(�.��1]���U�3/�6�7��\>�LÎ䉆*ĺ���B
:���r7BQ����'m"�bi��UN�@d@7��:�A�t7zgw�@��˶���sѺ�\I��Eu�!�q-x��x��Ԕ�s��Gf�;�;i��t� XCDia/%��~{�_�fI�=�M�T��^EƯ4A5\�e~�Yk~�����1E�B��.���+�����1<�9(�����
���q��8�m�Q���ȈXrkW��ҡ6��E��5�R�����g�Bng!���x ?��xce7V~���|~�T�&7!���ቝ8���#�h�<�k1q��r�-�y]1��w!z�p���	\���zO6� ��u)��b�+6�ٺav5���@�o�-5�U��2�Ql�`�7z�E}EB��AU�Eq-7�F,�b+��KG!B ���o�R�5��:Z�%�=F��EǄ��(��"���"���uO;��x���T�b���D��<{T9HǼ��9C�Cڠ7�pyc�2��6҄gN��X��ǝhFZ��<֜��|����tL����s�ɸ�i�і̹��k?��ڿs�\��R�A��X=eI�ʺ��>�U����/ژ�z�q�b��^R
�o,�h]�ӜU���#���t����))
n��rE�� Lo�ݣ���b�	(����^C��/�2w<���"��9�u�"��Ԥ&g�/@�����z���G}b��!d�Îa5�^��y��_���2{Jr��ׄ��2�6B-"�̣�k�5��R���	ξ�㉾�0i� V�4��L/��y1�$M��K�8����
��_��j�s{����:��v#���a���V�߻1�$C�����Q�?lR�v�!� 2���6�Ϯ��&�V\�����<ט���(eZ��g��L�=ٟ�l��#�z�8��ܳ�bh�[��l��*s��O �s6�@&I��֙6��l�_{x^�W�9Vf��1h������k>�@2��r^����M8�4�+>�Z��qXI꒧٨#A���6�0�c�����4�yr{�e��1�+d7"��u<�ZE�u�+��Zp����k8�dR��}�+�E��mP��2�-¹6�EB�	 {�Mj-�ݟY����ͳ#���/Ic V�_���M�ѝ��o�T��HEіh���";���R�)?��G��z�:_��5���&Z|�U����/�)�������Y�m��D��|�!I2K�*�m�פ�Z+����Q�7�=�:3���m�:��X�t�Z[8��jk���m!ei.����
��wSU��[CV��Er�J�c�V��ؑ����YV~Brk��F����� -Mh�<S߲��ڄ� �fV{�}5r�H�gVY�QM���}�/M��}[�L���Ww��g�7{�T5��;w�Y<1��wu�	,p/�В<(q���38:>������V��8�N��	+\f���1\�g_8� �}�8�P���%-|*�⎖+�f*Vd��"�c�kn���Ӣqa���W�բfi������W���{�l�D|[S������.Ɓֱ)?\@�����f����6Y���{^�7�f�Ȣ*hU������)�J�a Q:xfTL�I�f�~؍�:�X��2�NcN����1��Ԩ�|��P���Q7~��zt��f�Nk~�q#��pe�������t�Uߙ�Je��!���m}<�H�w�cN�JT�WY��5q1�ŗ_��>�1���`@�2l��C�~�Ȏ�z}b0�I����5��C���
5��d7	���V��=ɵ���T[��*�s�7��a���T2���vO�Įj_ݒ��U�yo��|Tm�Օ�Z	m�I�[#X����3w�A�����@C�¡��8��l��y�u
�K��8��^x�R�_��O����,��"��>8�(T���M�B�`>�X{�K''k̝ 6�m	�]N�^?��v>O�^X@�A�ؤ� mX ڜ�O��LsCJF�&C��	�AVn�z�k�6�%E:�W�dЈE*k��)y��hwT�o��,%HQV�t"�p�q��#(�É��j�@	!цt�^!s�u�"H�m�W��H �m�}���hj���\���G�n��I�+׮)9�d�9@")S>�23z�-1m�����`6�bT�8ȵv��*H
�N�������G���:��*�����o�_�OzQT�k�>V+ ��˖x�qf�3gZ�{[����2�;�p�mw����R��F�0J��E[��wF&B���9F���禸&gBa	xȫ�~��.E���O��3����sf�!@��wrn�3�]�쨦�a��xEd�UC&�/=ܶ�ъ��Թ� ������|�3T�^��w�ᆡ���������i�FQvU���g�5��!yz��$��
��o�Q����N/�/!<Yd�;:FP�I��@l�ǃfd��n�r���7�?��b�ɿo��� ��b�#�Tg7]z��7;�H�}��-��±�(�W�-��ƛ`�C�>��*";�'�1L0�+�sB�F=zZ��~�$,l�I{�X
��@L$�\���LR'�Hc�\�"�E+2�mG5�aY4ǎҗ��jse;f4+�B8�p���\3�W�Zˤ�a$x9��O|�$N��ٟ�I� 	1mI�䑰ن��VV��EqF�{�a�2�^(��%����������	���������m�Jt:'�̼���6�%??��'��u3�TN���7�'{�k܉`�Q"��s�d��M��W�PZ��'.R0�F+V���t̹}M�*#f2Õ�� jw�\��N��?������GY�cvx,�;wB � Y+��"��Kt��(�t������]�_J�C� ��i�V���07��VQc'_�V�t5�+��B7�A\+��Y��m��WA
hf�3LV����y��]�C�U��!�b;���8A;�d�O���Y4�d��4a7r��a����n�>;�f�8e8/G���5�^@m�T3b���i��͏���$K����ѥ�$d:"�s)����>�߬uĨwk%L��Qi�94�������e����f~�z ������L\&D�%�d8�R(��M���,׋��9tV(G�!�Hǌ��S�i���^'x�DB�:���D�]���՞�t�
C�2�-3?�H�x��麐O]���.c�$�h���Sh1�'��^���� (���3]}2���,�	����+f��F�1Y�`��!7C#����Ѳ9�n>W"5%��0/����s��kP�f��Pf�VYڝ0�iU�h܁��U¥d,ft�UpD��w���Ɓu)UR��Ȓ���>2�+I+�j�EY#��N<�Lg?fGdEIz�6���FC�~S�r��ff_ `��S�w�<<���ſ�LhE[1�B~���Ņd��y\B:�k��%�H)|_���Zw���XTБ���_)|����P��|�~Y�����������c���F�꧈������$d�B��׭
�!�m�^s�|�LZbi>��`fj���i��P#�ɘV�֍bSì��I8���P���Ш�h˯��0�0S�xB��8�b��%sK��7� ����K�~��nP�X­��5�_�D��G-@h�I����R�^���z=V��<�'�F�u#`�^˨hc�Ѻ��u�p�Z���e���;�q��4�yS��a��	ue���!w��+T� 0�_��2;[jq�_۔����*i�T��.|ʒ�K����O�ԅAjP��őI��4���o��z�!�T��$%��7�/������+���x��`��
��A���Q@F��m�c�����+��I��q�߿����k0ڳ���Lf���3$_�V���K�DMJ6�8]��G:�}/{��4/L�;�=Y�Ǳׅ����s�6@�Z��♙�S�h�s�!�給	b�z�k�!?Aд�.�.;3� �6���T����fOZ�;���!����*?o���U{$�E����,�sԘ���,�&�CAp%�T�.��a���6�m��R��L/ӋQBjD���Z6����Az�u}\^��q��"q#��-�I�i�幡��Y�O0�&dU�6��1�$����t�km����F1��}�Q�2e"�\�٥LA��7���8sI�j=#��J����t� �\qEx��e��m�G'�9Z�w�M �Q8�C�bʤ�.}ǧ)��o��� ��r(����V���젫�H�XKـ���,w%.5�#�NJ�%����*<�#��?� iP?)9zH���g�n~����_؉�/��񂪎dOi�H�)���s:!��Kh��?��J�����A�6'CL+�,���Y���D��"�p?�I�B?��,u::���h�V�O�4Q�#�k/e9 �����/��|�����@�S8��Opc'_9Ke�)��ESV*�WƑ����U�q��
$���_2���ȩ?a��n��BD�V	����]RX�<m����A=J���̻8���/:�3T��y;�L"�Y6������ݼ�����f&ܶ"��PT���j߄�3�e�bx�l���ʛ%D�G��2q�#//��q�����O����]��x%]n�x�U �B �G%KҞ �o�G�飝̹c7�	�FY����2�-*�\,j /�p�ˌ�3v^<"��c�[@A&�Y�=d���L3�W���#B]O��F���Y��Dc����8��ĉ��~N�X�N(��u��6r���G*��	!�����A6�|U�Y�4�?�I�R���(|k��s֝nM�.�NȻ�ѯ�X�7��4�D�g��`J��\�\���W�4α��lG�j�S�o�e���Bdr�K$ё�*�tౣXq��W0g��"}!)6[�bG����$��-�����71L��Q��ɺ���z4�_�;��_�B��t����j�vl���l����n�s�R�ht!n[ ��,�4&���g�	�d�=��ϱX)�*{k̎[�N�.ѱ�BK��v_D�9H_ך�)`�h�<�N��xy�%��~��$N|��)�"���8Np������xЗ��ە*nӘ����;_yu�ک|<��I)�hV.�hfmG�ξ��^�����KIX�{W�OV$R�+g��4�U�7�o �%85Ys���&/th���m{���Y[VMyf?�
H�{��k<�pA!~�.�sv�D�l�������e�y@ә5R�������"�1Y��Dl�j&����s��8An�"��f>�A�WAN+��H/vIPNr� �d^M���e[�G���|W+�l�R�l3�2���M���!G��>��l�/����W�,��,^���H��+
�`d��x1ٟ��a]�G>�?=�j둪:m�$��!�t�N�.*\k�~mS�7h���jr�ƹg`M��ܙa�q�59m�����2����T5��v ��J�I���v���l��!H��\B�-~�G?Q�� H����f>��[��L =�1X}�,]`l��3�#��T��!���e�[b���6�=6q�N.���\�b�����vw.�}h��73�y`��y�� �t.�u�񉜄���%P,�����Tj��ti"��X����e�W��m����������<�	�A�*���9Ø�eo6������ܰ_��p��b2Ւ�$)�q��U�,�R�(�`Vũ�T��ޚ�@Z���� GJd9;uRB�τ.��ٚa���4��D��XԬ�!w�_Zk��.��i������Iwњ���H��M�^j�o5;}$�}���a/mqcR�K���-�@*'��S,:��̭���b�b���74���O'z1���ݣ(��*�iws�Hi�Q@W�&M����I�:3����:���¹��G����=kY:�n����=xa�Os��'���&68T�t�]�IF�8��
���w%Rsr���Ϯ����%�rn#,W��&��.T �2��r�Mչ��R���20� GC�U�#j_���N�+YA,���.��}p��u���M�so�Jw$��F4-�v�7��ś�l���JD�#7n�:�׉�1R����,[%ֲ�Ύ���Q׸�G���1���ǂol�p;�	[h�1��}{�l��;*��4�Ϭ}tW*�(eGȠ��y��kY�h��`�>����W���x��߫�ք�A���M�~�s��Ѡ���hp�'xJ����/���st�l奷Ma%�G&��QR�<�,7H�N�2��g�&�/����g�h5ؾj(�a�N��m���ۦۚ��E�4r�����ޞ��@��{���Ҽ�J`�2�~{a���!�ܘ��JQ%���Ӌ�W6�Ťr:��Ns�U�[�L��$�u���]gQ�"�EcD��x��3㒳+!��&=b��$ľE�)`0�����V�����\�b?��d.�7�$�+�UF�\6����f�q"�������M�gY�����U��d�je�K@d�%,��gW%��~�Q4���ن�A�@}գ��$�
wGg�Tǐ���&�6y�T�l%wrͷX�v�51�!V�8!K�߆1ܺ��߼,�`E��Y�����k���4Zs��W�b����'�3�)C��h�YS�[�z�O�V�0�[́ıT��UR�}T�o2A�Qe�������h��H��gέ�w��}1$�����[P7��"��$�-r[��ԐJ׈����1��^��wD�4���"�{rv|I��q2 �1�0��N�CP��lT�i�K���ۋ
4t)_�g�H)t�A���1Di�.���J-唀�{�'��B�[{�3�����ȳ�(6���僭0=pHծ5#�F��)� D��o*\�c@,�d�n��|�"J�μ3�"�����5Ϊ?�)��-�]0�2n���v;��K�տW���}���T6�(|�iV&Y2m�ܪ�Z�R�|��ܝ�p
��&qFܨ�&�.����/=@"���S�i��.�D��T��=�_}�&Mn?$h�
nF���ץ!��p3�nХ�=*SL�􋺖�d�#cqͲ�j|"ahw�͜s�/\m���D�5"��f.�^P��)��[>?�=_9{�]/2|�������!|��� ����|&S`q³��՝o����Μ6��u8b(c��Fe Le ʬ&O��!�%<�NʢK����0���Y$����醋Q��p��M�F�!H&m�;-�ï�u���R�6�	}Dn��)[����f�V��5�d�1ex+��E�c�#Jg>u�s4��y��'�F�bw;�X�ATE�)�S+Pq�J��h��ڢ>�n���=���g��.�DQ�Y�R���e�<Ú5���x�/��;V>@�H�t�5�D}نgv4\�=F�*S2f��=L1LpT�u�.ʘ�l��<O,�T;����ٹf߬�zX
+�R!�+/#:E�3����5��0s�.+��~o0*�L&<��>�����q��'ր�Qs��xqy^��n�˚����k�3�"?�\a�ʈ�e�I��M:��B�x�2�9֧��Cn��Wb�T?�1!T&pax�F���_�3R�i���
ֻ�?-ea�
u߃�7�˙,Z���E��|�O'eeB��ĵ2�pw0�Xn���8�� nG�Г� `�"�F�<K+"�d��u�dx[#�W���V4�W�_���i�8>���tj�`U�<$��J�F*=��ֺY���q���5�Կd�.���w������
m,T��pF$�>��}TM��-�j�:�ñ�y]�B�������@�� �8���ju���`9�i��H(B6_ ��GHP�Wk���k*�G?�^��@E)��	'�0�*<�:��7�%׮Q����q^��?���N����>�A/�Q��p���oN._�oƍ�8z�`+)ť��[B��G�'���b��o��$}i�����9�~ϡZ"����0Q��yJ�V�<�_����l}e�o<��~B+��>���Hl]�ɼ'U�o�FVK�h<��b�����-Nߗ_2�����p����z�P�"`/d/W@�_�����zLP�`�7����!3|�#P�tլ��*@����uƪ��+�@7�*�J�4���S����q�3wA����r��ƭY�DY�4T��� ��M����$e�P�kE3�_[�)'5f�lau�#9��c�\�p��K���� �Ƃ0ᮇ)�A����٢�ibbd�"�Γ��E|"�CqIY����P1uH+'��Dd�<-*{���R���fNA�6���gI�WҞ�Vg�Fp',��8�5&S.��e���c��Y�D%�f�4Ǌ�Tx����^��2�_���h�c�wn�q_����n2��9�������I�y��i7���;��M̈�������~M��#`�L;�+ЖRX������A˼g]�CRѫ^
��&8E�؟�,�Zf!��`�t+�y�YL�DT�+���k��xs�����S�J�o�G3? U��Cl��,�ߠ�����lka���
�D��|��َ�>zd�G��.�Z��̽e�(�N��-��ˡ��z$�p��W��[�D��H���%���Zh<�M����!�3!���V�j��_��μQ����܌J�"%C"��x��nt��`��'�:���!j&n6��y�sBm��6�N%��ʂ��DK�A;C�)J�4� �f��8@���7A���r�82U섍|���3�$�fN��J������ ���6Һ��~�W���H��q�{�_U�L��N�4/�ø�j�ff �lY���}���8���E�_X/ަ��]�˖��]]ܳ�	�dh����$�Ķ����z�� �,x|ߜ��MY(o�;�_�O����k0
CY2}�ٱ�'ML�V��1"I�x���T�R�-L�Z�ES|E���m�;U��P�9�^?S�C�=V��S��g2@\/��񮡑�&C)!�I�]�������M���y J��8}F���"�2Z���ck�FqF�{^3�SL��D�9��9��(��Pfc�#I �H�p�i=|-u�(�Ȫ���߹�.���Wn����i� Og��kyh:K��Sޔ�a&��Q/W��,B�oyhJ��-�/gq^��L�AIV�)Qg/�d�ϑUU�OgY���wY��W�:<�@M

H|�1=*E�4��}֔��oEu��+[��D ��X�}5�2�C�	 ��i��� j��c+N)]�\��I�.6�k�i6�B]�$C��D\�-^/S�^��01�V��\��R �C�*��d[2ůN�T��4���,~8O�����~����(�+M�	|2���I���bY�1��G4b�衜����.�0ZU���$8���c1��B�\���Sxnd8YS�p��k��_X��iW�$�њ�o�e�XO
�AJ�cJM"fbOaE��<jE�X��D�{��5�F�	��tG�����O����A��]�x��^Й$���]6��� �����@M�m�@�^�w�Ii9�
s��J#��
�^�Z���W�qX]��E����=�Ӛ!!��f�I���M��cX[�#VcC`"������vxcB���_���R�08���?��T4RV��ŧ����E�ױ���4�&��AQMWt����P���f�_x�z�m�[� TA��$�g�r&�ų���`>�8}>���A�p;:>k����nԷGǦ^	�ե*�2 ��O쫷�����G�bH���*a#^�>��P(�2��@�v+�E��Z9���fn���j�̈n&�ӻl�n4�1�k6�9�|	U��&e�Ϝ��K[��J7�v�K�[	���V����s�ЛN�����≮� ľ>�<�� !��j--̴�;-������V�Hd+�c������Q�7ֻ�â�!3���/�j5&�`P�F�����O���z�����SF#M�i��4�=�����>ȣx8�� �s�[��!'���/���g�c��#���l�@]�����mPJ�y�g|Z�I�����M:�Y���>Յ�D	���p�y��̺��1`���	 ����^Vq\jH
��@�s8r�䎓I8.H�Ve��W���W��S���:�������3(;�=c�;�����<�8��=�@�St�<Hu_?���\y�L� ����4�{|���;d�!C�+F��V���P�����,��B(�JC�Z}ߩHF��_��ZǦP��EzS�G��a�J�v	�б#�~ �(�<�pc�Ҡ?�YC_ԣ��S�h�mh�"�e���GE�o���ގ}�孒)ٺy�B9�BO�>��Y��4i�L���l;*1)��\�Rž����/����O�ݢ)��w��P����l�B�S�vfoȆc�p�������{ ���&����v_�<�CreϢEp��D]:&�>")���`Q�%�_����`��7z�/�Qi��� �e �Q���^����9a����>���i�M����3��%j������7�Z�z|�hB�O�7��y���s��Uam�:@�LB����O4�J�{@n��ӌ0�
b[����b#����t&�(�8�Vŗ��������$�)�JGt�s�h����P�-n)1p�* ���?]�Nx�0��%��D�A+��SG(T�J��Ag�-�[� �'}ּk�$/��[,>���n���qb�&͡�>xo��id�mħ/�$#%/�f��j���e�:&͟������܈��SS 
���L¯[j�|�<_ �6B�	h�M�<��m�k���@Cw�Q���7l[e�ϒ�-o@=�C�D!N��kva68��ݢ����3� �����~{Y�u΁����+�hBG�r6�g.��I�t�r=��3� ��ԗ������:[q�+](a���W�
U�'�~D�Z�1�R4�9�nТ�,!w8���K��yN9���\
������
���=B��}��e��<�# I���d�O���^���qL���!9	��p�Pt����'��q�ǃ))?ZU{�Ւ�m�o�'�zA|�j�4�?��'��}�]Q~�������6�=��3F�����}mH�pp� �`��\\�Q�����\)��;$?mA.�!X��Z@2��r۫�,��޷���Y�i�}])a�w��9�{@$C~�E���`����~��d�������h5��Z���j��r/��<j�<!`�Ԋ�G�&I:�;)U�~�zp��逫K�@��m��OS:*Q�|ʿ�����Y���]�?��\�Pt��(�Ja���Z��W��o{'�ӂ���aU+,A�v,ī��-�sC[	"1�,��6d� N����&�ҁSy�~ՎdV��.����H�~����
7?��"��2�������L���8�O��N�%"ͱa��rhb����%
��ci3�z�dx�ړcMԨ������0Ӂ{��_��|W�XQ��(/��.7b��ƫ���5c� �"Ǿ_�,5)E��"��\0iљ�'��%P�]�����F�	����_��6�r6S���u�Zַ���iݫ?�~?z��=F�� e����#�P�}�E�B}���.e�L�Ayk@�� Ȱ�{V������j�v�x�5���{�o�\9ܭҲ��V��N��V�<g��"��Ŕ��T
�3���&ˍۓc�0)I"�
����{����lC�Vh�{5d�,�ut5��啻Qۧr�	��_��$����?,̹i�v�%��ƶ�L�M�@��@72l��.��Ac�%Ra�D��Ή��kԞ������@���ܒ٢���}�6��հj�Bf��|	C��G6��"����m��|�'h��*~Lm1��O8S���������Q+��7���[�:$6����qbJ�R!d���l�B}��Q���+*xP�ú�5�B����9�[0��4�>[Y��\�};ŅÂ�X�H9J�l~�֓��]P�����"ז҈������,�d>6���i�3w�� ���8�c� ��c��%�YQ�c9A}��>|�*���L�}A鸣���¸x��yό��M���Ƴ���Z@��]��*�}��sO[�%��|�S�A��x>
��-v#ӝ�F���= 	�W{E��VL��C��?�,�{��#�k94 $(y4�I��kr���	PK����Y!J�{�bj�T��U�?W�I��x�����;�
��݇�^:����xw��s��1����̗%���S��0Rk������n��F8?��Y��A�q�K�ZL�^��C����G��^�T-�㝈��&&���$���uY�_�����@7(p�~��=W:������R](`��Zl5:�������%�&me��<�6,;�mވijM[M�*P��3�C)yϨ�̬�t!	<kg��*�_����Ev��Ӥ5B�p~�펟JaS߰Q��E4�\�+������l�%�ƮBV�<�˼Z#�iĜ�W,{o%iN�U�LT�J�'M�2��:;_L D�Gļ��Vh������*E	�(���Q��3FTwr�,?{�h}2�a���>O���g�i�ʛ����|���+��"]
r�y�<
����n�����z-��� yt�"�Xʥ�^F޻���q��zn2R�B���iA6�[3O-�f��#�����a�Y����&c��I���7ȋQb�'�"K�os�;W)UlG!5�dE@Bє@%ݱ�#&Gu7/
�k�������X�Uek�ӹ� ��46����U��On�&@LA�x�Y8y�o��g�Dؔ���/����m���ڴ�o���k4eA�����}O#V%��P���b?��銾�h�{�C�ů�ტ��*����f�x8ݜP ����\p	6�9J���8)�U�Fs{�Fcq�G�ք�����3\:��ϞZ��y
��<0֎w��G�t�Dz��V%o�� '��'�a��`�Ê�����A{QD�����ΑH7g���v�6-��J���n���LHZg�k�l+��K�*/dv���a��t<M�q;��*nJ��ey��2dfVu�Ĵ���`�ޯ��L7��or�\����� ���S'Vk*�/l\?��������~t�R�7�Qo����H&nyhvTK�:'Cϼ��T�<Y�d��G~+�@�%r�\��JW����p����k"ҫ}'�L����#c�V����*e���*!"#��JviG��I�n����/�����X#Zg�=���v��pd�D���Ⱦ�yfOz���d���#�K�5�(����S�B��w[Yh�+���j�X祖���}W�2�U�P��g�
0Vݓ�r�[}C 5�#�I:m�X�h;IL>>F�]	�D��T��Q �B�`��r������Z���L�6��W�m��p<@�:����KWH�3����WҺ�� .3�������sPt�y"
�
%���[RH7�xî�VN��hπY�Z�o:�K�_I.���<f�S�hj��_4G���x,�I�n���;	~���tS��A�~h7�9�@�������44b}�`v��>��au�U�a��c\�g1g�[d�����1�z�[xA���x[�N�ډ���hy;�ɣ������A쉉�,��R�X��2�V���e�CH�=i���AM����PbH�ك��HC�J�q��K���d�>s�	q�El�QlQńѸ�7K�ٖ���:���)�惮ܺ���~yO��b�+
e�)G���x�?�T`y~��xB>o5��×LW1��5�?9�/d<�f�Qc��B�Jj�ǻg��;�
�ۦǸ؁!:#�ظs���fb�zN�_�P�z��,��&p����8۾�˼r���;]��X�,�g��a=�j�N	.��l�K��7S�~F*:���U��
~r_7�ٯ�ST�g�\��Sl�Ӭ��;���[d �o���ŋ���r�)�~(n����?^IY"5��M��9��3?���4�[��i��G۾��W5-("~�[&B�CUA#~dk�����N�P!?��2!y�5 eY�eњ�3h���;�4�� �;*5D�U��4�)t�Jt��դ�O�||�3SQ	^l�͞go|N\&��=]�M&��h8c����P�>i¥�%�o7(�RP��\ح��r�]����0�#�l�k�KY�sN.�3F���YK�&V�:����R����A��S%086�_�.� s�W�]_/B#�ɇ&�ΉB.q�����H�U�F5�6��jՎ�dȪ!ViLܨP
7-���k���v�b��5�`��nx=�K�P=�&j0=�70�',k��� ߳�u�"[��4Ǣ�����\�r2�R+�X�z�p�D�S� (�M q������U>�y^un��L��-M�6���,��:��޳R5|�%%؜�T��-^KpS�J�w�����X��pZ�����#c������SLyӥ�)�6�M|��օ� ����4��!-I�V<@������X|���*f�M+�ss��zG  p׷݅b������A����W�P�[�0��ybL8KddA�kt�l�_/�������V������PW�Ay��la����<�~�x��S*̛p������=A���_��=�W�ҡ[��XKt�q^C>G���a�o�MUIQ����
1��9���IAE
�m������[�n�Z ��^CS1j��Z�`�K�m�]���}6Y���� hE�>ђ�2e�3�G�_��5|�d�ߦOtrwO#*5u���(�Տi&�r�g��4�����X}���^5��q��o���D�\cP%�XrC����\.[wO��Ԥ����-�7���V &i%��= ����"9���{�Ng{靦��b���qZ�B������4������*Sp ��yN��An� V��v2J�,����B���������41Ч}���6�\6^�. ���qH�tWR@|�A7&�/���(4~r`�[�v�,��v'�u�}İ�.��f���4��5�7��;�hf���k^�Q�׿a;��*������b��B�P��O����?db@�.w�c��v�r��'#[e͞�#�\u�Y< ᪤+dh	� h-�c9���$#��%[r���;�e $��	��P,/S��ӔT���;c�R6��m����Q���� v��7�<��!�hAg���J�Uq�1�/��t��+qEsQ[k� �&^�ש>�Q6�+?TG����wQǇ�
����D��������HG@�g��T.P���R�FG��n�^D�N��{dU�A;?;X@]�9��<1�7f��V�B�3�y8�v:S~�̅�Fdi�����h��*��gH���V�`0���~�Oò�sY�-�=T�W�(G8�����'lϛ���q���{��qp���<�w�%���FS]����F���f[�2�@[4ܖ:0?f�ܩIwC֡�)z.�O�a\, �\�Y�Ҧ��&�^��z�Sxb�扑+�#����E(��xY�"n�V�a3.`S$�6�ݧ�[�
�!��AJP�e�Љ�����9
�*(�(���Oh+� hA��(d�u�^OdIjnN:TRR<	�E�Jk��B�}��L�!��B�S�RR����կNPV*P���Q�m��Pj�,8������X�Y���#}����n���27Z4	�Dk˹�͡܆��0%k���E��j[�U%�S�!܍���Y������@+�
w'kV
��%�ާ�`UQ��}`Ҡ:VH����6����F�:�~NBW!`'u#���-�!O���}�a��/QW��fװ3�H¶E��R��| ��N8��P�!�u"�䂴���S�(g�e�+]��!(�i;c�u�^{MqD{���#��n^��4qE�4�%��PyN�[޷V��=��NS}�� '�Rf��(A��P��i��C�����)��|�_�86�-�]��������4.!RƢ[�ܨ=dHM���`�Q�^l2W�q$��BC�����kA�ޕf5##
��_�Z6�4��[��3����K��0#�G�D��#?����q�������U��PI�1`�p�����mn������=�tN^�V�V�K��~�xzn�����W�O(�
�wu�Q�o�S+��4�^G��5S����fAx�*���{�B7U�߾���	}ɂ�$�c��)�Z��Nwe�)�߳�����?��`/H/`�޶MŹ�@�+�:ʀs�����o,�xsl�+��O��߷�F��Jf:R�sF��ĩ��J���J�=�֤�=�x���픚��S���_�����^2�&��*��܌��=��[�mѺdQw0x�^l��\x���Zii��%LY�|�����嚂q�KD�\�`�3QmM�?$n���v�4u�\�U��:=��݊���v	ٮ�v�?e���`f@�99+����(�F������D<q=��Ood��t-��^�.*tʌ:�o�@��γk��4��1K;b+t~J0Ëc]��xo���5������<��-;&���0gXpNhА�:Ι �]��92yR���Wwy��c͍�m�m�2zK3���!fw]2;��K��A�C<���u��2���;��4,p���[8ͪ��/�l ��(T)w�f��i+��"PX�̖X�K6� #R��8:vݯMbV�����tpm!O��pq�Ղ-�#[��b�RM	�s�
l��cⲰ�+7{)�t�,�T}5��./�:c�GĂ�u�%���(�օ#1u�ӽ�L���\¿]`����!���g61�kh[�T�]��3GZ�y�u:�[���,��gs%ۮ7"�{�d�<I|ѓ�|��%#�1�!����;cg����}B<-3cw�B��<�),b����Lņ����~�(1ꊬ�W���7`���gz�����oOb<��*q����D�Lek(�PS�[�=��#��k����tn͎��vcw�:~m.������O�J�'	�����QvOl�;��J��C�H���Fo\a��{�q�o���H�>�W
���@4u��$�}j���d4�ܸ��y�Ų��e�*�ص^�f�J��lc�^y���E�i�W�z�ʬ�v#��y��&*���lV�*`��}���x�Vk��<�06Q b6/Eڍ���&��^��k���ZX�>�r)��F���c��H�D|\L��U,[�qP?���_e��?$��RN �?��*ST����=�K.�6�*4o����Q�-@?z1#��<�k��F��ëGiکR˒@-���^�
�}��̃�NP�ǈ�*�V=-/}�1N�\@�������N!m�xh��^��18��Q�M�ɏ�c�:�}h�u:j�v/q٧�
I
|5��Y��6&R���Q8�p��{�r����i���x +��34Ӟ �1Y���b�4?�<l���z/���-k�Z@�L/j�q���I�_8�ğ���q^!@��[��\�ֽ�M`��7�A�2���z6��E�퐳�ᒞFV���~� i��OR"/iY�����0IW(��{&&�ռ �J�Y!s%�;>.��1�ߥ��O�kΝ+K���k�|{�]s,�T��1�z��"g���~��([�[�)�q#3�(�v��d= ��ô�����(�	�>����T�������Ϳ���$�g�n�H���o��u��;Q^��/��qN�>��e��k^s3o���>�?C]�6�0�=+�ƚe�;�4@�R��42������>�>تl�����óR��?P�b�!��fg/0��`e~�·k��6��xY�ƶ
at�{��%4dc~�e���v�lo����eő)��:��x4�8�[L�&�oH���Ce�F,��V���׹OƋO���b\���/��5��m�h�_桕E�ּ$�L�x9���V����wc۸����ϔ�i�dv��Bv0Q�xͼA�w�A��0�%��O	��OT�[ގ�����g�^�.%��+���z����'ٵ#5�m9X��y��vN�p*[��n��T����F�c�3�9��ſ�1��ر���+5���{p�!NՁ=�é�'�)�h�h���Q݁ͨ^&]��V"�|�xh`��BU� ������� %6���gf������3g����.��,Xg��$&�)ي%q��H���T��� ͪbģ2G�W���������M�P�G�ڎ�K�|үh�����㎋u:zxZ�r�siS4��S^C��y()��73�����-^+��_��Ag��� (U�����w�1+Q:"j��A��W&��� f���n�}kb���%y�Ӎw��f����ս'lݺm���~$�Α׷�C;�4rtj7o�s����}�4�]�(��ϳ[ʺP� *��#�W�^���嫲�A�������5%�~����L��/�tn�̵�i$5Zo�I��!�
k<�%�Y�w G}����e��'����͑Y�Z�?v���+r���pz�7�u�DC�[��0
��3��<���$���xmX��;$���'UțS�6����8�R�6�����`O��*�d	���n�WIJ�9��l�<?�-�_��B1!�̠���-5�޹G���=0tA�ߏ�h'��o�q��<.3bis�(y=���E��H�J�_�,�@���3fU�������ޠ���/��x��4/pt��6�x�\��� P�@��WT��2�MĦ.�ה�E,<mm5���9s�OL�f��R��l�cjK��y�DT���+Vs9��41I����!��#[��X&��V������{{��l
�_o'��Qj%T�����6�bK�6ԁ���Cn�Vf�?pt��m�b�ks��s�0R��~9գr'��m()>��pF	N���!e�D���K���X��%܍/)*�s`k3ㅼ(wڈ}��b��.���KX�3S�?S:�v���]�4�Z̍��m8o�YC^bʨ�\$K��֜j*(�������k��}z�L��=a9f0���˴�5kB2�7���'�dBJ�E��(��Yp����ML�;�kp���$��m��y���<b@f�g]�:����Z3hU�����Wv�D�����4�޺����� �٭k��,լ~���nVm��7(Eӫ�2��P��5�*:[@*?�[�k���9�-��JM4ʿ�\O�+;��==y����n��)�҈�o��35pT�/D�usG����3�������64�/������;�9�j��<�ı�����AK�d`׫l��P����?��c�sJΛ�3�9۞�.o�+U�:�Ρ���_)W�~(�=���q��ݴ9���t^<�JĨή��e.��N�OFr(6���9ڴ���}o1�`�S��u	(zf�4:?�S�{�~&m٘]�u�(�{G�g�����h�,"Gʴ�FR7®�u�"0��[��C���ܛ���!��<�4B8�pS޵I#9E�Cp��a�A�K(�	{[��z����Cg��+�Z����bv��:b���|S�$�h61���r�
��!+��8I)��i&9_\�=*hf��Z)h��-Xԝ��'u%�r%� ��y���.۸6(�"�i`�#&/&)q��1�im���ǎ|ej/	����z�ԏ'�_!�(<$�Q�RSO��0���%8E�ݸ�Z�us��E�~,���؂����T��1��G-� (d򕈩50m��M|�f��&��%Q�<��l�r�Z�p|r�Km�<��'r�T���t?�+�{G!gP<�Q�Y\�_1G��-���堶��"�Uf�Hb}��0C[^n���q�֔>i���l��R(U>{4�!��ۂ�Sd���S[���RrDO����^�j�CT��O�ۡ���i�X�+%��	
?���q2Qh����0�E��*�w��!�@�ay Gfe*��E�@��!b�1�K-�7�11�i�]i�\�(�1����p���t7��1p.a�Z�0��<2Q��g^�����d�#E2Qa�p�F��Z��ci�͍Y���5Ҋأd3Ii��x��&NĲ�5�k�!�}�y����T�?����h<��I�{��_��%R:3�-�$�<y��U˻�W��u8/+���s�^��0/r8��*����@KІ^�<�p�#��� ����bZ�.�@�Y'�V��Y>ꆾ�є5�oU�Cu�ſ��œ<�9:������/�Z����u��X�h������h��x�<JqWV��1Fy�C��T��9�� �ު�+dg~���S����RX&�����SX�\ b����o<���V���A�M��������l4ِ�Ͻ;]�e��Е�#.XZ���t(�fw���h��ؿ��˭�>�i��ʌ9��c�Ֆ�,��e�<<&{踆IZHO	��z�@7��}/�6��ß�Z&�o�I�Li0�ڌn^Tg'D�(kC�_�OVS%*�WXW-i�w���ݐ�Qs~�_Z'�`��Ykǔ-��ߤ�Jιc~�♁;��R��&�hI��He����[��k�7��U$�"�<7�8�L�N�lW�r�ܦ�j�EM�A��<����?��k\�����y]��
�f�?rh �G�o�Zh��0��)�l8k7d��So���{J�Q�Qa����Y�㍷����v�u�bD�<����j�X9tui�Ek���R>�8�1#cV�q�qb#�=�ӂ�P	�L�s���ؗΘ.��� �څ�j�+�K��]�'���DoV�3N".b�IO����z·ϊ�VW�9�BH}­�)�����Æ�6�$D◀.�n$$_��"�eQߛu
lB�Y�x�G-���b���y�lo�gDy���bOiB���J�(e�s{�^�0!+�^K�F��r�ѓ��T7�bͬpP̄Ҫ�]��s�
��+��DSk�թ7o�������5�՘�!���8u��뗂�5-.�ı%}v8��S�m��
����3Ɠ���m&�hj6*ױ�E��}bt%�<�xV~�R[~��������m�T��]����Z1]�S�����쑱��n^sC�����(�W ^�J��k��~�W��%�ĖO��ށ����4I��ٲ�ܕ�<�atjc]Y.P�MD*)��G-�n<��{|F�&��Zgo��ZI3abP���L]a)@��ù�i�������T�]�q �f��M��^��j���%�DG~������<�*f�O�v �.�ꌋ�\
�� �}�� �0�[���3dp�V5*��lM��$�h@���g�n��h
'��{�U:G�'�EdU������S�	w�l�j]�ղ�x(��kԈ��X7[���	�0}r�uA�ź)h~D8Q������n���l ��oY3�[����7�*�7#֍��yp?��b��2é�9���֏eъy"C�*�[
^��+�U��Sġ%x�Uah���KM9��I�ޢ-��G��1��P,�SX�e[�s�a��J��;	��1�o�y���		���}�3��F|�,fN`�
��fٝ�B'��63�����0�dj2_y����g
N��:�0���.A�aG�qn��\Oؖ�+0ы�]�ZJ�!Zf��׿Vv�Q��〕�Rτw�7�_�����ΖU�ܪ��(H��2Q�(� ��X����N%^*���`�Vrā�y�FL5L�RtNA|��4�\Z�8��g�
w�?�s��	Yū{hRBĺ�q/��]ӛ֐���^����Od�p�S_?�c�`��#W��9�B�/[��m��)�ri��rF�2�Қ�@�oa�dg�[.�;�����Dj/�t�_W_.C����T,��2VJ�ssA�!�Z�uPd҆E��%�6�͛�sĐ���\O�7}�M$�9?|4��E%��^[+W�_�?rM�5
�CV�9�m���ؖ��8`��~�����e��VՉHT���uE����s_XutX$|�T֣��.�ι�T�(K�C	��J��X��/�F�#2;h����ׇh�!8m�a�oSC�Z����$��phYf�{�@t�`�����6zl+�_7���D��P�g����W,,CԞ���*��_�$��w�e�gpѐ���u��n.D�_"���H����B�{N��Rg]"S�f��3&j��_�b�_=��[����c�`�Wc��(Ydӓ��<QTY<�K8:W���͹�|�1y���u�e���mgp��f�5QS�?���~w���h}��(��!�.��$W�Q���18wH=6a�`����S��{%����p�
�JR6��-�/��e��n'fu���/���	�-�i�w*`Ym�}��-�({x�O���4L���ux5$q? ��/���:-ө��m�eJw�]�@�n��͒�K~I5��>	����7C>�Af��FR����s/�^�h�w?�2x����؏=,�<�����N����< A�L�Y�Y<a!a�h�k,��kQ����O��;}b�\Ɗ���q	�;��,q� 8]���Y]C_�,��g��dlq�e��b��%�uڝwzOn�"t��)*�F���MV�/��}\����~�ed^Y�m-!t��7&~�W摡sm�*���?�ނ�bl�7{�����~�` $�Ë�,�Xؑ� |asP��E�=��5��ғS,W0LEܩ]%X�rW*���ɉw���T�<�A!�"^�=YB6�>u�.Z�{�N�$V��Q �%�TO�^{�N����U��rS��۠v�2D��p�"���"��hQ�x�{O/���ǥ�ݻ�����	|�|�_:���|�
��5�����e�nd8so�E)��
�
�����6�[ʟ'w��~���F@�X�N���/���2uW������dm�WW��fH�l�c\5�C�"E��qs�B����o��+bZ٪���j�����(z���C�fn܌\�n��
��Ni�`�ϓ��L9�FA;i��?�����)��t�͋�d��f����o�xd��E6E���F��H�D6�;K��y�t�߸��9�\����R�h6e���${E��0���F+H�ٵ��?O�+yψ5rџSS���;�G�f�����J��g�
��J����Tⵍ���yp���6aǆ���r/٣�}�
R]�o��=B��h���A9>`�8A(ި&�At�����t�l�T�BMGB2�&I���#-�x�ŭ������^>�����!���"�)��Q_MKv,��Ъ����4�ʧJ�����d�J�&n��o2M�/&�K%�` ���G��� �W=���Rǂ�"�
����6)�I�����yX@#��H�t�2{"K�ͬ��ky��Z�w9�2h����zgb�0>�i���s�z�6=oR��|lA�V\:����;�1�|�o#�XG�*��If��Z@��J��C�����
����\�[��~��]*�u)rR����U��-�AQ;[gN��8���$�\VuD�4OsJAB�Ёm��g|9�N�0�["g*����;��?��)�F'IC03uL��4����RH���B�x#�?��IǮ�;�L,�eWT_�ԏ��F��D{,��x��]gOp�*�L�i�x��m�,>�|%g�3�w3���@;-7����[�;/8�j��23?X�މ�����L%ݖ.�]����4��1>���E�:�4��p]I�1���� x;���z �e$�����fOmIn�>��vt�� �Jg	��6�A�����z{�OɏáZ�I+�s�ζ��e.F��(�S8Lʾ!-�O�2��,�Nѧ�%�:�6��/�����	!gQ����������)�����پKа��*W{��g���ʨR�f���t }�@a�q�B�eHiD���i�ojG�m���Љ�W��7~˺�t��ʚ@)-�I��q����0��w����k��^F���������ږҩ�=�!�6�t��hGZ�rj ��9Z���M}��7�p��ba�Q�A�����k[��}|]��жˮ��B�1�x���A���B���Q��6�H��W������$����x�q�6����fň�,m7٢�3�Ӣ�lj����
�)f#�P6n��j{P���M�A���*��S(߁T��M(�頭^SOd�	 �P���]��ށ���ĵ��L��3��8�&�k�U=C�x�=n����ny����kqI$�kѲ��rf�A�I�u3�֔�Q
��.dse�7��,�/2ʘ*ŀl�:�\6��^��GѫyVj��u�	�At����og�0�0[�q��	6��K���[�l[9L�e/�����sH��g5�Lw��4%L�;b�x]De���^�1簭"٪5����+�4n~�4�<>	zK�*����nB��H�9q�J#���"���KK����Ts�y78@��}���i�*� �7n\��_ ���u1Qdi=�%���f*:/|���.��f:�%x,偻���AM�/�d��iSR�� %1�֚��"z���͈űF��o�A$��@�F,����k����)4:��|����3c���?�vґҼƨ��K	rM�Nu�P�Y}���@�SI����@Q�eݬDu������%pLP˰��	E�n�'�@q���r��� ��!�t��+��QY��"�&prL~�):wd��c�m�_��J�%%1ǱM6f��Ԅ����W��k��t��YK,녬H�^�W�����C4T(�u��]��8�#�>N!����3Fc�<���i���TJ��~���r���K�0��w�%����]W��������8�"r�+}g�\����UGB	�xj=U��͂��R�f3����@�\PH�$En&�����^Q(&�c�X����R�w�8�_�[#�Tu��Zۊ���0D-iF,[����`��]D��=_=v���?'Ae��b���CU2��x
M.� �&'�8vy8�n��Jh)�YvC3G�����&3>����,�Fnt^`5C�Z�8şR8d���b��ئ��h���6�>�mV�+(�Ǿ�bM֏%r�'�T���cX@�/���֭hS�@!�Z���t��W���Ln��t6��W��+��蓎b=Jٲ,��t�I] H��y0�d�O�!A��4�65z��c��	v����̟M����g�Ǭ�ٍ>�7"z'&y0��Zdd�����l�`���[��lc�kz��ﶣmUd�$N9+�D[*�~�Yt�<�BB$�#ǝqe���ȐWi>xKмe�pz��Ǳ�b K�0��jJ��l�S� ����YM�	Z��=��E�a�x�;m�+h?!�=��BL����c�C1�T:;��j�]�=a8?��yUQ�7�/�%�ۍD��Y�wp©B2EH��F;��Xh\R��:�2.�1.�:���0�(������`�M��o�F6�î�a|�Yk1P�A��;֟�+��)]@{N�o:������:�Q~ܺ�QE����;�����w2�?����U>�zw�"U�	�N[�h�>�A��ӿiI鼗��2M���.ė�Z��bI2�����9�}��ŕ|/$��s��f��`�/-�?T4Or35C�aR��U����9���Ȫ�F�=Ey�K�g`j͐*��_37``�*��ݚk\�:4��I_�5��=�3�Z�o�)��u�C���m���FCW���@���ᅊØ=�$E�d�bq����aB��~�`���!"��5�t{{�0�k5a��U|Vr���%h%�?ۣy"T�p��5���k|�;���N���btYy"Y�O����:;/:�=��gX��W3kg�����}��̇j�
D��(&�j�#p����).��|^��m�NB7 �7�c*b�̄)�A��~h���lgv��������~�f�Vchq­u,wȉ8�1+�ž�ET1�Y�u8oQtEz�_�i�n�fM����Y�i�9B�[���zPҘ9�Q�Z8jegoTC�� ����`e�22:ofS3�7zRC�s�]�����/Os7�YTed���Mb˭M��qW�憩ۅ�t�R�Y��$�p����e��WEQ �ܤ����]?�E�2�G��jd���镔ö�px�i��^)�=J��B�m��2}�p!�� ���P���{纄���f����X]�˴M� ��}GڻI���;ۉ�JjtӉN�a��v;��qQ�Z*l�'�>���i4��d'6�>U���ڨ\Qre� ����Cl�2�I�'	��.�ώN�j9k�E��$А&�q�z�C��9��&�źc���a��y���]uo�ei|D�d���f䭘I"� =�}vӲDт�X��x׻���$ޭ��g
�Ĺ��
�0��.임9q�d�t-�6-Fr�>���[�% ���[Y��%D��H"�1��h^!@�x�F��5j�S��O�dRz����#���
��z���(�ݳ�����x�����'��|+.x#�lZ��nu��7L�Έ��_x����<S�v*~ ��pV��r���2�O)��r����r8k��,�?���
���`%��|8E��'�FmNI�j�]�b޶�|�ĀOʬ?�*-fZ��n���&��V���e�j��XJ��L(����- ��*e��Y�����u){��d�a�R��	��%�xMl�r���������FӑA�P%~3�(Ï�˙쇩U%�n����w�UWl��Gp�Q������7޿|�[/�A��&/ͯs�Y�M�H����hA��$���U�2�w������1�r�GU�
��mu��ےC� T��8���^O����l��y3!}���Y�ɓ�����D	z9�����_x*�u����C8O[0q$I��f�Ϥ<i ����{�4J�N��ns��Z?�`��Kh-	���6��N��ߖPB@
J�wX����	"ʿ��rz�Z�<��73Dr��SxY/�����E ����
��5_�95�
_/0��/��7$��-ɂ�JP~~~�'��^Hv�d�e��gf^i�׺[d� �
�Ŷ�Կ;�>�(�9�q���/���?B_��9�s��K�;)$f�[�ЁO�kU�xK �~9��`�1�%,�Qf��BPFD�\`;�H��G�
�1x�Z�
���kr��1'�HKC���5#��0���/pdJR��Ps�'E)�r��9s�\�`���y��V�$���#Q@T԰�R�ϧZ)�{�q7�׭�l�tٻ�R��T�����ҊV�UK�AɗE�DQ�)O%��5�U��tن��`,��aV��vJ�/�.�ϗ���4��d)�'�רO��o�6��8�����f��3��3~_��Z�r|c�9�Uх<��[�e��k��bo���P�Wg��z����l��f{C�����!�_�2L/˺uˠ)�`"ق&]�1��c�Ex���.H.x3���&7c��R!��6>��q'�p4i]�*��a�a�[��]��'
S�h!�A�~�L񢻵'|8��Bi4M)_��ɯ���Գږ�z�,I_k4�-����~�S�8Z���='�-�s��Ώb#��	jDD�����'Q���H�e(Qa�H���|j��xC�w�P^t1"���,6(�sU��@!����o9WN�Bѯ?��3DRض��RSnWG��#��G��$Z�Jƶ�,�ϗ�2nob9�W'����Ƕ4���~�/���?��N���g���,z;c���^?�g�%���[��3��H���,1Ս���ыiy,��Fjt����W�	�i�H���@���aB�����s�U��7	a�/C����1?e���CW����>�1�\��ZZ�u��p&K(I���%S����\�̙�^WV�4|��#˨�wв+��W�'8	PG�i��I �OE��	<�����f�k�C����k����^�Ⱥ�6�K��R����y�c�ٹО�~C��O ��@	�Q�'���e�*�a���.�~��&��1q.�_͡N�e�������V������lҥ8ٌ�XSv���dr�iZń�=�M�)o3ֿ����if�+^^��H��>�A��\�3�u�J]�%� �`0E}X��>*|Em�w�	2S~��t�(�g�fn��*Γ��vu�TD�,;U�6�hS���%^x�`�(!S�4�C�
V��+�\�?�w�{����N�����&�"cMi|u�SLm���v͐c$�U��٣���W���2�U�9S�&��I�e����^�0�i&���K6YuJ����䯳�:��+��p���|���Y�;��p$�&�P�Ą���P//���wNW�l"�����zØ�=K/x�d��Җ�����6�H���������VtZ��/�2�{h�<T�C�!��Ux̦iO�7�PYzXg�F�\�V���\h�֭O]����c���}q�����a|�[¢���h���7�%��w�[TiFD�4�H���p�u��y�CC����4V���{ŧ*!𮖣�/���^���!J�"�cj&�U����ޙ�-�1i���5�73qȵ���A]+U�(����e ��WV=ǛToL��L����?YS�6mt1�n��R�H����@�LI���C���Qw�s\ZnYh�b�Y�h���n�:�7&�r�gH�s��#\����Q���ʬ�ah�9�(C(�%���z7ȜĈ��?h�W�>jY���d�9��oZ�K8��Wp֭;Kփ&�}l�g�cX��o�m���J����;Z��Y)�uA�1�l��8�AI]Q��@���Ԭ�J��Жs�]ϝ�pyD3��_���Ԃ+'� �Ê*k�K܊���Z������� �v�	T�FrM�{����Q8��ߘ��K�[��L��COٵ�'m�*�c��|h�ܷ������jȂ����l�ț�Do=�S�u�����	��u�?����5s�Fŏ�LrP�\�ƏٹƚW��m���[�BA\�u����_�m��y�:^�SI���m�M#�.��ڍ�2^xzmF��B�G��m)�=�w�����qǋ�*�^"٘��v�-�U�)k�#Uw��q�@Ʊ��
�pQ��tz�}�]��й�2=D�<nC��k;L�=^���Q�h��r��R۶GXb�<��֙��Ys���K�ߖ�Mad�r�W��F�[��W`|�:�V�)~;�K�*-�#p�7�a�����O?+?��j&��'?�8)DR�� �]ۄjy�������j�a"��U��Q�����zv��QNu���q��aǇ�8����~����?�#���.ۓz,4��.z��b�K���JDVi~�F�:�]D�U[��RM5�(���(�;6j��+�H<����~|�l�8О(QZ�9��7�&T��-�oC�	q2�]�F��J�N+�=0��1u��W	/����h������iW!|cעy�
^4�Nc(�B�g�2���`~��C!�`�4/ � �Q�Ѵ+*���E��᫐�G]������QV'l�.$�K<A7�����ԏ�����D���=�L0��^7����Z5�� �Yf����R5o��Z��'��&������49���_:�QԢ��pͩ�w;�g!2�ά���:~�q�o��@�[i]co���Ã�e,����%3�s�Ϸ�̎�0Җ�ք)�n�.R�^�:<��
y�@9x�!ä&��&.S�C@�o�w�F�C5(�қ�C�@we�X�Nk�1G�d�r<�9�fM�-��Q���<ަn�š��K$�޶�A�XE���2�t$��B��P�@����
���Fs�׍u�P�@U�u8)�ː���M�VE+nGѵp�gnW����«9�	2�彊V�~�� &�)�C�lT��&mW�+��1�2^%?O�$n=KPD�ۮ����������;$ �W�a��Z���TSr:�'�S���s�	�K3By�9'����<������w��:g��<�//�o������*�VB��pt#�o�)6��
B�;D�T�!�!<ބ��e.͚��x�����������9պ&ռ�;r+�)��la&mׄ-[��L�i��q�����x�t�q�Vbq�J�8
�v������`�Bɍ#H�� F~��!j�h�@���H�D�P,�E��y"�K%P���j��j�f(/�d�B�C��Fo���*�?3u����Ιm!pf�yk�Ԟ�[�p�j@T���ҩjO��}����4���%9���!��}��`/hڤjdy�1v�DuJ'n�
��ǥ�W�cͽG"[����1�؊I�kS��n�:1o!��wo���Ў혿��*C���/lu&P�;XL��)HC����C6���� 	3���L����i.t��J��c
��&��	�J�%�W�����dK`J�m��98<������i6��0����&)Y�kZS�s�#ۛ��L�J�	��jK�fL�mQ��&+1��vu���C���O1G6�-rV�$�d���D(١��~�W����B?����}R�1~,&N��Ӄ� Hx�	����	ް��i���E�\E�����.�����a��(���R
G)�^����H�C�uv��&�Ñgsuo�2%������+Z��Q�2Я(��2
ŝ�0`�����{��X)����I��Iю����\ g�9'����:~���ϵ�#�q[����6�?9�E?D�Hr�>�Lt��@���'H~U;e����S���<5���s���}DW��ᣛ}J����*�L�(c �e����]i���C��y�\����d��TK|�U��·��Q�
bh$������=6�$WR"�ВP���"�s�מ���C-�/�ҽż?|�lp,*T+�}\��B['}��sЧ�Fu���e��(8sVt����E�*��b�����2�s�D�a`�[��uw���2.���!�Ȏ�#~�wG�ir�f��0�����Y�5��Bb!\�/\�8+D�x2�V�MC�n�$�\g���fwC��:e�~ywӰ��4Z�)�խ �'1�T'����
�D5��4=�X�Ƚ�'F��O���5}l�i��Ş�(ʰ��L�ts�סFU�e�{(s>\�!���oG����9���	��6�aIߗ+��,��8��Ʀ:$��A��C#�C��)~W��}y}	fHr�L4̈́_�`��k�Uicy�N�g�;Dӑ��i��/�@� DGMQ�R*�.�cS��Pu.W@Vh�7��22!̀��	O��P[��D|Q�U�&��*�:=ē�lx�%�+3��&Z�'�MvFہ��1�[V�cݺ���W�P>�+f~}�T I�l�ԗ�P� �P����5c�<�ʪ:vC��f�+�Lz��y؍/5��Bzd�8�����g{P7gb?7�@Ɂ�Nb�DB�]N��^�C�� / RT��G�����
�i�K5%�����=��(c}\�����1�o` ���L\D$`�C�p�d��%|(\�r��K�qi�H�I���<����'��:t����Aq�"bY%e���$���8���f6Zxsx>��OY����aAR�O�3j���������K�A�m���ǃ�YN��tnn�����=X��b*�&B���-�/s��|��7��<o��/,� ��T�?y>�N��Э�^3��m���n>���7:�Eh��uO�ʪ��d���W2��ܗµ%������~5����|۷a0a��IN��-���=�M �V���,hhG�t�]��*���Ŀ�[/�ޑM��>7��������P�����"�n�����%�*�3i��}�"s��<�w���w��C"��
c4����)�W�"L��h���9= 2��Jx����c�R�Dk@���.�]rI�c���!	-{?�WС�M���? }e ��;x�����<�mF�AM�=`�,�|T�� �ħ��z���.3{\C��.K?6H��]	��.I�-���N� }�h���c�uK%z��Z�mJ��QM�
30��8|*;��|"���~��,�wo�m��L�9��b֞��<�V��m˒��% ��օ.PLYA[��j(~yN�@IA�F��O ������ƿ-l%lgc�ͤ�����֠����&W�yy*�;�_����Q��ՌP�l��׎-J;-|ͧ@_�3g{���᳦��'�`o�Mmhĸ���1}b�X�/ʻ��ػ��Y/Qd�������k�}�¤��=�d����B��}�f_��sޥ��Q�=Ս	@�W�3�s�1n^����C#�X�T0�����#N��稶�}��X%׼��l�lW��S��E*S-|��Q�J\�r��u7��� Ċ�&����EN�Z��Kj�V'���[��C�aȴ��_�m���C�Nܱ��?K�[j"�[�wLy�$�Y���1m��}0{Us�<����Q=z;�J��PUсy�<ϒOl��.!�#�D�~4���b�pIe���d��n`�:n��L�7��I����9�פ'�]�����v�W�$��j����K	.���G*0O	����b�`#箉�XC�X&Wo`t^ۨJ��Bj\����0)<p�o�{����Z��Rݞ� �\��T����/шI�#�άxY��z�Nm��~�?��L ƴ튫{V͊�ֆb�R�GHb��١�f�U}��
1�����u����4��9N���w���/����,1O����ә,7�I6m��v��,k3���*Sn��Wx���"n8ϼ���]*��"�����E�DS/�'-�?�F6�Mdvؑ��r7�-A�'�6���9d&�5/~X��k�ȍr.i��L�s��JY�b�
7�g׏�h�Fdw�m�he�U�x�,&�\#�dē��bFBp7�_��a�Iw�/��JN�M�^�QN�`��XP��qN�l	������I!&�j��m�.l|�,�lT�/�l��b-����NÈ��Q�P�߉�Du:Û�Px䉐�(m${YB�k��t�E��v&��m���ɟ����)�BG}{}��:�>P�*�El��S��V	��@�	�G��7̑̼�?�"!�-��B4U\,�������(���Ȅ2s�<�\�iqO����s�O9&��}��{��|N�u'�W~Ձ���q="K ։ߙ��.�B��f�hA�q��.\F(0�1����!&�-�r�/���s��&�9�U��?���J睴
!��K�' ��a���%�^$��$&C�7��eC�S��X�J������ܲP�I���1+I}DWZޚ.�жQ�Q��0|�$�^Q��o�H/�'"ec7j�o�\I�ʯr�h��t�ޓ�~��(<&�7IJ�Sxb�WH��m@�+�êB��b���߇葽Z�Ad�I���s$B��k/�������lN���AdK���1�3!��4^��7<���8����h��?kv�y6R��S��z)t����1���<�$z��ƴ-�s/Gj+uT����[K~7����Փ;�)k��Q ���>M��,^��+1����ĸg�U�Ǻ�����gNr dv)�=�}�wH1�����n�ퟙ�	k�G��ܖ���D+m�>���"�߬��������]�\6�X��6�Y�x��I"����&H��IUt~�]�I�aT�o�
iB�������\#ϳtC�J�(�r@��T�̾j~L#-#�DHX�0K�*W��y|�&z
�7��\�A�CU�*���СŖڽϘ9�Gf<�m�	.��S��yUAx�S����R���Ӣ=�-�)�6{�����|WDA����(���ܤF��R�Qs����G	w��ѣƳ��G+��|�r�(F#W�z��A��A+4��㵬X?���y�E+�L���dɍՀI^�O£�o>ߦ�� �wo�ɮ��^pz�?�72<*���~�^� xF����`��W��,�Nc����a���3I�����r<t�9��}Άf�����v[|�|w=z�!l��BI���NL��B�6>��U�<����I�T����/;x��{Jy:��԰i�����a�aɍ��zk��VZ��+&� �L�~�T#:ݻk�C���i5ێM���?H�J��'@�:�xt;�Ud��[+w|sU�P���Q᎔�[��ʎLF����~b�Ƅ�*>��[n��Y���1�/�&p{&�O��6:q+��P��܋׻�!A�o�j��7���='·0]Ǩ[v��-�[���|��i,�ñ����PW�`ܢH��+�Y�?�����t�hD�0T�