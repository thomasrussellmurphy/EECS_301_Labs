��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_����m�e"kxu�Uٲ"#oB2�-g�j��h�p� M T�(�P�+M��&�[���+"�:%V_��	�Ξ�܉�����_̯��֛%�����A�Y��Y]b������ju��e�c"VoH��7��ۆ9O�5�ҋهO;�������w}7:��yFP~�%ti�_����q`�$H�,,��Y���^!ط�R�[��ʆ��K��oAH(��m�Z��Z$7���+\n����hSS�*B:a�(�u|��<e)���qL4X]V6�2\�= Ҹk��Wg0��l��u�O��=>�j�	����!0_�:?��j���q[`It����ծ��cM+E���P�xܲ�}U=5��3t��n'�Ќ҅�
�X�q�F}��`���+_�f�|*��[��ͫ�Q ����9�e�$TS�]g��6�u4�^�T��Յ��@��c�/�i-`� >$�J�	=�l3f كf�]n�N;��lJ�j�%���|!�h�~�{�i3<��tk��{�'te���T�b�Ы��&��D��H[Ū��c0GRT���(��1�f��PN@z�����2��>lْZ��m��%��o�� :�۷t��g�������*�Sw$�����uǃ?{0�s֟���51��f�hZD�>]��/��|��9M���(� ̑������P���O�T :v����c�N71
ӌ�Hл��7�$�n����3+X�ǈ7ծ{�L�Q&VD�@����^:���c�l��))��=(��T%k�Q��!rz�[��&�k���&\� ��7�����\@����ZN1(ˠet4F������HD�v�����۔?	1�O��W���r�M�s'D��G&���roCZ0�Q��aR�E˙ь	kA��6�ע�'�U����f��䅛�x�;�qbA��Q_6���b�/��q="{B���R�N����1�:���� ��y� �-�����q��6.��Y�Pg���D��F) �?>>��"��2����{ώf�ţ_�tH�+��w!T;&ia��>��2o-�P6�%i`�2����.��Ϝ����t�r�4OOF<Ӊ�vj���R���L����<'�a��Е�DV�Q�`� =5���ew�V���MG4ʉ*ur5��t�/�)!U&s���$�9�r���#�?�Q���;0�| �-'�BO��ϝ����6�)��9����p��ܕ����Ї�3]�u��':T��"* j��˫�1Rώ���PV	!��h���$3h��l��*&�_]�>Q� �Ӫ�h�vw$���?�uU�i�����r���`���G���ݦ�"̦��i#�jJ�̽��^�yh���\�0�=�1:�ؔgL֩ߘ�����N{'���eu�&���LT��\�0}��C7_[��77�-���9�ˇ�'[�8�Uۊ�eB�Dy���! �H��Ǽo�:R
��d��=�U�ߵ��D}?w}BDj��TBa���V���o�:���+Hi�7����]WlK=;���p85���όH&���rR��y��N	���0����9�P��هU�8�_*��:p e���[y��OE�׮�����]�k�G?,��/6�ƺ$f���Z�cJ���I(ڱ:�Y���=���iN^m��[��h,V���?S���$�^�R��C|�h��4��NN2ȧ*!�y���y�)��DT��߽`?�ۙx�ag������~l!�;�u�of��͂��J�ϐ	�*e5Q�Y���Fk��Z�� 33��9�l���	2:�A�|���}�����w��}1e#'*nm�DN߶��a}�(��p�T��eN��X@TtʓNS�_i�&>v��t���[����=e޸�u�/OZ�L�pUj�2�����g��gg�rv�PrK�ObT)�t���Xٸ_����� �o���.|�އ�/ƙ��QC/���!ZÉ.�'/-K�d'�B�817�����w4/H��1�BF��2E��۟�zae�?�cE�	;�I��j�����a�)�UEY9�J*U9o�3��{%�elP('g�z\F�#���O��H��)��������X���{e����]44u���i�G��2|����*�D�N3���i���6ԝXh��
o���&��XL��#��5h�f�v=���4�f����t7(���!�T[�)�\N9]{����UӦ%����=�$