��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|/K�^!�� �Ϊ�I.F3�h�]D���� �1x�ϓ�k�K]b�ec���9�̑�2�۰�}EW��E�aǧ�b��S��+�/Aė �d��׫�~^^��y�4�4pjTK��~<OS[�EI|�ݾ�wi���tW3|��.�O�#!��{(�N[V��/2:DY��6���T�'��:;�5(8���$��Eʀ%���4e�p�;��a����^JN��Z0����> ����Z�� ���1���C���Ղ���Z⥃^��մ��%���ݎ���
E~�(6���B���$�i�D��%����?f�G���Cy�����J���ǩ��5���z��d�޹��L�t���M���TD��Z��oW�����l�$�+{J�M〮�
�qH�37�t��KN�s�$D�^��E�޵�Bl |$�[�Hʽ�y^I'V7Qt'��ѣ|DA���Im9�-���Ww�qG��>�soҐ*��^h����[��<�Npz�沙�����@�-���\(�fR�i��rDz)�J�}���Tw�ǳ�u��%��	�w(�U\���Z����u���%���9&�c��h��h em��N�(� |���i�L��t�4��b_���A��7�VR��Vr��R=�f��8�%=� ���)6Gu@[��i��U#�ޔ�-OS��Ӊ�v8�'�w�l.7�ʋP<�k�<"W���	2��X˵��
2��0¨��q��	Ы{�P��m�	���%��K�O����[3�;c��D�Q�I�PQ5��,��ձ�{Pb�#����3���51�Պ��EAyl�������xZ��⑞־.x0����[�g�٨=b|���j�|O�<�]��tԠ%��h�����>l$�'RG�a'g�ա�����������N�T�s����a�
�Ȱ�e��Ӳ�����D�9Խ]��}��~�5�p� �U�s/�i�$AW@-5nMĨ�U�P|���Rs�
��k�`%�"o�(�汢�ߎ?ի���tDg�*��3�f��h<9 �,���d�v�0I�KWI���B�(W���[jC�^��b8V;�ů\fAG*���{���fu�Y�$�s�z����$�i\���@�C0��z�@b�	�`�4a��c���%I��a�r�_�v��?���S�H@P�H��ݕ	�y�8�]�O�T*x�x��u�hq�D�l�X���g. �f��!�#��2�V�W���b�L�>��A�V2d�OI�U|��=�$��Mx�/ӳ�^����S�ꘆl@&<�lBv�9���F��K?ǙW��U�y�������/���Zc��g8�W�INe=��~����۱��ZP���l$S�|t>re�1�#w $�y����Y/?�$��o?4��q�9�����j����q���[<yG֧ Zl��gR%S�T�	��1d[9��F�Ni�6���'=�G�ڂZ�H�\r�&>�,�!��o9~a;���
vQ�`�ȝ�����&��������I�RV���S�+d�DRY������-�� �=���=��>��*P�m�q�CUpá�K6�s���
1(ǯ�te%�^�e�;qŕ{�����F�Eݭ9��s�\F�j��ܵe��;�_�[v�2ʅs�rr@�*�8uy�x���h5��
�tE�jħ����0^�����=�f8���'���)�ն���Ϡ�F�0�k���M�B��X��
ŐD�}䠎�F&(�k���&;U-�k �@n�sX� q�*I�G}�ՂF��m�a�����|���$PZ�K0`)ʬ}��
�y�C��cxE�{/)G���'ؒ��]�z������B�QUA��6��ñW���AG8gX� i3�D�Y]TO7�'n)�Q;8$a"�����6I���j���9��INfjy��k���&y�~x=��������[��H\H��s�w���5���Uc3��ƴC��!��+� /M��g�$?6�
_(- 8�(��Mʐ<�c=���~>�����v8�3ō�c�����=_���JX�U8��ؐ�Z��Pmwp��͏�g6}�p��M��w3Tg��Rq�+�i~?7gZJ�t�"�	��'-�i^lϰPe~Fn��M$ڙ~n������o�-��v�:�	T�)۳����ؘ����3a�.��,��k�LfJ���I(��7�����ˏ�v͓�_<���&�J���$G�ee�r ��`�v����u�]fU<�?j���G�QH�Ƭ%XX	g���n�(����ۛ��w�_�zJgZ��.�-����o�NN���'�͞���S?z Λ��a�R9"��]��<?v�)]I�L�&�'�;�t�Ч�|�ߛR�ޤ���|�~"�
��k��0�Ҫ��j��If_�|\��f�{F ��4G�>�2X�I����&��nss�갶f����u<9��粚��]�.�W"-*��+H�|/`\%e���Y�(z�:�ru�ꅚ�GN)G�P��%��0�ةҗu��!�������^yS�V�'��d��������1>M��,T���qme���{Lwe���ĕa�%\���E�]a!X&�{{����rW���
VC[V����k�Q�����V}�l�3��1'��E������4�2�>:�t'������{];�,Xz���w@�~"��P�*���t���G��΢/��e�#c�6u����\�(`��iL[�*�o	.�u}��$�H���-��N4�l��"�Dî�y��V��0�x�R�i��Zr�� ��v�s�(���̾��#)��ِOz���l M��3CD��1�7]0c(@� ��T�Z�ƣ�	�P�0_0!9�@���,���+�@||�,J@Y�O	T,8��p��C�2�q�f(��2ǿ��/(��'VyAG� )bs}`��1 M�/��;�Z Ȍ��l?j��	�3�i0c)S��օ�O�i㺻���.��yS���+�z��D����Z�n4ï����t2�o��>;��i�.��)���b�_�(;��7��&X�4�%�v�)B��C�92G��,���շ�w���G� �i!%�X���;� 
�2XC�~"���#>���g����� �Q����6:�.��x��(��õ�R��eˮفq�n�� �C})�r���x�Dx(�K���y�� vBF�%[x�휦���&�k^���%��6�kˍ��Ķ�H���0��O�
���ٝ?�� ZL=�>��}����/r�.��xA �ѻ�pd)M��v���:k�ΜmX9�М�#=�6�<dR�"e����9S4Q�l�!S�{]����3��g���u���S��P<z��\ш�h%��Q�x��+5�i�{]B@8��ds�8�wFe��	�_��D7�(4�\��]
E$�&���/Y4��ZO��vZ�V�)|ذrϮ����ٲ���$\�<cwW�*�$18p?)�ἦ�҃�*�C�-A�{��'�~kat��ٿ�fX#V�9���m�  �<P�ҝW�b�
���06�3O���@F�C�֠��yg�G�����l�4�r��h�
��q��`�y�ԡ���
�S��n9p�n��N��Ea￿�;��"ͬ�l�������V 4?|]�6+�q��#����щXw>� ��jZ�����^��c���L�Zw{��Zk�aL����x�Y�:�S~Kk�,��GQ@�L�UCσ��t��o\#c�þ�! b�	��2�"СU�8��%�q��X�I8�L]�DE��;s�"����l��pΠh�����b�鄥`6�ҋ���6�������x�`^ ��~��7���3��1v�a�{���US�|�[�B*�s�ݔ�D�Ԣس��%���Z�):]h�
7�T���H��~ê�h>�W�1�c��V��S��\|��<���l� %L��J��l-�!���\l):*1�I�O�u��Bi*�00;�7��h��A�S��Zg��\�a��ø��^�]`'��"�M�X����Eq	\�-��t�����lⶌJi��W��S�a�Ԕ|���p��H�-قy��L��iY�ռ��.ʳ����"~tT�>p�%�
�=Ϣ)�r��vE���w�е'��/�A�N�d�҅}jͨ��Ңn��Êұl�Oo��i�đ��5�8�$
˦�%�Ԡ~<TB\xv��d�LD��F/E`�X�jj�}�å">B��I�,�ڤs-��q�o�;���*�~"ej�S�XE
#;�l�k���+�w}�i>!n�@9V鳌�"Wc$Vnt�S&<��\z��,Ȓ�m�܋d񖘑��CY���5�r|5aA2�D���,�#��Ua���yc����m�T���{;�E��	��?�c��gi-	Z�j������>fl�:���U�����1�'Zٵ���6�qL����f:ٲSԨj]�� a�!��Ё, �PU[j������^�2���w^xrg�ѽZ��G�IP+Qv����7�3f��1�_�[�4oW���ݔ������#�A������;e	{�}UAg�ؠ]��IEʝA���;הR���מB�W<���k\���底,g~b=�̘�k<����b����M��o�){���|�\�qEzU��dW��)__�u�6�M�BY-�U�������iN�C�_W ;0j�wk!NO�Hͅr�_���i^�f�� �V��P�#E��rr�n�e�U������v0N`=��X=�R$��#�����3(��.��m̓<��ᓲ�O��0@N��u�0�O�Y[�d�����7]�i9�#�|���+���mW�#���`H�/u�x��W
��df�f��Ĳz��à��J<�Db�CP4<�2Һ;�6^xJ^w.9���v|I�V[�c%�QBg�)	f��>��cnD��FM����O��YaYe�z�=XBTm	�j�|����ҍ�=���g*@���Q1Հ���H��4/�3 G �=`V�-�vG���{�&&�� CR�3�s�b��T/�w��C�#d�>�]��9�y��K"�ãh(�8��:��#|�3��g6���ţ��g�.��e�y��I&C\86�׿�=ţ�v��IØo�[L�i��ˏ7��2im�P������?SD.��X,�S"u���˺�(�,ث3� T�u�c��K~hG� p��>�"�)P�z� º�Q!E�Fޛ"n�{����;7�d���9J$�U��?��U�骯?����E��qZ �21w���ѶMAD���#�#F�:!��ݿ1tR�k�%��x����h&U�v�����$��(��HdR���4�~ت!ʑDw�M.am�w�21���W�hJ�
8�QIj�"o��|��'��R��t#9�uI�+�v-��"�v9^%��US;j�ћ�~S�';�A2�����g� b��[�L��T�iW�"0"KN�Zr��x��h.��Qj�c�:g��נ}"��gL-X���R?�
�q�cG����2�ŞA;ڇh��OJb�.-AG4'�jv��hkKi-Kuz�K�M��ǎ2�K�HI�k]�^<7a�5e� ̷b���­���[�H�$V%���t��֚Bݲ����=t����  �b��lSd����'�d���gB� �|��q?{l�^M������xlH������l�!�1
:w{/��PY�>Zkح�8�)A��=���*��ꇑH����"4G���'�B\A+S��|A&Za��,R�y����5N�> M�S[�����m�l=�����Ɉ4�B�xv�څ2����N���O������g���<@$�y6L稌sR�a~_y�Lk��$hb��a���bwg}�^����;��|/(��ze����� �z�2�?'~7l��@�@�/yH�:]����|}C��'9���� ��ɱH��)[>ڰ�Bz�Nm��+йR)��S݈6Z5�L�l*B�������W�}VF����� /)�c�L֛c~�i��궺�w�����"�h����I�t�*W�٫��:�1e����2<�ٖn�99<�Ko���[��&�;!޸&� \%T�o�)^��c�#�v �k*c��i�8/B��ar��e�~���S�DU.���*�MM9���y�f劗0!��������[��hRE`��H�����{ψ
4\��v�K�xg�w�[6�h� �%o5���1�n8m���	�I8 @M��]^=&�ԚQ����CT����&���d�Pc`,X4Z�c�};���L��h�:�K�w��A��h��=�<�
Q�Ɨ:�B'w��1y0�M�.�!T�
�%s��ɮk�h�q�� סe�/��?���8�;㇘g�
���3��bc{f,J�gw�2ނ�����]P2u���4�f�d�G��Uۄy�W�_׫�Pi`�l�.ڐ^g6A���%Y������)^Jґ��U�B�W#��t)��޻�p� ƆPN;����մX��o�S�+�8�r�QI���� �	�TVP�-��j5td��i�X���4�79��>�5`[8D[V��V���DƉ��8> 
��	Ώd�{�}����sh|�r�>Y�{8��������}vp~�9��%�0R�.|�\����h3s�]�%˚l��Rӱ{�4ZZ	0$m�k�p�#��Ϸ���o�py�Yw� ��Sg�h~i�5c,��r����j�W���jf�X����+D�����!1�%�NH���k�W�mG�J�N�?�)���i��k��ōx c_u�Vڂ�ٵ�m����l��J���q	G����>�!�K�y��Z���H��h?{a������^���P���r���0ԫ|s�§���d"羜�ir������.qx����gHU!^���(/+�`F[�+h��OX��W��yG�	I?h���ׇ&dλ[	�m��C߈/�.�Q�i���\T�_5~,C�7�=H�%N�������<#�W~��/{��hLlbƑ.�oc�T�0p=YNԙ+��xȄ9L�#|�̭9�C(� e�3c`��E���!kl�ݶ��z8J�o67=ٹꤩ��#b��ۡ���R� ՙ��O�a�l�|��Ţ�p}���ې���apoT5�j�n�����j%����o�Y��G��[m��-��I���z.���ӟ�mDټ���j	�䂠��v��r-�:W����5vR����~�i���#���<8�:U��ZÙ])�}x���;1���Ā��hY@3��=��Ef[�D�gEȿ��ư�kz�.��"�`&����Dv�Ӵi��n��Q^��M��M�)�M;$֨���(5���L�3�oK�TA�� �<q�gZ�~-����� �g._"R�D�/q����Y��o�Ǒ��j ����nu�J\�M�0��3��˥��	
����33��ѷ