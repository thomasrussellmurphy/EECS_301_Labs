��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��&���i} Ĳ?��K���"�`?!9��T�8���W�Ō�SF�Vđ;������W��{���}��麄��Q{��<�?@\������p|#�0ѓ�U���Pi���hw4ͩ�x9�k}A��ïq��a��A+��[�*��&C��G����8�-�0�G��$�q
f��(ڽ�C�z��������z�H�k�VAGF���02��̿�[Kj-�GVC˽�I��S����x����6��|�n��8-w7&�|�:}dM����"��u�1q�%�T���m6Ւ $�Ǿ
���s^C�*��P;�w&юgQh��\�S����49q#���.�dߠZ���J��2y�l�Խ���VA*�
R���<o������˚�R��q�.��&��P���<m�}�|�t X���(&��i�^'#�F	2TZ�$�N��x�!�O��n�I<������S��t��_�h;�"��F.Һ��ʊ6.��C����%�4r={bON�_��9i�.eOY�"�0ʾ�J�GWCD�a�?診�>�2����'�g����婘FEYu
&E�G�_�b�4��Zֽ�qs�!��z\1��w6ata��P�)�׃?ꓗ>�5�ZJf��?J�A#�J�����
,�*�4�(2{n��u3;��T� �I;ʽȧ��`��y�E������>y�DlD�Fl�	�$ps]v�g��^^Byj;�쾺�����=��n*�*���ƺ����P��n��`{D�R�4��]![}f��ɺ�����JPL	��3���2�HH�\�	�+ ��K�4W"M��L����)C4�:3'ɦ��q��MH6�e27@w�
�+���>[��t3�����/Rݞ-f��-1�V���c�'c�U�!Ԍ������k����9D
����u�Xo�h�])��<>�M7��ٕD�o��[6G��M�'�Q;�����%��lu�3�u��Dg-yV��{s.:؂�:��ح�K�S�ޔ������u�+b� �q�Q������+xP����b�-[�#dg>as�|0
���>b��������I�(F ��$�����m��p@����<��B�������2�?cQ�ﺮ�V��Y��is��ħ9X.����WM[����Cr��ݹ�]�Aj�UR�&��9ư9�Gt��vb�jbm�38$��"��6�7�#^}�񇅩,d6d�\m�ty�;c-l��tq��J҈M���)�R���Λ]Y:v7������u1۞|<�ю���U`7pڽ�a
�>gCӊ۴y[ �qH��G�!�F�o�G���tPX�^��R���:-��b��'1���?+1Ѭ�b�߼ʉ��m���
�V��w�B�F�Х����Z?�u���n"�.֎��YE����B�����Ăzݏ&��S�������P*�c����
�oqx0���'��0��[�a������綖Mn�4�!}D�X?�W�e�@�`��e��Pg��C�0���-le��܀�Ԕ��6��?�仢�R�R�7�,XLg���_�Vma�������42���Gz����id���}:�XsG��k�n�î7���%|��g�J!�'�PWCLj�
qU�m5��c��-͒�~�f�K��b�0Z���gP��U�c&/���P���w�Z�."[ew\�[cf�x:�Y\��B���]x����〢1�6kX'�	η�d~@s��J�sk������ɹydd6�@	򦴖����#?�䟻���)���
�#����[��w����S��:�	� ����o]4q*�"�Y��}�N�S�?�17��R��D�V~'������?�`Lx����VM�)�J�"�*��$�:&�����h3���u����o�����a ʱ�W��:4	��ս�q0Fu��q�D�]��,"M�7������{�4�D�y�~Z&ӟ����?�om�S�¯D�:�׈������@:I7�R�e|��:93Za����"K���ݼ��tV���p���t�v���oH��|� c����k6k=Oh����ˁQ�j܅'p_WU�00^�i�19�sq%��"H��l���Q����(�{4pc`�U+��Q��@ʍﵳ6܁����?� �/�~4��΂T�5��]��a{� xn'X��ە� -*�^���&�6�B��[8J�W���aebl�-���Q�+Pf�q�*�ո'Q$g��P��Ϊx+����a�_�e�-����xn�1����[=�r3��\��2��ύ�}X�������x	5�ܦ��,D�S�J&�E���T�+���z�	u��!�>%�rVe��N��K�4�&�~vb��"�[g��;��&Q��S���}p����8�ׁz��l���ͪ��{�T߆�Z]�M#����o���PУ9gU`�G���B�Z>nv������K���	O	��11�	�K�-(���<S.��{�珘P��)/~��z5�ܩ��#���yT��j��ӝ+�&���)>�F���B?����H&��+r@PQr7�"n8���T��<1&S���__�:�pZּ�g=�s������|$Ց�R��(��8�k���LT�V!��];&�+��G�1xT��X!��շ����u�$ +u^����(yh�N����i���lɷt������K�ňa�~ %�o�r5���"(�Q�>���*n��G;g�_��f-���4�2?��2��r^�K���6U�J�ok[jֺX9�0k����l�Ig�ܣ������a�s�垾����ٵX����� U��9gG��n�L�6��ͫtg ��a��3,Cd�K�@��q�@o{Jȯ�uɷC����nik�.�2�U��ik]걽�� ���ҵ���N\���C+yC^+2��v�G���˻	�b��CY�+��HgE%?�r�Z�k�� �ĕ]�Ѿ#6q�5̲�?��!iG�<Z�qjb��~�~�����a\ʗ2=O���_8�m{~��*��T$'xi[4IL��1C]���՝����:�d�B���E^o]�����	q;��##v�c=$��B�o.�V�����KN���P�}�*��i��:C�����a"x�KL�^��BD�	�G���Ya�Tm�>�D�?�9��k�AL��%��Y� �@�����ʧ��&��l�8��]����g�)J�]|�׬O�R�F胆Ԑ�ݓ�
ң��"68��L�ŭ����M۰~�!����o�ǝ�����*��tB1����YO�C�an��̽?�s0�J�����p�vzS�@pr�����UN۟�-�J���B����t�'��4�:�~�u��`$�@d��2]܏E{m���|Ɯ_Ŗ-D��Q$SX@�ԍ��~*~P<���mr�V���\�ޤj��u�6��;d=�o�[��>�V�;�t-|7�d���?�ȏ�g⃏a6�Ҫú�:�����(��S�^'�ʐXzT��陂M������J4/L:���u��v�l �<�43Z!"�J���HO���Ax���>H��q2���ж
�#i��(f���h�l{�E
��(!�<_�&�ʐ�
Jٖ������\pѨ��c$8#$y��bU1p޼ ̯��/,O��y�ե���"�p�u�_��"�Q�b��ׅ�Rwc��AHBa6������_�D�pت�=�ե�
�g^�ĉ��q�<�_�3HL�<�:���S�W)���;TK+Ac��iN�NmäiK�~���pʨ)�w�i�y�~��X�<n��B±����"q�z�v�����M��~��Ҵ�!�@�]�����Mf����IKru�S �W���x��d�HS0hd<$i�5��ST���m���焁oKј-�L4p�bֲg��:ۗc3y��Y�7���z(�?('&��Je4	=��Ƹl�O>�Zq�*�`���Վ �>%e��ώ��Dm��}'�ӵ���Γx��%�8�B�$��DL�
��h�z�o�Y����M����k�OE�=_�H1~��0R���u�Jωu�6�����Uբ�<���5`����5�����F&�ۃ�F����mWL-%��Jx�Zn�xt�����B4ǰ�k�T*�`�6���({#����h"�n�v�e*�ܧ\ު�B���?�LT�7ϐ�%!@�}��a�|����b��;-|Y��Z��i�SS��;�
��(	��̀2�����ڗ�9\p�4a�a�<�Td!��\�<�3�"0�^�'I����ޗHV#)A�^;��'��?3�c��Z�n�u�x"�c�HI�*�c�p�
%၍���%o��M��?�tw+j[���m�o�B�1��|�Cͳ��\)��z.�.�}7�8��Ҹ?��篒u!�en/?!�}�	o�vL9p�@uŋb�&�0,C)���B�^�Y �9	[�s3����hȔH��
@a��L Ήuj���շ��8*��Ω�����l�G`��?��nM�^���������W ]�7�\x�%�;�AS���wp��;X�پq�Jh���5W \)��N<w��ۤ}��F�l�ݎ��n�ʫ�|�g��$w���BV�
H���6/��Q���Cx���!;0��J��?yP�T��.>jf]P�G��cLP��?_���%��X����_pC�-�X�atx�u`��g+]EFC�o�pj�!��s��TC�r����:;�I,�(�ht���)���5

yKd:8��:�_�t���� �F:~<�Bk�%����,��;�$�t�2��U@b
�A��2�&�F��
�hp�;��b�5�vs��m����yy������D�k�ڟ����d�{��Zi�8�/�Psmv�%����ɤ��?�}��э�E��7����Tף!5�|oB�R�,�\�w��1�E)c�n����B�h5;K"�!���DlAI$k٭R��(������߆`I�ŵ�?Oy����~Y�nv��e�B�F��4F�3K���b�g-��f*ܯ�h����>Bn��Z�Zg��Z�.W�u+NPcT�gg���m^d��G&�$K
nsp��"��pjl��;��yZ'B�z][f�8U����cyy۠�C�����'��Q����7`��x��P����;��$�M΋4m��&2e�-?;`r]x��?,�o�)�ew� �qWs�����Lf���dؙ���b�{AoU8�~������~K
�M��E	��u��|G�5�����-��q��e���k���)��#��I�"x�7��A'\#"��79i�7�3h}l���z��C�ն;������ǽ O��ܱJ���Q�\�!ݬ v:���!HW!ڑj�B�&�Q�tq�jr�A�W@jM��V���-����H&�5k/��bm̔B�w��p[��+;~�$�}tg�V�B%p�g%Ny�m���%t-LJ�3579+Y�P���讪����4tZ;���{��z���fݖ%k�1 ��5���ǭ�<����
J	VS����#p��R��ܖL�4�$�pH/}+�qgF���q�?�Q�J)q�����w,/�%�.�Vwe����h���m}����gB*��sJ:����@j�
��
�мi�0�#X
�ˋ+l�78�=���h�Z_�����Y0BV)ʠ����d@����B�x���瀙'����,Sˍ� �D��D,�-X�+`��s_�@�JQ�6�dc�kډ����&�5�	��!�ԿL؄6(�;]4��y<���L��
�nG����p��88������@��J��YY�s���]n�.b!���{d����.�{a:P���7X��w睲�lN�v��1X�A���2#���41-��,�ִ��Kazw�^��-�O:��K���l�bUU~�Nݳ��#7B���DJ�n($��_�\�.��D��r�S��~sMTV͏7/p��Z��M�bm���_�2��ʹ�L����u��<������[�ѵ.���[쒨'�6a�1�s w��oE4�{%Iq�������̄��
?�(�Y�V%G*�P9����Z�Gc�[a(S�e�N����%���T5�����N�l�K/�z7�D��ƶ�;�=���U#���c�DH��i1A�DN�S�
���{��nβ�Uf�bʃ�X��S+��v	�]�M:���!��z�6��6cB1͍hLn<�G�<��;��w����;&I����8���)y3C��ӴB�!M���|v��4��F3�W������8��q�P��̩<T�=��p\2�i�w!�=�����"�$? 囪h�FO�2o��,�N7lhe�[���Ev'
���m�**L�n�"��q�I���Q{%3���է����>�/�R�,�3s8㵃nJ��i�W���I�ʨ5A���k(����=���c�_���'6��O H7Lz�k�������C}��^��΍�֯N��fN�,*x!_�-�a�ݞ������Jw�v�i�fI��bAY��U�G���rG2��W��I�އ�0�4z���U0�gs�$�gM"t�A�\�Ec.�����qm�p�xR�� D7ИT�=Z�͎�8
��������D�������gg0�pC���]�O��H�k���@�B7�1�T/��\k�Du�y=z��{ߌ3m�LO�S:�R!���ΗV]|{M�@? ķ��َ4CM��(��H�R
6Z���n&�x�1�_=߯X�R���y��f���$�1IB������,�����) *R���*�$S5գre��u�Q�8�ʲI���m]�0Z�?���6�u ��͂��7�d��\�U�Q�ǋ�@d5��?� q��	�	BۆB�W��U�l����nT�<H��W� �}O���>�grn��7��ӌ-]�[j�9 #��ɤ�2��p
r=���1�-��t� z�z
1x�S>�j�J̈��Е�	�'YS�X-C2K[.�%!E���ֳ��o�| V��@�_S�+A�RJbA�G}�H[/���V��W��,1��?��u&y?y�Sf�'�TvF^j"x�!���'SY?��}TV���ͺ����O6䱠�Ũ��c�E�LD���`K��,P5�+ߑ3R0��,w�����P�t��O
�Z�]��7�YClv.t-$(�ӛ��֟/
��ˀ�g~-wv���3!���)��fe���bD��4�mB��1�.�*��_
�� $�����q���>�Eʆ���qe� b�lΠ�j�s��T�?�VN���YzFG�K}E]�mZփ�������['a�콸������
����
��P�693/o �8A	��x`���8Z���6��Ӄ�ocQ����ϘT���u�y�/Wo�ϫ �*[�{��{�̿���$������3v`9�0]���"	KW�j�����f���/��-x/
o%�W�˓�Oyg|��{�W� Wv(X�9���㓃�(���ڊ��ړh�ȁ,��o�r ��=L$H�s���M0�v�q@��'��~��A�yi�B %��1�"x#��NG�3�O��\���h�>@�q8炋zR��Su��������4�)d謬�qc��K�(�t>G�f�T�V�'��ؗD���oć���Z�<�N�%�-���p�B�%�����R�S�V>f@��h���/����s����6���������y���w$����B��.:��zr,���î�)k+��9�v�>�B���V.2�@��d���/�A^�C?�A_��i?���h�|L�W���ha�|0s;�ߙ�����B<뺵4�bfjF	�h�pYS�\�o�-�ٙ�t�Gw��{��T_�����v��T�(��M����ʏv&Dt�x�nK�`�T�z��}�	�Dy2�1I�q]���)Z�> �������c�=�ky-/U]?�0+��T��k~Coj����#N��&eI �xO
"�1���M����n|d�3G+�CS4Ɏ�	�)x6D�%�L�$'3)��FkD��_���Q��dFs�S�Z&Ҭȫ�����߃�O=���O���3oh�i�@[����&���ؙ�l��g+�ōf2��8\��?4��!	��ۃ�Ğ l=ir��)u����,"<��x]l�$}i�S��,to]�4�mE��~?w�����g�!7����(7��黓�er��u��'w�uŖ.�c�x��{�
��!�O�J6���%�9�f�,�)F������<��Y1U���r���Go�����4�U�A���K�����T�R���"i��C�����X�y��bdl~��-�}��b; 4�Z��C곉ʁ���m=S`� ��핊^���R�^���`�i�-�����~�&K��fI�o[��/�[ ���rkm���-Ya�J�Dy@�/�=��nF|��:�$��-֙�شhE/����?�U�$�������.��z�Ccq/x)-���������Pk7��Ù�ȿ(8�K8K7�%P�^@tui�06C��|>�ً�e=�m|��_9��୭@,
d(kK�خ�토�@1�b���U6o���V�8ټ��I��� �$���B��[3_���VV�+���3���I�YM;���t���k2����ky�#'��@��urFL��~��A)�i'����ޣ��"�<�~�(�'��
u�r���� '�$�� ]�H� ,�1Hݨ�'bVۉh!N��x�.��%h"t�����29+aK5�|��wdI�xe�k�T�����w6�N�#�~2�L����Z}и!_�6�s��j=�?�,�zЊ�]���(�'��\g�&`X��ǧ�s+�')�ѥ��A���mz��˾+���XMa�
��4;�L�*U�6�������#h�R{S��>Kj>�Wk�/���yM�!tݯ2���W�{-�ʦ�c�]�	��(��[@��}l��M�@IQ>K��H�oaK:�)m�[��5%�	c�M:<B��6���0��E�>833����Ә!�l��^y{\4f&�D5�f
�[��:����DJ_dOY�O)!Z�<>��g��ݗ���Q��Y�x�B$ڤ�lo�����=Tw���w?�1���L�!���}i<�P�k���L��i��c�����қ�j�w沋\�S^*(ji�6�ϒ�+bx�j��F>3-��V(MF�a�m^��Tr{B���$�sA\3<mj���創8�D�a��<4�2Qb��ͦ`X�V]J����O��T-���V>y�B���z���Y��ÚIq 2T�x���_t�<�/s�#�<�k����LS��e��pă��E�]8|>d��Qބ��ik�Ф��Zn��3Y���h��*~7uV�8�Ml�"<D�Xw�'���J�V:[f9L�����ڽ�>�$��@,��?["3��Z����׌H�8'W�K��)� ~h�!¾r_�Lz������i�Z��s]��0ĥC�w8Ҕq]�D��*���� �#��Yb�� L�I��n!&ځ�I3�lY3��W|��Hɞ|���@��pܙ�qxa�y��6�M\f+�,�ƫ�@���fHn�T�Bb�VbF�:�5���?��`<f�}CQ@
۟�̓T,�K1����b9yt:�� ����ϋ˧E�թ`�pD�����$xE��?^]�
؂F(̖���v�h�R�K4gO��������_����Go6��|�W�S��x'?�vp$�x�4��XX��5�vQ)gn�Ń�a���b0Ph�wش�1�@zC��7"H���e��̛���5Y�?w�_	i��#݇�A�	V�*��x�J#��@�$�r늖?=!�7#:�=/����,<T��Ü��3]�t珔(�t<�ܹ�������44��~'tD���W6jJ��a�@tq�eT�K�.,��,A䊍�����F��C�LL�8xV����Z�\�xA`7��c������E��L���:Wtb�o?9CFXAq����������Vt_�^�@�8(9��2���qy��r�����4���a�~��1k4��}��yC��A?�k��7�V���_���^�g�E����`Rh�#��zO���2�I��2�I����L��)R������y<�%���oFb�c�xC�l6}�5��m�����O��:L�0$Z����[2����Z',���niGp\�g��f���P
��xn�w(6�<%�_��V��t1N�6ݮA�P$�^J+ʧ.�8�K�i�-�-��7Rc崀��_����?ҷ�Sʖk.��d��O���|1����|���>�g�ш�`��+u�Txʵ���.lk���x_)��r6�S�)~۔�x�$�sԑ������-KA
e��2i�)��"#�s~�����"2��ZHq���>ɨ�]nk��|Ǵ���0�!���@���h,������~�w��)�	O˟_>�-+��;a����#q�k�zvp����Lvu�1�k֒��}o�;W�De�>�!4�)TOo=�D��i/
1�0�5���w���U��GTZl ��W����"+��8Q{Kt�֐�i\��Lpᰥ�|o==s���f�S�о�4]B6�܎��[7�ܹ��I�:���(f,�80ܙ|�Fۤ$���������3�E��qg��+�� f?� ^#Ǭ�*�͂��@��.��O��z�zw�Uv������[X�ߕH'�/�'���
�5H��+2Q�jP9�_ �X�ǥL�Z,�йe6b�t� W��� �t��qt�`�]IM�H�nk���!NQ�*).|�j��a��eЎ^�o�?�"Z�2�s��9	�*�ϥ�N��8y0^���'���0��Tv�D.r�>�9��.������ˢ*9��}�mh�U�L�>tP���f(\֝�a�^�4 [n!��.Q�Pߜ���q3��G���g��^h������a�-/������++
	�
�+��r��ٖ�챷�7a��V����6�X+d�5S�%6I�9�	l�{2��(�;Ę2����m���-Y�xXmfg�Y)�b���Q�ؓ��o{��E����P�*H�
���2wD��ж�:�̣�?�9�5�ʽ����i$8�s�z!�h�V�]"%�GfߧDtS�'���F+Q�U�,>%f��81Ep��쵂�`���Q]奜��o6&��X�i�+�	/W�'��~�/�s�m�?K`Ǉ�D;=��lA���Q^��"h�D�	���[<�0�#0ģ|���x�)�?"��&�����9�5������|���0�>��gy�bu/�L��h'�Z��L�����6��h��SGD�6�a�&�S�����$��Ũ�݌q-Αm��_���j�6�1�������}	+��zz�������>�v�����c��7�SA�V^(qA���V��<����bv�E�*\�����&�XE���=����9��>��Ru�2�θ5��&љ�S�����=�T��l�,����]^�pv��R[�Hގm��*qJ ���ꋼ��y.�HΩ���A��"%���[�`T��\@��&]_�AaD����;��#+��>Sб�-���fߞ�J��!����[�L�Se@�u���YE in����*�����D���<Qq�Uߴ�f��ܥC�% �Dye����;��
t�|�Қ���A���D�>��N�K�V�oD][�ʧآ�/�J���5�v�4����=V@P$�g����i�_Z��5����`P���m�+N����R�����L���2Z�ƨ�4�����y���1����A���Nm��>��P��X½)?K�L_���!��Ҡ�����f�q�j�ȟ/�k�q�-�\��韹�JT��
�l���P�~�5?۳t1����zpM���%X̛�	&^m0����X��1������=ر1�zJ����b��{�{�O��A���Տ����	��-SEU�ʧ����ׯO�uX	\��Ct-�Q��jC>�I,��e�4(���v"���/م*Ğk[�:Vνk�ZD[q(��8�4�K^DJ��g��iA�!Qt7m"M�Xz�竾�[�h��Z�/{�8��v´��O>|��	�5��L�>m�k=f��H5}e=]�߯#�<�J�;�Yċ%�C�+4�ע�d|����48��ݥ dO��{�Y،,`�e��:jz!��'�!�秒Ϟ�$����c�A���`�4�tJ�g ����Ż�Xb�$`j>'�+�%��~_f����I��~
�c����Ί��9��JC=�`1��Ym��"���m�������|�ޡHK��Lh!��f��'r�p��\_i϶rې�����т~O��E���zx��m>m�E�UĴ�4ke�<F���oH4g��$Vܩ�`t+v8�d%����kfK��
yƷ�V:�ܠ��{���28�q�d�G�D<rr�	�>���0L�(��U��N;^Au:8��i�/�o�v��fd�ǥ���R{[pt��R��D�b��c���z��S�F�>^f���)�(�E�7F�'k��h��꧂�`��>��i^^;O��m�n�4���UT������� �5T�����ҍ�cҧ�̽� +U$����MBy��Ai˸�ږ��j�D�bӡ��5��Z�&T���j�Ϙ�#P��zw�Q�3+�Vv�րj��>5e⟿A+9-��t<��-�k� �cIU"��B���՚x*��@QP������i.�+����?0�3�7��6���I)qc����]�ڛ[��"y,M�P,M;�*����Z0ln�RYg��4-�r��(������l� <@/)Z�]��+<lO h$�.����,���&=�NM�~�^����e^����0St )N����j$�Յ�����K\	��I��%���Ɣq�T����w\�$}T��ʵ����/i1v��y��Jg	m
Vل$s��ǻ��K03�*��]G_����8�>YQ�M8�D���R�:�ǻ��64C���Q�
�#j߈���f��p��N����W��i�(jY���@|��^��X�W�B��K���a���QWU8ق�T�C�t,�^��~qO�>�D�GՅN���!J7�8'��'%�=�P�D�i�ޥ��Qw��	*�Z�i݄y{���\]:���ҙ-R���"H����?HmÔTo��Ǯ?���I�a�nD��`�4�wRq�ou���!���y�Է��C��������.���J�l�YKԊ@�y}j̎�HF`X%�,���Q��2�ƞ�v��|���K�)>iL@���v?=���yM��>W?&Ț� av�c�t�_n���mx�fFʇ#-~-��*�A}�2�e�LhQ4�H�����+P��LJ��]����sTJ�OD����8.�'J����p�������� ""ĕ\���~�CZ��ӆ�?%���5%�<`��d�觐k���gNA�Fr�(4l��_~4����B�'lM��+�;@��k�
�G��x�3��:�9=y}��Q7�������)ebI��ѓFT٢l��p���pLS l�`�c������R��~�}�v�g+m[{�gM7���\�g3>�������Fb��c�x�=h�R�e�S]�ރ�﮹�=L1h=�tPb�@3ǚ�[��>L�=D9!/)�-����W��Q�VJ}�@Oے�E��:��B�`��3�js���ܐ��"g�̤c$,�i���R�B��V60�(�Qz��c�;Z��9�]1s����H�����:3g�5l��6��Z޴geM���SI�8�wdl��-9����=�� ������]2�i�H���R+��[�w���f�F����x�t;8:n��K�'"ܘt�9=��m�b��?�<�j��ٗӮM^Ҍ��b_�#x8ޏW���
���^)���WeA�O�78	�vz�i���u��ՠ����6ęZ_4��"w��G�X�.�/F�ܹ���(XRg�)��q��m�P��HiAގ���ЧWΎ6O���&O;����t�Ve*A�ZIm�Gâ{�HC��A4l�,��f�P�M2��A5<ә}J��u����k�f�����B<4�-��姄?���\A&����賿2S<�6��Wp9�c&H�=���91�}Q����77����y+.*��||���T�%[bU`U#�9Zi/H��\�"X)i8qVy�T��RU ?�$�*e���v��9p���� ���nܻ�"�w1�4���U$<�Hȓ?�+v>����]5�S�q!>*݉���L�v�h����(����������ƄnZ�s� �+ +�0��KogJ�*��7`�4�1s��h�uv���f�r�z9��gdª�����Ǣ�嚪�������9�-6e��H��v�WK�_�@0�25ߦD�ay�����n�j����2��Jw4�9l�� U[��s�⅓��g�CS���C�`ZcS�fnLv�A��1?pjW������Լ��2��h"�;o�ʟ���IA��D��9����T�t��<+����1"9c�*p���v��Sj��4��.�a�Y��۶]߆	_�9�Rg���j���W&
O�ˏ��fS��:
/j��YZ����P���%�����ʉ�{0��Ot�F�L�8�������b����B�����R�,�'�PYV�<���%l%\F�ʳ�$�����(LZ�I�r|!��9��U�h���b��8�����^�y�'�&/����CҎ���C����)�x������C��Z��ɷH�S1�q�&�v |�N80� t��+w,�y�iy6R�M�6�}z��_���N��ZE>XK� r>�' J1l��N��ep�r�Qv�<�'��މ뙡T�2�sG \<��d��i�B�ƅ,�"8a�T�BL�]ҙ��V�KvH$�	"1T/8r�s3�������.�����t�g'~i��)��h*���RR�	H����?e� �V'B'i����¶�K��H}���Ɨw0A�17) {��7��{�O!�a���*�"t��|�[V��=
+�b%��|q��u�ݿ �א�w��R9��k���18,C��>�)\;~�
8�P�r/�~��,/*0��o��/,�*��. Nf6�?�1@^TC1&�������"<��A{l��xb���ڂ,���}�����ҡ~ڽ��˴�B�+�t9��Y�L�#��[P�QB��h!����f��� ��Pnr���t%�����|�Q$��s����(��_M�'ܺp��:Sؒ��Za�.�����z�:�<?(=~��C�N��@���*���>���`��/�����v�Eu!�����:�.��@���m����J� и/($�ċ�XY�j��y �V��_1�bX:�=EN�6,2u8��.s��*!�A�dɂ�m�O�ƃj�)����;U_j�HQ��U��P�hWC�E?R?^��]e���_}Db�zX	ؗ��&0�`1����Z%0�������V�m��1w�l�4^�����|.���R7���n����B�+E���5�a��h���ܼ�p��\�-�-l�4Y��1�:71Va�]�0��k��v���N��!��CU�`$�qO3Bɤ���xɰ3�P�R�5#qH�!�$�մ����)6�-)7P�X�_P�ap�Yh�f�m���<�F�9eho�[�������	���s��]�+� �	�� |�[E莻<�اࢉ�Y���_p[�� ����a"I��(�x莩;hc�("u��}n��}��#�C�w�o��j��������Xf���9D9�Օ�鱍J|���cٯ��R�J���1/#��&<�ٺ9�v������^��]I���f
��������Y>#n��7mN�i��C�����7��ED��~J+�Ϙ��s�����;wՇ��F������to�9m
.zq������^�Nqí����g �8 �Ո�RPyqޗB�FG�d�o���6�x���3����|���tӘ$L�K����ۚt1��6�4&r���v��@��J�z0��!Ut���[�w`N����&&5��#<c �z��q3)�X���z,�
��y)}2��}*pm�[Q�?�Z����D�+�j>-��H�Bb�u����sЮ����m�rB��]�w*�9�����ag.�W��R��Q�P;p���q��$/�ꗠ����'1P�#���@:�������OO��-�{ZU3�O-Sge`j}D��8ؙ�]
��v�t��Ǜ䷵�_Qv����RZN �V~��v,hI�5_&8s��ǂlݯ��t���<+2�_�;V�#?�	��;B]�Z"���;���%�3{�2qC.��.��5�"2q�EK-�E1��SQndbjx�U�ƚ����R$�׺ڏ*�� ��0�yNJY\����K�5�w@n�<V�0p�	Go��t2��{��L�aAOX��H7�w�L�(T����E��.L��Wt��6�).GV
a�7̪���ާe���lХ8z}��*nn��E��
��.�A\0+���[�P�ft�!`/�5�)�U"vP���7�׽[���0���x�Kt��ӁJ���H�A�O�O�:��:r�W3���:��WBm.tߙ*Uޭ����"qVs��DYLi ��aX��\-^!>���u���_T�u�C�k���(X��
\G��
�(?�Y�d�rWG�o�NM�X�2�V�a/Q@_u=�nz~g��HM��?��f4�������HQ"�2��.}ÑL\OF�ƢU�@���Htꔝ�}���C�Lw����W��}zq��p�"P�<�¥�����@�b�F�Q��G�P��܃���($����+��]$�Ѻ�L���nI(�$��G+/�[FI�_�Ԯa��� 2?�ވ�k#���!�3G�P�sny�f�.�����[�HJQbFss��(a��!_,�x,�x5PF�4SK��߰����t=J	�J�����A�A6тv��60�,3|v�v���b��m��ڭ���sp辋:f���ǲ,5��u�Ќ�����]^�£��	�Z�T{��c]��8BZ��Of$�֘�zb�aM�x����������b�S��MTFSJ�0;@`?��1Sİv���CBQ���ɮ��˰S�&�b?�]f}]=���⵸0�d?�H�"(���j�����g୤�)�߳4�/�9:���Y�Yט���[H���k����ˎ��gB˩Ho�o�{B���kD�ة.Q����B56�e��g�mtE ����:l��M̝Ps�N%ۜ�х��q��(�d�EǤX�G�s�}�ƻX	!d�4t��I��3�w`��<���̺�бt�?ec���?�Po���S1umWih��<���M������Ds�6l��2���-��{�O�>�FY��c���1񣰇2
~A�g���
�b���B(y+f�f9��� ��_y����J��9+����{�f6.�H�A�H��.-Z�z�ȨO�y��|�y�����k�ٰ8<����F���G����N��A�#���UD��/�C���a��1?��˙`f�>#��W����<W�x���je���t�'��]�c$�`�b�˲�t����6�����C�(%ͱ���c�U`�N�E�Egۀ}�_�� n �O���p��f6��bn�ߘCCH����:�;����"�w������_. �r�Ə{�d�ʔ��X��l`H���P�//������g�W<����<���M��%�,X�Wo�UJ�=k�nhk���_}UR	���q�%�'H:���0�	p�Y�
���B�x����Jϻ�$���<B��Kh*��
�|� F��OJ�o��������LC�y��A��r�����Nu��f#<U�^`�LO�wd�9�a�8��ų��r��� �g��T��i�3~�|.U�(�~��m$}W��D���"��J�F˔�qV�5��G�<,o�x����q�W�b���[�@�o�j'���(ju��;���mw��P�5��;| ��i���S#KfPO<�.��k�D8H��s�'����$�\y�� ǽ8r�E�I}��.�6��rsm��`�?�5�7�Z̍xVn���#�2�v��O����)�eqc&l���)�4ϕ�>sg�He7�c�.��l}�	/�L|m{���8��)q����E��]��AK�b�{sH��Pj�P��.$���?��2��C���@��X�`������N�-�e����5s6dd�+@Ƙ�\nyo�ۉp�F���2P�5�~�h����W�k�#���R���(C�G���O^��J�MH�fH�=O ��v(~�O؉��R��Ձ���먔��dmk�������]/��J��k�@���������ݲK��x�q�F�.��`ҿAb�Ff�fo�\���1���pZԷϙ��3��UL��w����*��/����
���Y��*�����
?KSg�|���!�S���Ħ�~	r�V���*�bfm��>��I~7}����b�R1���S'����1���q�@-V�6U��qi�ed"&�??�M����e�'D��u���@2>{l}R|�&i8��%�k�_���[��AVb���՘���a�j}��nT���J�o,���zܿ�W-逸-~Vy�d۽�ړۺ�}QS��W��iN��+��*Ǩ9���q�i�Rn_�ct�S::B	GN(,ߒ�A��L�|���n�n�W�F�,�������;,�Wc��ɝ��P"�І{i!A�֊>l(�Oq��l���
a�[�G�J�AV�����H�ח0��"��s��� ��O�.�r3
��_sH�x��hd�U��*���?��)�3��b3�,��%m�/4�N2�]�r�̰υ���I�Q��;Qf#����`$��rD�4�tѽ��(�\�~$���eZq֓��p�L7hA(�i/&�b'/x#��`mX�<~���B�C\
�q��5�C�</��%���?���Bjp�}�ڡ)*a�@��!���q�?G<�R^�u��J:��]��"S3AfB�g��	G��6(9�r�!��I2������f�/��\5�E��.dʤ�v�����j�A���:0�hi������E��PM?귫t�i�ry�N��&����Rg�ݑ�)���/>�Y�qȹ盐�����E�%��s9Y�(��L��+pۭ�[�n�t0�TPO��f�C�❐����=V*���_���w ���]�w���;(⪰��Ei��1nJ�׮^��GB���9_s���ˍ4-o�C��/s�s�q��U�,� ")�V�~�3�{Iڬ�	V�	�<�@�B�gJX���B:3�Q9O����"����Ԍ�W���d�8N?�v�̖/��V���YN�M������,�m;	<H��30g�Q��Zl$o��ޑ
��ᅹ	$��~=�?�0����]nSc�rC��������։D�Ye���yD�ޠ>��O,=w�I=�瑐o�Q�.J�P�3�I�S��~7G;�m�XT9��S��^b
�x�㲧�|ն�8ƈg¢tX���9A�-11Z�=�L��+��2��Q������U-�>'��O�*f�]�B�|���<vʊ���\�R���ѕݮ?C�! �fr�芽3�А*�f�\m�?�A�H�?tT�������7:�A2��J_���#抿!Vt��5��ZQ��=�F謕�{�y<�\�-�����+�6��-��{��ˤ���
Ӟ�,�XX�5q3���Ԩ��Q<�9��$�v���'������� �l�-���Z"�l�KD�٫��P�;6�9-̹LQ��� -��C�X'�3�g�芞��-�K�P��$j�]m����<S��Ҝ�XօkDPU>��1f�u���t�^#�����9�ة�c�K)]��jM�2����|�C6^��Y�S�i/�:nMf:,?��7����+�� ��ʡ�a�-��1�y���j���rI���B��]ˀZ[�i���F͏�#3�����:���XH�Ky��C�ȹ�I�X�_E��C�\	(�w�H�_<��gt�T���[N��qY:�8�\c��I+F�ѩ���ftI
*�u���̂��!�J%�NV_\L��7���&7@�oHg�O�^��֪E	�~ Jn�����D,�T�i�����)B���p8}���f���+��h�̄����I�pFlH��vG�U:ʶ��j��V^/j]v�E��G�,�j/��K|��C�ǌO����r^P���p�4/m������-I�M��A��m�^��!�t|lQ��LE�A_�('}�U�V� �/S}jn��A,X�Hl�.��}��a� �K��"Z�-�C��#R�9���1�IRB���]yu �6}�1�=ܝ���Q��ӼƋ�A� �v�]\���5�n�H֭OX�`T]����I�a�_��Y-�^ӽP/��?�Z���]X?�σ����	�k2vOY�	�Y��>0�Ϗ�x��u��DSw�?[̽Ԙ<��+�<66@#�d��J�`�|��Tv }k�M[wP�kE�AV�&���^W�)���<��\:�[�P�y����~E���I�X�j뫂�i�j7~���J�II,�ͫ!ɳ��?o7+�Mg^�Ø�E6=v�5�ȣb
�� ���mE �L͹���<v��ƅN� ��=���V��J��TQ�28jEnC� ��I=_X�����w/���JԮ6@�\����=�_~�߉��^g�?c=�@�����_w�:~�I�\H~X�Eܐ�M�?FR��^C��k��'��fM�G?��`�$�fNd	+x����ۋ{�o���}����R���q7���ä����?�绉m�k&���8�B���aE����Z�G=�����8>�=O^�)�a�q\�&���Q��N����9-Q'��Nv����@�}sd�h�i�?e��:���L6�Y-�=��\���ɿ�dc;@d�S��M0�\#�l\7�g#��쭋�)���沌)�]7�|�]�!��"��'\,e�.a���2n�[�JE�,����@�SUP�������V�bR�v�!#Qc�g �p�
������1A4N�&ïQc15z"�^wq��k:?S�k�|HR�\�Ҵ
�~�J�u�:� �GVlf�LO��D^���|�'�nt��(��.����n�,��㏄�(�ն��	��D�$Ϟ��ˈ�@��O%��u^�6ѷ�Z�*�����zK��d��I޵����F$AgAų�����sr�}���p��D)|H�q<G5�� �@����ŉ�{�c^�0�Y�Y[���އ�yޣ�0�4-.�R~���*����ˡ����Fp���t<��� 6U��s�=�[p�w���B��f(��hK�g���n�­�}ȑ���p;��II�����Rng� ����Ho��Y��̩&l�p�a���ғi�E���F��@wȡ-�{�A*���g�[NU�rVTA͹1&պ�ֱ��o���!3x�Uo����ğ�����D 0oH���>	�b>����?�K�V�@4��I#�i�e�I��"�[$���*p�K�t�-�K�m�
TÚ{1��)s|�%[��*ks�4�Wy_��}��:�t�	�բ]ލ�W7K#�	����=x /e ��).8c����-�Ga��;J۸0�@V���"c[��6�+�������Z�l�����6�Z*	q>7w.�t餠�[v�������&jw�m���uAXS�C/�bA'$��#gN����\�t��}tMb�N�����Q�@�Yx,�b�b��ud�}����;`��ڲ�-Z:��E=�%E��,��q�g�����jÎ堁���aQ,��+ �i�vI}�x�y3/��9�)�YQD1[�oh�[X�%�$���CB�9,�u�w�2Nc�Χ¸�[�[{�52�&��G �t��NsO�����Z��5�_������t ��V�Y�	n�T�Eh�A&jo���.zk��8�-��AG�0W=��;�c,C	�K#�|b���Ǩgc�M�7Qٕ�y��m^$M����~+X�_y�68���G*����@2�..e�-5{p3�AK�޿
J�7&�l�������JM��[�|������o��Ѿ�;*(Kk!�~��'K�D���Rx��V�Z��ڌ 
��t�� BPK=Y���5�'���T���d@����7��*2� Q�v�,Fm�H�*�8�b�N�-��=�5� ,Lp�o��3q�Y2�������W'˫3M���a��Y�<���ޥ���i�LZ*�%N�Ԩ��b���$�Hw�$GA�����c�?#-�C���� w��� ��X�~2d�Z��&�s�-��r���4����V�~����EO��,*p8���+�^��C��h���V�o�RM��A�$��)ħc�O�BڷAg&��g�p*r8����r�X���Fر��ճ@v#d�v@�	̧ @����d�A�s{!�"��֤�T���(|rA�D�X���q_�tLY�uR!I�~E�$;��>Q�[W�n�V�"!���:�]re�d9	���Ͷ�Kk�*����_��7���}��3�wUh�c,PB	z��7.�mD8ꋞ%3�O8��A���b��T���_�.p{�R��Nv�������.�'+c4)F X!���������U,��rb���#ߥ^4*�ih��2*��@q�3*$��hq��o�i�o��h��\������d��Վ���ә	X�(��_�i.��Y;��+g?�n0WS�'�싷�5찏��~ ��� �w��4$1t�#+�Cشٮ���'=��}�l>�����qh��WX���@n�0�hI�|f77�9q���ţz�%�e�����=���闡�xT�*�G�����hr�����2�ԅ�L��S�������j�"%W����%� ���3xV�S�:<�R�#prv8��
�L�+�Tj>��[dpޢ[Y7`�}��%]������}J��h����I�M!3\�t�I:�H!�C	z��12�o����������G5��V�!U�O�� 8�Ya^���O�3�P��y1����uq��*rl���(��R��uoƔ���Y����O%RϞ#��9
D5�./��M4���\
0,���g�2N�9r�+	�NAf��ɳ7���ʒψ}oee�1e{D��_��+�j)�O!�P�G�t���|����/W��j�.�=OP	/�%�y��N~��:�}:��6(�+[9:C�>�lh�zD��Y�	m!�b-��x��RA�n50&!T��
���sQPp]��}�F���S�q���YzL�ŗQX������N���w�={#R?jg��c
D���qh��r�(( ��HThS�b^�t��X��7�y��*�Z�b@gW�؛�b	͊L�uj�-!J