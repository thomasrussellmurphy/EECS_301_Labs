��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���2�U�z�[B`�#�� 3�����E��R�=R��1��TH�G��N�����` �۠���<q��c}�޼Y%�(�"�sڙ�AӛXG�{|��AT��x�PL(�]������r�@�h=n�O�^����	�{K�*�q�a�T�FV���:`��Q�օ�H�m�Z<A�=p�Y3������ϭ�;�jHz�#D(-������Γ�Qk��c����{p������y�q�K�Ʌ&�o՗Vy��P�N�*��}f�G��g��&�W��$�R
����a��㯅�Z^<9:�G��S�kUZ($�%��]&�A��Q_�+�\�~�4�Z�:��iI��`I���E�G�&d;���;u�A���|����"n���П�d��D��+Bӏ�}��r4:җ��	���ORP�|Aua}��V_��Y��Z]^@z�ks�yE��04,�H����c]a�(%���r@Q4xOh��!�\�������{�fTD��˦�.}�IzQ��%Ns�u,�Y�,,�H�s���%��7J���H�P�իL����⚂48�g�-x*��3 �F�++�%zGvZ0	�����.m�7�s�7U6Q^/�)���e� �0IЃ*۟�������@|���*���hBb��YL�%k�9�ΏLK��C6�L�<�n����R@�Թm"�0A���9�K6���1KvP�z�d�yn��R�%
j��\&).M6�� 怉���B�~//����4P��a r��~���o��k�{i�Х�Z �%�Q� 	1�]��� �#wb�����{��]qfU+O���Q�C���~e�z��f�zSf<o���k�ݝ��lǓ��ϣ�G��9��Ђ��8��v�ࠇaZ�<ϩ���z�:G���G6�ɫ��Z��@�p���7���0�	l1��~�Dq���k� �4k<���S�w���MP�ewa>�2��y�`B�X��!1\HN��n�u��:2O�븕lR�$-P���V�c��|�Na]���%�J��$�O�A�3@��K_�����%��F7Lׄ��^d]�R	I2u-�y�n���60@jV�^�>�=�/s3vy��q�L�!4�,y�y��$�ؚ
�ZLPŧm���N�k�q���"֒��o�o� sN�Ίu���J�o{w55��uu��w��J>җ<�An^@�!6Hf�hb7J�5D����%(1�V���m�ӇOC�ˣ��XD���A������
l��R��-$��9sq�݅��eWYƌ ?���Y�����V
@�JMm�C`��;*����e��	���[�_҄�7���4T������8~��EC�V'a3"�6��q,��[VN$�C�	������}7V(��v��[��g����FW-׌�zc,7{u�Mgx�i�t7�ב�z$K��ksP�~��ɫ�CD=���E=dX�1(jz,+Ñ*$L]�ț������N.i��?2��
 ��=p�j�/O���E$M=�M;alI�J��V�S��D�W~�(nJFL��{ʄ~����%!�E���b.����$�B���A�=gGl1�­��0��/��w������[ ���.�T��=<t�?�_�������
��5�C-�	�v�0��Y.�s	|~(��|�?T�RV6���$j4I6\(�,5���)zP}�T�����f�ڛV^01Ś �x�8Q,���g%P���z
��}f���Ó�yd<1=�v��G��,��F�|����E���w��nn�ea�o46���<Mt�d��у2�$��9��_�j�ފ�u�t|U1k����
��&9�ݖ�����= 7���l������]�/�;+�^`��8!P ���ް�V�	o�<����zO�r4�0�Z��O3-����
�1�+�7�_��)w~lx�~/76��c*7���S�����ےRe䙓�4�L���/��,-��-�}��꼆���j�0����iW�M��=�3e�&�L�Cy�]������Х6X[�^:��:��@�j`��[�|�Ƿ ɶ,����*SQ�^���j���B�܅b_��yu��2 ���ב�*'wx��j�2T�q��Nk�b��V;[�·ݸ7yz� `ݢtb��\����XD�me'o\��,Q`d�g������� Ҿ�|�^v��@�%ݯ�	�^>��XA#SY�ls��? �t�دPm2��R\¦�i������Ya�Ӳ)��s�ؐ�=R����y�K0�2y�:�x~�]FCŵ5��#{]���G���[mZf;W�H����_��g�f���N��$�!9�ucf����Y9�����ex`3���a�1rW�(���V��(&u��*�y���Q�I�����e�e��
��e��b�#��m
�+U_����tԑ|H`J ��.^�OE�-}@a\,����Vߔ贖�������{6hN!!@=.��V	�sQ���Ս�@7�����I&��=X}����V�4�( �Q�q��f���|[��J�Vd����"'�փ`�g�<�`>�ɶx��Ƴ��v���yѿ=B���G�o8�*�et	��������e��vr�r�����ޢoo0�>ȫ-H~���-@�Lt.�޻UB�=�B�kjE�����(K��ݛ�c6��]��hZ"]	�X���%�'���rˇ3-Ш.��j#�+�F�ی���)����D�݁��Fɴ�h:'���U/Jt�ٳ̡4��t%h�/�Q�j ��5|ƿ%'\���,��������?E('q�@���xL�7���BR�lds�7�B��@ك�L��V�����2oД�	������A���Z��x$)�$�6�
I*��Hhu��#�r>;(�P�
�k[p�xΪ�l�R��Hּ�8m�B����ˮ�Y��;1���ޚ�:�09�`�T��u�)���d��!�T�P3��[��o�!ʯ�^t�w RmmϠ�M���(?�Uyܭ�5'��35�wΜ1_1g:uT��Jt��sWP����3�$J	c1�"�	��ꏥ~��<_V� ��O^/	f�ڠ��]yO�u��g<bEw����iO_w�>����"�{]W^���߯��ߢM7I��Of��Z�,�nv�}�5u�}e��s�m�2(\P�a{�{`׭��)��S���.4���cr���-�ƺ{b� S'���@�.p�{}����K�2���KvP�R��7.Y�����/�i_;t�������%u{.�{�e��'W��{� ��s !�
A�w�v�K{�	n�8youZ��,�ȲE[_���J�a�SH���ɩ���Z-=gҏ������M�����a[��@Z
��	y��Y������(M�
�*ƽ:e�cE|���5޵�w��]ޏ8Ip�%�z���E!��ʈ@�^�U9#R�>�\TNJ���鄫3Ǵ�mu��/@��ae%��\f1�m�*n�	C���m߸X/���k%*	V�������@�)b���?�mu	舎`���� �`��yP�h0sU<|K��b#�L���=U�09!��}�!�<�db���B󲆗���1�a��)|��Yң�'�6�n7���>A�e��K�S�b൥��:�ͩ�� ��VI�fK@�r�=�����2���4�n��օ8q��!�r@�(GޯA����q���%�{
�����B�fY�B�@	M���D���!Ft��)�����&![�^䮒�J�G����y�n�K�6m�Z��Q�ې�CF�O;�b�_HO� �}w�&*���&���#�fx�~g��E[�.C�c�4��-�b��.z�U�|N��w8d:�=�eμ額z�[m��YͭGt�B \�����Wl���$K�Y#z�I)�/�[%V�Y��(��!s�Y���@	?��̣�Y��7���4˧�{�Ңo����Z�ɤ0A����C�L#'�&���y���Ǩ�R��*<WA3"���b�i�$���b��^����qn!K�[�A_"%��څ��YU��$.|2���U͒����m-
�Г�[�8~ �/3��0���g�{����SE�7���4��H�#,�ψ�ޘ
>p2J����?�
��骚���o̍t���Z��-����U�#a��u��0B-�o�#�������,�u';r�� �t�1�f�/��ȪS.'H�gʌ�J�.'߭���t�(A���	1]��G#�|�����͊�(�yo�?]�0�K��ˠ탏}��*��`����2=��:�9<9\ׄB&ypS�2U��7V�ʣ�/M�P�֌-a�ߕs?����:p�bN��?g-3�ͩf��p��j"9��r��Wq'�J���(#�9`��	`���B}>�2����q��gH]A�P�)K���u�r��;�	�yh��g6��*�|�,C�vA"扗ʓt��iu���$}2f%���<��B�(`�� ��/˂��Q]3(�b)�����g�)��]Ȭ���2�2�����J��-�Nz��q`!�*_aK����]Du^12�ʻU�1�Tz�S���q��p{�V�{%ͮ9 �є�".���,@���{�c9�?yn�l�֞�3O�����&�F��J}��v-qNs��G�j��Z�s�6���{�!6��mDR{-o�y��y��1��W�q�{�����K,�5�of�Zf3��~w��s���&k���ȈZ��[8/4�.ԡ� s���F���p�1�@cE2�xFę�;����9wZ����/t�o�-?���g��w�{�N��s����YO�1s� eTi՞�����6��h�eq�*�7h�-1�F�W�=����\�m�R���\�<��~���+�)�;��xȘZ�װ;�VI�0�#�e�|v���N���.�q���)��f�S��,��"�{n����˩jDn���k�;]%Bw^_��ے�l�cA��Iyv}���C�nޑnI8-]��%�g�����Eָ[}>o\��u��{���׷�׵�X���{��F#Ir��r�1�,�;I3p�_��/��������{�p�S��_d;�h�G��rV�����	��
�X��S/fg^l՞Mm�h�о�/�Z�"�f\C�=ʙ�Z|�}�Vw��u���D�L�[������bfw�z��߁��f\���*�hu��Y���t�c�����L?��d��o�6�_4�����e=��K�Zdrl�uT"�d��h-Jp�!hS��4��o�3����9��zhs|F���d>Z3����|�x�T�gt�l�3A��x��x�vi�Zڲ�sI[°�F����/]Ӡ2R&PV X�Ǡa�l�K���?Z=�5"��ډ��P� �fz$#�_,��-II����p �j��3�;[�H#o2T��Qk�P�R;Z6�r:L�\�����,E�<�7!�%E�K�q�i(�����s�e,�����TÙ���>.�kW��� �K��S!c&!)M;f�n6�L��a6/��SR��g��r��ǎ�G�Ev�+�i�Ү�o�p��?t�c�S<�^��S�Vc��d(�7���z��HvD�0�+(@��N�()����"w�?F�O�� �\Z������.�����Sc�+z�"�N�QM��I��{�l
RƠ�V�_Hnф �펤2�����"B�	UߕL%�+��[�D�����-v\��u1������{�E�W��	�ɯ[V�w��Dɠ��\tQ#xR�B�z�QU� /�Jߝ�i�9��y�Bɍ✹����ͬ��nw�AI�{rI܊ydj?�eaʙ&0��A� �x�!@k���U���M#�0g���l)�aL1^E��2)�z0Տ��%�a��BLi�Ɲ8iY\*r|nI�n��Fo!��aӗ��r��~�o�]�.�!���D�&Ec5|u<.�Z�]�p��T�4�r�֌��(�~�hݻZ��<��oߡ �3�@�3���QȄߊt� Dcw��e�;M�BJJ�o_u0���I��Xk�z+���77���i�\�C+|6ϭ��躝-��V* od�A6~R֯Jd����S�t��;��7&+r�-g/��7E��vHY���+�mh�SB��1W�#��PE)�ҼՕ厞���Sc�W�����O���F�*�:Yk���&(��Ev8�����~HKxQ��\�;ʽ�y���OR�U����IC�
��v��3�ψ/�j(�	?�01��J�� �m4� A�j�\�T�����"�� �P�f�>������b�c�ky��f��|W�s�n��݂ "g7v����^�'íq1)�D��E���z����ٮ�P�+�:�����1cj��Q�)gs�!�B��9��0(|֏�4$
V�:���6��63���}�L������/)�� *���Z�
��/rl�@��<�.VR��Ђ�3���i�w�]�����N'�;	%��Ŕ�}�!�Zp��	]aF��Z{Σ��	@�珑c��L��Z(	��]FN��CC�֜�n�mu��:\�!�d���@xZv+I�q���Kg�h�W��(��?���k����"CZ�����@@1n��f	�����a�T��~&-�����~��iG��f�����W��.>T���)�-q9�EЍ=�Ɍ�u�I	pl{,h7j��'S[��.�a+� �-t�li�/%l2�v��DZ���ڟ�](L|0,z$/r�eu1�������������0V�ޢ�	�����"��D���Z
%
��-d����X��y'�`�c�9�B�`}��+JZk[Tm�!�Te�5d>j�����\3��B�'\\u`��Cia	F�%A��Ӽ?�>&��P#��H�\��F���p�cp�Mz�ڝ J��Ԉ����إ���O�N,Eo��� ԍ?�F�BN�H�f���w�G���'�G�n�N�D����:[ �!��ge����CZ�tf�,��u,L0"��/=�XA�;=5C��;�Ml��X�$�@�7��0�P�-�P�{��;ȃ�x���?�/(�E�nԃ�6sl�ǥ��,m(S���P5H�r0�OӾC0!�����B�lA$�>��!z�����i�ۚ�����D���0�i�멈x���|�9rwDQ�3�wt�U�lV���ч���"����i��-��4#����6/�ubk�e�&�������1��E��'�U*�|��=$����FK�.�rs�k��fd&5i,�ʴ�R����2 A8ٛ&�}`@�� x��
�H�� ؑ!��� z
�,G����._�`_��f�|���o��k1��w#���֖���Y�8e���Ftl���o_���=.�'�w�Υ��0�����D���iy�eh�����5n��8�4d�>����n�F<
���D��a9:�ˌ�N��_���+t���]�v�"hJI���l�BM�҉Q��Ns���Q؆�1����pI��=��<Ԥ3/�
��H������Iăr/�i*7�F��>_ބb/+>ɶTaO��� �>D�o����8�&����ҁ1���[�@f�/�J2#{F�a쭆�+���@���c��L�yD[��e��z(��%�@�"Z�g2aڸV�K��uiEi��K�9�d|��q�N�R����

�C�r��ٵiߛP]�ޭ�0�����:�[��&��3_ڐFY�����c�n+��t���{02�͚�B���k�dH���n���x�á��\�Z�-X��.�g#�/W�����c�"�^4t�|}@;�	�[7#ʵ����e����i4�f�
��q��<H��g��GWֈ:N7)QVp:bU)H�_
{�C9�>)��w��%�4-Z�tA{����ɀx�Ȫ��姃�W���*��\��do�2P�.���@WM�4����N�b��� ���8��\e��J]��=�� �y ��dCf�i+b����5G0�հ���j��0l�I�~�v�Š��ї��1����y��Jb�9��U�}���DSa�{��$�L5e���Fe@����k;��ͪ��V���j��P�Kn��صMI�ĸȆh�%.����-��]�-�F��Jz`��7K����Bt�3�_>���Y܊�mƻ�=�b���ͧ�w�`z�.uR��'�=�[N�1Gf;� �w�-U\K!�!��/�b�����{���_\��LZﴃ��jjg�F��Jn���k�ƪ�y������64ق��~k�c�}����G��.Q=���\��lz֯meU�[���r&��#�z�2 2O�H�!�E�RK^D|�;y�ͨ���)oW?N��-a��v��<ћvK�8i{oȅVP���Xc���0�O,�;
Bd�����&x�K�1�_%pljj��Jm�u��b�5��;~^��ʛT�ø�����j.ђM�>���n��L*�X��eXN<�[*.�����Ī�R3S�\Y ����!8�'��i�wG�؏yyV�2��D�%O]q�(6�Lm��x����t �Ek��,-_��4os�bWL�c�l��Г���/[;��J=�կD���h�`}]P����U��v`)rz��R9�k���ro}P�u]1�&�#�zGY���T�a<T�&�~� ���J\F�V���R\��8��N���A�;�z8d��O�t���Rn\�U(G�Zq�=�G�b��- z�vc���%�.L�G���C�Q��F|A�W/��GG���4��ϑ��׻��k�^}z\D��y�	Eq �.���ǞӴ�	�s�ýQ�	�"��T�S�[ȉC�Ӆ0T�S�b��+�}��l�V���O���2+�YC'����H��2�T�'H�h�eZ�^�Q�r��.:[ 1"�	�n���HA��Zrl^lva���]eC��K,ye	! �r�	V2�0R7�}��uv^	>(:�J���K�-�t��<JUx��ח��� 4��\�$��0�j�ꃷ]l]@!�Z4z�rJ��n�c8 EZ_H+��;�����v�ŧQY����Ld}X�%�g�5�h�u�'G�7X���d�}��gAFK	r�'ܖ�V���8�հ�|�x���V=䙍\2����8p�p���*~�Rt.��2�l�shiR�+p;o�Na}Z�<iH�L�|���`�5AN�o��b��V�0��q�����=��Բs�-���z��R�7�����#Sܫ^eCH)�L�yy�֑N5�-�0 K�#�j�4#B�8F��ͧ�c�@�d�o�irf��!��9�J/�zXbW̆��8Vl�)L�Z�9�;Sa�Q�$(��.����Q�ю�<�⴫xP4�лt�����dD��g�wt�d�k� �/�׆c�5c@�;?䠧���K�L��mM�<_�c�}c�$���H�5V��((���^Y�:M�����}� �׆���+��O�3�7DW�+��8N�|T�����;��8�EQo����Da�w��/dQ3v���볙��u�� O��/�K*LZ|�&���
g���\�-��L,�2F<�$,��[�$�Ge5��0��4:J��4F}�X��u�PQq�iw��`RJn�EHjz���t9ê�-kXA��-�s�k�:?�������ڛ>h:ƶ�%{S.ؐ��L��S�ø�4k<p��B�ee��b��+��\f� r��Q��Y����pd�Bΰn�"BZ��3e�	��HM���I]�g������.��BO�<�: �[P�sJ('�7׎��86�D݉��&��z��%��{���~K�@��mCI�Q�@�[�1���CY���Q�o��B��4��h�h��f��V<Cl��a��@5����X�S��tAޕ���2���O�Z2	S��ڽ�|����N/K5޷w̯̃���C�F1�v[Ō�(���%�=6�H���� {_�Ng����(ݦX��Չ���g�Q��;1�a2���O�#O[#ZB=$86Y���0
7m��^,=�Ғmˏo����<n��h�|�����2Ӛ�w��,�c�
e��&�d�GO�N�z�zC�XX���;�ů��������������$���Q�P:LA$!���I��@��+N>L�_���P_fx�h�gиL������6j�H!��Ķ�*����/v7�e�bo�ˇ�LOV�iOɜ`�*&��-�c�wR�a�[ۦg��u7�0G=c�N�������x!�/�Gk�����<��x>ke��&K�'r�6i^�VJ�T�Y>�=8
�G��hz�+:1R�a�����"�E���@$$VXQ�bzx�a>I����b�˄�j�Nb�9���ؑ\ʳ~3IJ��Tj��yѯ��!51��p�_���Ŵ��g��ۏ�dL��.b�#c4����N�"n�X�V?�O�@`VY���M���ҥ������^! d��(��>�J��;��9����@ �XO�?�,2D����|�t���g+�)͏# O=��}���ӵ��%:���K���ܤ>d�O���������u����w��eR����ߑ(9?�9�,:�����[v�
�M�st+a+b��`�m,����e����#���vо���yӮ����3��i'F锜��؄S�"z�.
MV�={U��������8���
�^����s��p���=mRf�tY�D��n�gj��_��ʎ7M3��e��������`����A�i4 �7h�Nh��eU��%�w3(��$qq��.!�7ީ��j��:���I0�3*���dsE)t\w��ĭ&3v$�J�Ak�:Dp��ɴ�<	m��2�Wǃ71�������J��A�Mw[��?(Be��`�S<怖�p�� �<4�D�zek�9WR�+F�p5��}�ܽր�d9/���^���{4�Te�q`�mR�!An��B�Bٓ2�!ۦ�7�%)Lx[M�[��^8��^�🢏�MV��_�Q���XM��P꺾'�t�e��G�6�̔ӱ�/W����E/�`��I��O��%pyV��S����/mق`>}�bxC�T:k^���
9����Z��s�bQax�j�Aq���	��3rA��u'���.9�QI�G�X\���{�NR�f�`�N�(���t/'~8kn�_�PL8^��� B�w�'�������L<V�¡�#V���\�x�^Bo���وw�CLa�Q��DFT� ���F���`S�x�s[>
�������0d 6� ��[6z�X��{��]��#�������:ڻٳ�H�pP���gБ��0�����B�益�o���U9lf����ɻH�I�DcJ�j1�Һ�g7���LɁ�
��g]B(��7.�Q}� �z:�)�9Oa�|�7�U���ڙ:JN!rƖm#�j���v|}B�Uح]>G�S.A�Q�����#:T~ᢗi���ri����f����F��&U�H#�,eR @.��� Pl�-�:���~�H�|�r&��&bAm�P�)>�W�&�A�_�TX���uASe�T����&ܙ�q�δ�Ǭ��'����OAMW�X���Bs��_-;��#�]2�!ws�n#/����pB%"��e�3��wgݜ%^��&&q�{ќ�L��g��r�k�@M,�����7ɿ�§� F�7�z�A���aO8���	@���+��o,��P�h,��e:��زޣ���[��R�9̧͞�N4��Q�ų�1�Gy��)��|n$)g~[2�S�_T��G7V�X�ٯ0Rغ/�8>5(BW�o^�x�����,��� P7��Ϭ�	o��+򩮮g*C��AP�����Nz�s}A�����0��%ܼ>�c�K�S\ԣ.s���N_�ٖ�"J�� F��pBV���>&�;O>�4��Cd��)ut���v�ky��V$��(j�bK��x9.TF�(�Yz������bC�k2��������qGE|�򺪹�[�AM4�$��j������F#1H���W�u���������n�Pݾ����b'��<���&Ǡ^��0��c�`$v��_���Y�@��<#V��V�-�و��SP%�H�6Uλ䄠f(l�v��5��a����k�r�CU
 2�-�����ݝr:P���R$���t��j�j�ovw	>xb!�c��DNv�?�^�]ԛ�J���`	��q܉$�(gH�����&&<�L�?�kT:�m|���c���x��2���O����iC�8}/�EDQ����B�a�Oq�>�5`,F0�)QS�i	h$��Ju�_����}��]�-[�bb�{��1K�=bfL�m��jT�ȫb��x�ߨ2>h�N���"�Ox4!ZXIb�c�kg��O(�Nm�u�b����;B㨴,�	��\�}B�o�F�YF�I˾�2��~�OO�Z���J�B�*�r۶��1_ƅ}I�L�0Uv��g�R|�^�x���Gq��A,��"��Yׄ��j��8�c��[}z�T���%!F�yXR6�m=��Д�ID������q���R�y76O�د�"���|�6�7C������y ���&��t�M�$�Hj
uF��n��2��v}E2�����R��Vۥ�H}��E��$8��@�قڡ+	r?M֋�?�v v&�#�@%�ڵ�"q[[H�O�KP&���W��|j���i0_|L���뢻�M1g.�b���»���Y���ձ��(!��p!��w�&=�ܒ�R�(Z�^���{"`qa� ^�Rx%A�T����ډy:�F����ɻ����^���n�p��Y8�B����
P�������Q��0=
hF���K���7q�;�s�e'ng1J�G�Q���&�K�S
���:��3�՞X&Z/��:�E�>h�i�{X�F��.d]��f��v��׼�7N"��O$T��r�}(��R�!�O����W�����y^�[:gR��q�%�V �?����į)��wX�h���� �t��!�&4�ȼ��o��K@�m��1����5ӆA�	텵�L�-��i�N�4Ǹ�߶1�4��n�W�ʣ�FI&o�uȻ���$ ~����,ﻀy��o�jj;�5��������IlJ���
�q�4m�~���:����:���/�D��1���ӀX�e����2(~�i�Cƶ�4��gJ��nZZ�FyEKʑpͥ9��6ew<�=m?��ْ	/�����$d�A�7n�v S׍�N�w�};7��e@�QB|+�< ���d��a`�w��AY�1�^x�F�!ǾW��������bĒ�x��T��i��P���0g�, F=5�B���m��
�S]�ѐ�x@H�����fL0�NߧB%V�0O���e�˘NGؒ�W<����1g�JR��$@���j�l"��v �I�me�+x9L���t�=��%_/�����5�dbyO���D0T��tH3��z$a�,�N�o�M���L�]jM��Z}NU2'f�Ɛ3�;�Μ�!O��mZm^���'坛�g�'"W��II�|��G�,:�3�Fr4	{��ISR=�֔�C0���{�͵% ��rk+m�О�Z�h>t6�P>/����t�ʅ�����b�$u��/����ڹxzy�d�Kkɨ�� U��b�b�&�H5n�K��Ӻ,z�+C��X��0J�r�
��� �����x��9��g>"�C;�V�ϓ�������Ku��v�<����#����2���I�`3+�����x�t��s�qi�J���~f�-�N�"�n�ķ�T�����9��QS4&`M���e�^���%P*�� ƅc:x(ls&nf���7�Ȧ�W<�TL�`���D��5=�l�c�L{t=lm���A�`zC�n9�ήZ�����ža�5zi� ״U�_N��`�4;i,�`���/j��%x�G��R��G)��U��r�^U!�(-���M�ط� v�\G�s���,H�2�	�vV���a��X���nھ �a��@mQ�b��<�o����C+��ID�����|��9��/�0
3@��,B���6�I�Do��Lov�/0E�x)����dHS��b��\�_����k]����Q��9p�vߎ��Ƥ<i%h>���	�iz\�ؼ�!���7!'lk )��ЮZ�%X��^�[�d���FxJ���:/oZƿ2Y����Z�?�����k��o��ym2>�\_":t�e��hy�l�Dʄ�[@"�A�j�'�wm��Mgc"�Mn6�_ۼ�����A�[81�[(ӊ,�]\*hҝ,�@�^�=<�:
�~��0��������y�[�i��}���@_����
��(Q3aLn�q�x�ފ��{M���i$%��Dm?�j!����1�O;�K8z] 	�c�����1d`/_v���y�I������m���#��(�&� ��*A�:6�~C@+s�Sʋo�E�ken'��c��������\�Š�����������c��Bҗs`��18����.҃b��wq���g�p���J]�U�e�|?��¡���;|�x��}fv�FJGnA�����>��(�Āeؠ4�&�E;b��(cΝ�	�,�M�G���`hsx����xR3���р��v��a��@�����_�1HH�C�� ����E�E��'�)�8�6] l��ճ@0�3;l:����ը�;w�#"�!�x�+����ֿ�d{��)�K�Z�������Xҭ��w�D���<��燝O=	o�����1~��I/�S>��-OL���]�7�{s�K7����$��CW�@;�Z�e	�L�G�D`�(˲n�do������x�:�.d�@Fr	_��B����	{~N�I���ʶu�<l��_$����k\��l2�co�qY[�z��x���d�>�����t5J2q�k�oTՙ�.Lx̩�_���u|
�q�`.)2�>����磟��r+�Pr"A  ��RL�b���)S�Á�`��^�d��Yج���쁦10eA����v�
�����ދI:��O�+c������]�8=t�RŨ�M�ZV��&#@م��$+����er��.�2�o����d��J�#�&�T�V�Ԇ�	�G�/���p'�����|��ZX9Qۮ��>�.:���Y�*`�[ق�ر-��i�ҩZ��p�E�<�̼]��ѷs.�^��#�:��oa��%�`p�﬉G�j�E#�d�*���Q��$��vi��!���`�$� %����ީ s��=�ތ� �A%��z]e�0��@�C�"��#\砗��\S�y<��/����(�9�u��;�JS��'�W�Y��V9ي^f�:����
r�%��Oi�M\aK���%1�>�8�V�H���������+�0����B���}<���R�"�Ո��}2|����.ނ�a��Q��q!���Q�U�!(6_�H�����9��F���Q>\��PK	ֳX���<,R���0�5�Eē����/����q:{�^�e8z��K��=Ԣ�s����`;'1h�6�2��|��T��cU&���!���3�=�����8t�v�L�j�9��OΖ�30��- �$W0T�b��Z�N�!5,;i�6�A�b[)4�E�+��6�2��2��:��w�,���5֔�z��?���PKb+��r��(��'@����J�$����µ��w�2�7[�#�s����\<	Q�6�������O��F���]P�љ�g[ŝ��[����8��.�(E�M`:S%hH�X��0��C�^�2z�\��	�=�񣿖^�&'m��q��\.��~�E�G߿b�5J1`t�cS:�6�<�z{�f��K�{��D�V��Q.t")r}�mO
��͟�fE�#D9T�q��JnS���i�\�4$
�	�&`\hb�fYL/˟��u�fw�2F*��|�б5��\�ܖT��"-~<�C�+`�O��Eu�������/��,"�E�<^AxU��Zud���R"n`��rJ�[����yиpk�s�HAʾ�s�����X��'�XkD��4~' ��E��'2�9�=i	����Nk���|���sln+3��i�YD�V�^�'�,|u����â<�\A�7�U!��� kB���B ��+�]�ύ�9�'/:J�5j�]���m�Ea�^�٬�&eH����y��	����s���sSC^��yj'������+�Mh���D�"�2 s��;dL��5�B�JP�ӊS�.]M=�����%�攷�fKƽ�jc���<��5l%����k^�>x�ݡ�dP�]�[������H�!�fc�Qp=z��Ƥ�&K����|fb�U6Tm�8��m��L���o��D����/Fz@��^2��\3ʼ�*p��ˡx���!!��}�>�0�z`^?H)�|G�7Ӕ�����P�x��)w���w�������[ۻ]Ny��$��r�'����Q	A� d�׭^�(�N����c��*;*}�Xn���d/��c�9o>l�YT�!�xZ$����0���g8���q2��^�D�Z�	�	�$�f��$6�=%�CP��N0�S[��R=	�9���{?��\�5Lw�d�w�d�\�J��O�<��j�����7��G�Dk�p��S�������U�wq��oCCן*wM{I����q����,�G��K�Lz{7I�m��P�L��t���������8��B����:�ň!�th��"��tD4L'����<7b�4�(k���z����a1�7-�K[�?�U;OfMY��T�/�ܱ�Z���}�����îQa맊z�~�ےs������������w3n�
�!ӷ2&�FJ�I���C��'�#ژ�E�զ/J�{$^�j�M�'��A�����1C�[�.x�����7�hxm���l�p-I�ikM#�P+�f,�$�5~�	�����f5�y��ȼ��t�[�k��������ڷ�R�8�&0���a�򱓺
�]�o-�N.'��t$$��}+����������vϮ;k頋�u��.]p
����{F0=���[7Z�&ù��q��UŹ_�3���P�	�&�Cu[��0,� 湺w���E�A!��tR�Uc<�`�:������r�c�	�qb�{�Bމ��.��!r�i�����ɋ�C!& >0�{h��RT�3�����Jt1S�K:p�\��ƙ��`�_m�K��Η��Ә���㶍<.���Κw�
���
��yԈ��r���h���:oǳY�c`����+,���'x�$�J��\ʓԑ9��r��U?>[b�0����\���vV��ކ�#7��u��:-!8sl|뻚��G�Wpk㑍VV+nt@n�p����]���$vJI+�!��?��B��=l�o&Y�޴z&O�'�NhE�?3�i/k� H�$)��D߮]���3���"ɋ����q4��Ao���:P��{�m�qz��f���c��3Ѥ�����C�8q	s�A����~�;��*�wO�j;j͒��Mүx���>̥���M�,��;u5�+ �$�aբp�p�6G�� ʠZQ4�N�sy'��M���w%7gn�:.szM�t�h9#PuX�.�XYTM �6�!҈��W��E:�H^Wj���=�Y�3�=����Á�AOj�p6�:�8����kq�X�l>��d$B�_����,$4<��������:n���U`
x�x"�ht00эɘ���={م����郾)���+ U�
�e�T�5S*��\� ���~(�b~>��C_�G��9����E"l��񀄴�Mgҕ�B[O`�g�'}�]n�2ah�N���^�!����@U��#�
ԅ�r�#VB��<�%�Õ��Ѳ+��(ҹLC�և:�(��oըh�e|c�&��A�R�h�a\(�}qO�����������
F�z��H�@����n�œ���/H"5����]�E|13&�uaX�����J�=2��
1}�HT� �����>�J0A�W��ъ^��d/m٘I��l�+-�b�#��n-�q!�x��x}��'HA���G�Uq�_�۸{��`S��:�]�Y�Y?.n���3��V4�-R�����z�;#�<-�c�!ưN ř���������L��q�x��c��1r*m�i�`,�Έ�N���"��p�I+����+�Qm�ۮ��r�ˏ핍t
�V��h�Z=��-�(*�82���>���!�=�pz�.u���2԰V[��g^P>���Y�^[����k&�W&���!�L��+�h>��FR�X������t�Sƽ�o��)o��g�Z���^s�pil(j���\i��v�:���G�b�߲�d���]��!�JM߳�9RQz��/��G
P��?4%�8R�h�K*m��3�|���G���R�!/EJa������e�$�09d��Zm���.[��	,^2˙�I���,����|� ��� ���3ݨ����ۜQŜ\'+��y�c�̼�?9��Bi�y:�����Lc�>�F�a.y�1�`�^��o)|t���6�puS9���\ G���
��K~-��S�tw"N��P�[DǫR/EX�;�� ���/|q�m�w��,���/�7E�F#*�J�����`J3�nD��-���Ѣ�I޹꥞���kh�a�M?���Q�F��w��F��b�8\u��%o��z�6ɶi�3j}����~�W�j�H7���b��w�=�
�JIE#9@b	���T�®�%��J������*�H:Pdm�AP{��F��75����C(A��q�����MT͌�^:��h��-W�#j�}1�sL������Dn��o�E�l�� |��yY������w��˲���a�	�3��o0�n��tK�bD�G�O%&��w$ɗ���}H��̘#�J.�7�����)��ı�3'��U�d�m�6�:<faF�����W�/����0�0Ddސ0b�tMy���rPr����T��	�Hzm(0`�/�Yĩ�<z�ٹv�93���U�p�:ϋr)�Y��t�sPU�庽fZ�_!V���_vFN�=\�����,i�Ѹ�#y:no� �+�K�� �V�	d�T����B�#����z]�l�U���k]B���Y������'cб��c@ߥ�qr�(:�A߈09�h-0���/��ܜ�zo�Z��V�W�-X�i^9�M��
���
�F=p��	�/��Q"��������1̗�B��+�m�)����)ŷ(���t��_;P\�2���K��<�\Y�mָ�t�KBJ���&�3�@�X�"p�Y�C?�n��OiL�?Ֆ��yӋ# E<����Rֳ���/z,�_�h��B�>�*ହ=�A��H[8'�~�V�:-�zשY,ҿ���29uบ|j�?^�,��&���	���8{��c� ������5�c?!��,�!�{@��g=��U����)�FC<ȿp�FR_��b ��?K�WQ#��"0g	�`}���g'kf�I=�S�y�l$i�y|�v�(O�ݤ	�Y����mF�+S���'��I�Li0�<���X�n�5���vc�*�,��]g[�j��!��5�����ma���^��ۚ��7ǷJ�	������L'��s�����G���C�:��*��Jp>z������LX(w��}n�[��yJ3�6�)���M�@�|�����ٲ�q�ad%�@�[����>-�"�h�,֌9אɤ��\Y��� ��B�K��\���%������0�jʲ�/�*qS)=Y������0�d��)��"�!
����SV:�L���!f��������7F1��MZ��I
�oQ���ڰ���ji2i&\��Z���ZQ�?�"��`��QmiRqn���6�[�V��O����V&��D����q뉫b9C�-7���
�G}�[G����^��4܄~v���jo�/����W�~ �o�YF��b�P�����8*�!� �[�c)�?ٙR�_|J�ub�+U�)�Az�[+|��}���"�S!՜�3��C��N\�j �,5�Z��-����8�8�6		#B.o4�R�$��<$�׬)5�XF��Ħ�a��/�XltND�QUGG'CD^��!����0�V���ִ��x�C�"��E

��=/�����)2�쯪�v.�Z`wK�3��O^cq㋔���>�;j��	G�~�5��p�-��{S�|E�9X�emȟX�f��U�i}�Փ�Iv�f\b�M��a��ߩ<mޚ���
C,��9�rh	<�P)���� �(���l�`;54�/OP��c�v�?u���\�F!��Y5Ա�+�&��GE�(�3�.�� �/Nbiv�pJ���sQX�SL��{.z�(�ͥ�7E��Zl��8|m��p��7D�ȳLc��}�T�]y	Vqz�qr���W��c�o�َ)�mߝ3�XZ�����,D9V�g�,?�\5 �n�	���#�U��8��W�;���᭠�ZhA+��X�`V�Y���+m!^��#[��\��U��DNw�J���4���@tj��|iYL.�N%|�s��I�SW\�U����A�/w��!��/b�[]ge`C/'�n��|��K�w��á8��t�_������r�&�?R���h���"s��^�o2�)?1�&�o��T���J��9��i-o"4�# 3к�܌��f�B�{�~7*�2�>��YqaL�]����I0N�Eס)YqyO4(�S.�3�q�6����=dlZЊ�v�8k�g�5_�T1Q�ڗ<g{1/��ԝj�h}���%g��~ ��Aqk{���{�R��j�:��d�����&r{xcq�K-L��د��o�6��)��\���m���t&T�Vs`(~Z���;�"����k�fp��[ܢҡ�H���!3:���2�2,�+'�:X�ওO׭��r��_�
\�-����g�b.�R�n Z.����������,`�����&����[rm�v>��:*!�d��G�4q��5��� u$���{�ͱ�x�b�6QS���0t�e���OV���۞�T��e;������/���5�'NLL ���Ȑsb[1�W���a��l/d)"Z*̌&}W���>5u��s��]�}���R�� hA��#� ����2)tT���oE+�	�쓥6���V��?��g��	��߬H#�-p\[��w��X��9>�?A'�?���w�`�78��/}��ce�Xd�N'�&@��K1!D܇�wn�&��F�)�N�<�)�F�*V�������euЅM�b���x �]j���ҙ�t<0a����(^x�t[���0��B��o<�:O�1^�"�^	���́�f۳^����7 -�W��:��]�ɕ���d�"��L�{z�%�5�v8��f����ݣC�M�8zkT���H$)�ʆfl8ᤜu� ���G��16>��s���""x�}n����?<XN�3Ua��^�mdc�.���c�4��� Z��PZ��e��������)���J�r�:�?����-����u�*�X��93e��zB�4)^�.&��n¦0w; ��B�B*0���}Q��jX	�����8�y�u0����OM[�!��T#���]uR����i�4o3���@o+�ߑo��ߗb�Lr�.���g?�gE���nR=$ �5��1���	d8�cq�iX����w��{�	���a�.�/�0��c~��:�/���#H�t�c|�k~���B��jY�%�#X��1" ?�N�V�Iۨ�)24iq
Cjb���DK��
���l�ca[q	�Ns���/ϸ0T���NNf��w�1D�g���*|�n�
�3�L!Z�:�j4�tA�d�N��o'�s虡�r�(t~od�Ó�k�=�	-�u�&�~�%��n
�"���G�b/ɸE4�#�n����پ��m��;N�{�����v`�E"����{a����TrĞ�p���V3@AvN�ػ	���p���[��k�� ���#�w�� �����D�G�%�,�U���u��T?���՚�SF���g��V7`	�I�/��)̙����K���-�,�dη���(��Xi,NA<�5�(QaTH��t��e��<M�c�2�Q-ʇrgE�`& mᯢ�$�*��<
x�����zX��;���;�,��ZAԩ�E��/t�ɔ�X�O�\`z0e=��pa݊E�H��Q��kLj�w-p��j#�{nL�� �w	�˜S�ŀKB5NWujm@R7�J�K��!�HT��׬!�v��%�S�ǩ�{�1�3o�2�=��3>�&��� h���y��� �2е.�~;<�k:mSh�|�GmyE���cup� �IK ��;�ᘬ�l�@���~
��uE0�[�.�g��%[�F���4Ϗ�do�aaY�Ni��n�T�7������)�q�b��!����|�4#^ %aV�*՜'P���u�	�U��R��@�	����_�QTuL����A�xY�1r�e���;�U3͋ɖLD�2U���!�a�I�/m#�z^:lw��h
?���A������.:E�Ι�����`�A�z}M|o�̈́���[��$g/$�Z���`9�c��i��b���b�U�~�XJ�x%c&��K�v�V�o��0�3��d���Ʌ��b��uW�SJqֵ�}D5|���D���1RE�)GC��
���^��EG��݆Q�x^ӣV�j�%�#S�a�Ko�5`���²w:���/lp�]�ؕ���X]w��{�0R� �n�u�Ɏ3����#�(�7'�a�a�r;�'2;� ��L	mp���긤,���#��^�Ϋp	�����M�LUK��CR������^?�(�r�����Uλk~G_���P� %��q�����G�4*ۤ[�=Vi��7�ܿ��Rמ�0@�S���W�
�%�}��V��f����1�O"��P�N�*���9-�����x�W�Et&��@y\)�G-�A��|F�qc���f�l�
�,@��Q�^Cg��-���[\P.����)�U�[ʍ��'S�|��$�B��?;�y��fU� _|j3ɋa�V���ap '>6G<f߇�M��u�uH6���j�I��nW`J$���o�`�����;J�Ssd��(�ͪĕ�ʨ)�N������T�w��=�|��e�����5z#3i|z���313$��u��fǜ~V�K�d\��QK��yo����)��n*v���O�U��	̭�~��r"�w}M-� 7V���k�޴�vɧ�~UՋ����%��ϭ�P�����i[$�+�p��u҇�K�.���z�wyJ��~�߉D9Kg6�x��?��"4[)�C��Ze�yˎ�mpm
�$X~��Q=�ryB�d��)J�0J�@.� ~|%�l��|,�;B,B�ڏS��lU�D�1�Ҧ�\�m�|3������Zr�Z,�*KY�BF��|>�c����S5P�,�'	�ՠ<�(^�A_c�R1����|�r'X/�e��r��F� �Ե
����(J�?;ƃgfz|���&t T��6�4`֟�)�M=󟼒��[ ��4Se%G�����2"�1�i*0z�2����?x�پ|�_����E�����T\��qT�h��e�߮^&)F���1#��;��vԸ�7���������0'ϲ� �Ŗ��O�v*���.>�b�M�c��ݶ��GKBȄG�;ՎK�^�awd]/�/;���O��>�Z�4��C}�~����?Ę=tz4+(Rz�H�g�v������{F���:�M��^�U�g���E"|�����e�37%��)u�ju�)���ؖ���m�dq���Ĥ%�m�6p}b�hy���q�9��8$�&�V)3���1X�X~�8͒��:K�x ���S�[đ7�hv`>��h8�ˍ�.{j�)���8LꞺ�}�6�������c��#ka���|N��`W����j#`��Ֆ��N���Y,��� ;���TIgQ��:Ԁ��¤� ����nlX�ǀª��G��sEԯ*[�v�U�1��y�:��a��c�A���}�?n�sU{BsCe
'�~�y�R�����S�pk`��C��p(�c�9��O:$��	�T��4��/�X5y�.j$��]��*��-�(�o���=�4Ϗ�xO�H́_�G�$c��ف�p嚽ϣ��������u�8��Ṥ倉��H	Ggu�4�	�P�ُ�Z�'ibGgÈ~l�j�fJ%}}6�umX��b���m�\p�ȑ�yuF�A��s�~7
�8��ꮟ��uP+B�pҤ��Ю���X�;Ƽ!V�eJ\x��Zea����JBv��ܙ���"֖���Y�D,��E73�|����Q���J�� �C�Cj��m��3���H(�g�s�vP�׳��cB\��'v�zR�Q�����o��B�z������)zkyۗ,�v)���఻Z�P��r�I�XI���. VO��k��P/(�1�
~��OP�ϔ>�]HG�n�b��u`�䈜�+��.���z���������?�_6o���)���v^_���m�!%���_�H�m&O1�k��{���XǠOJ����l�ޯ�]5�Oy@4Y���4���C�&/s���5��v(s�i��O,�S� WN���z-h��6�"�}���E��WA		Фgǜ�E)H�ukm	�/�{`��)�B.��y�v�D�� Ю}��w�5��SS�2��:g�������',Z������4H>�6�Uy��<�+!X�Џ�%(1�����H��K�lj������(�?�A _'0D\�-]ɡJ�]�i\�G��2A�8k���9��y{cQu_v�M���<D ���ͱ���Q��������ױ��j� ���!�cv ���o�ֹ�S��ϲL�C��́8Q�|h�/���qёinx��tϫ$lǂ�6%�j��U*~c��<����܌t$�z����e>ۼ6%��Ù�AͲH�L�I�a�Hq��)A@ >f��#�[��~甛��b�5��H��js�WW$M��w�Q�?��������t�		k�v���<����4��ֳ��r��>��q	y5��:U$�Z�
V#T���71�WD&i¦�����o rA�W=�T���%T�&�|?ȭ�χ�i������x�^�Z��I�=����m�[���x�?p�D ��|-�Na�+}��5��*\�H��S�ʊ@� �Rg�������X����`ݧ#�F��f��d���&�\p,��jH��Pz�e�)�zj�QQ �?1ຢ�����j8mӰu�.Æ��/t������p��S��}���KqO���E��P,���������;�!U"��	6�dq��d�Vɏp
CVI:Dw�<�#���4��Yׯn�9X8��,�ly1'*𩥪����Z��Hf��מ�g�!A�'�KWF��f�Wo�t�-�,<�'x�A���8�%��
�<,�۾�^ؐ�E�d䢛��)���;����R�Y�5H��G<İ�_[h:�X.�`"�g�����ˣA�ihi�  1}ᐸJ��m'��&��~N��ZY�s�F��Y�£B�j�k�
�	�$����<�x�/^��yᝢ�%;e�z�)҆����ߙ��' 8� �Y�����X�RVs�q-�d�������6HX�i���N=f`�ݴ?�h �E{ȓ����@<�-������D�f�V��o#��̾'�;1�t�oc���S�p���'�q1��3��pV�Ϝ����l��_IO;{_�!o�������i��ߡ ���|��N���E�������K��֓wrl�I�b��ҒNt��i���x�;u�L�}n$�z�MG�_�ew�_6��T����f���u�,��D3
�:���I���AP���ہH�Q㝙�I�*���3���"�
��p�,;G�����C����A ��CO%�Ϣᩄ+8�M<y	��wb��Z2&���BN������b��^��w�D��JP5�wK4��t{�< ��y��w�x��I F�*�B�"yS�i���.O̺DW��E�j������*b^I��G��P5��}���Fsz{�A�y��x{�!j��ڕ�T}Rm�`RS�����ˋ^��^v��a�iKᄲ	3з�صZht��ȥ1�7O&M+t/�p���j&��L�[�����<�7_-�pR7��u��O��X�nkٔ� GP�f�*@ 9.MvS;��W�]㕦HIX�E�Y�ӆ7����V+$��tL32<������i[-lx]�
 �F9H�w�����4_�M�نN�?�84K�i�3�z���cԓ�u6B�1����4!3�,0t�$�%$�ϑ������=��]�m�@6f~b�� �>�"����_���n�d�� �A���l�����Eb]J��"�%j��[�������WƏz�P^q��p����适���H�*|����w�*�ӗU��Ľ�y#��̽_��0�$=:G1J�4>g+��4Hc��e_p�� �W +Y[��)�^@a�݅x��~�F��M���Ul��a�pH
$~��*����
F?W�$&��˵����=�s�[V9܋�wq-78̈́�B(iz����A-Ͽ~U#��=�/lt��l��1�Όn&{�(�O�"EH$j��>��d7�f���*]�{�ϫ�}�m�')d�cH1sp��|�����6 �ƛi�������[{�gO�DQ>u��n_*u׶V���!���폪��c�C#%�j}�_�����5��e��.@�TQl�bmO�Y��$�1�)��W��/��-�0���9x#J�	��U�$ZHX
&�Y,���{=�5� ?=}yof��y]`zq��r�����J� Q�� 
������$�B�N��A���!�m��q1�o`��N��AX���ڋ#����{"��b�^$Fy]t>u�-�qp�"h#�~�������F�"k $�&���e@������X���7��CѴ|���{����v�]!�Z���$�-Ғ\u�̡U��h���N�����#�;�<�~��X�b�_��JLmxĢ�ě_岤[l�k7�������(��!bY./�6��"I�*O��HBK<'G+n�ٯ�u�
����?�ӭr@�P�����m��z(�grUu��T"h�fp�y����o�E��A��n��5"x�KmZ^y���l�G8�������G����4��H/Y���:���L3�.V���Nٟ�K�<9B�	�k��c�Þ������C�۪>�B-Gv5A��^�\Z�cɵ��@})�� ,p���v��]�l�ܶk�L7��T�L��.6���W�B�����"�����b�F%|}OˤB`� �1i���\P�ѥ����C'}�����参 ��5�N���=�$a��L��>6H}��ӝ�����Ÿ����mC�rX����}�.�1�5�÷��Z;�/�;�>U�ݝ![��|r���9��q,Ju�;t�TT_ߙo⇈�?x���8J��)5ĳ�G������4 �E�V�Owo�ni�o��t�����1%��$�"=ieO&�����	������,�*���4�Pn�l�.7l�w*D��/Л�L��N�Vu���_���?7���V�5���hk򁑝�sm1�	��W�DH�����wL���d_��4��D޺�v��C��Dq���T�r����nl����J���y�~�ΒcIb�}l�������ȱ�j�?��[��_��_]0��#��v�F"L��wQR_&kF�@���� �Ba�۵y������
�ݪT�+GV�t<�O`���^��x���M���GPd&F
�
QҶ�\	E-fT����ŀ�Q>A���qPHB��,�M���՝{�,+&S���sB���&
� {[�u0)���;���S�L���x�[����ӻ`�V���?���!yy�	��Z�����[�dXL��yyCjz}}�����Vmk�unu�{:�.�R6L1I��3j�����'�O�-{��oH�;��@�_vT U��4B�!~z���t}4(�^��Fb{7�b����X8X5���OON(t�/F��������O�[#w+so����p�"�	E�>4�C|+7:�Q������'���<t��^��%�E�SdC�������2���v��}��ʅ�Y>�k�o��&n�.3TA�$�P�^��<�䠜����o�o�<�l�Qr�*�7�I��d�U�V�_�v|�xB
R�G`y�߁�T���X\�n�j���E�9a�<� I����7�%�P���5j&�ڍ���<hC��Q��������F�F�����4Q����	6��c��ٛ�񧃟D��x]��d�xWlp9�̎�4Է��f~^�iŝ��;h@h����O�H��,4&���OH���D��p��WQ���-oRۖ���N��,$h�����~�(�T��}�tD���Q)��>VōE�0<��"