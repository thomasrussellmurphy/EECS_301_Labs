��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>�m��`K���Ҙ�ƩV=U���Zݗ0b�����B=��N -5}a�B_���LT[�1����]�r���s�[�WΥ�U�a�Lh>�X�2�I�x��ק������_G�@&�cפ԰�~Ό��ص�ۇ�?i���^���˲_�P����6u&�OA�餳Cd�SG�dڈ���A�?�֍q\t(4̖;>h7�p�7/l>���dN�u�F����`tc'��@��u8r.SC�=�q���\ ��HCxA=���tR �-�4��� �6���x��2�t		X�p��R���L�{x�S4ڐ�F1�M�l0Q��]�ʕ\1|�6�{"�^c͢�r�P��(��>eQ'Ʊ���C,J��%d������J �'�Ee?��<y�JlM�Zbr�[�i7V��Oѡ�j(_�$ ���8�&W��}zl��cj~��"n�DK\{�y16��H�g���mT��+3�*��&r*�wJ��y¥��Vľ��s�{Ѽ�g�O�}���d+�1�uFjK��woɅ�kz�펝�����c�/�U�i!���6��?�/z�����D*N���V���X��W����H����YLH��{��q���K�!ݿ��Q=�WR)��\�I����̑qnVL�2��В�m�1@�!A���)��>&�A>6	�:WG.���X�\����᳁�*��'A9�``��VK=���Հ���}.a����r�fz6F��΋7��#�)I+l�|�[��C�3F��~2��c�jo�T��9�a �h�籂¼�w���'OOZ4l�������!m����k�׬c	��C��L*�8���MG���A�a� c��F&AE�����E���vs�N�0�pɠ��7�����|��{&ۈ����J�m��n��:�}���iq'�Ŏ	��v���P�IeD�����	 �a��f\|�E9%����8��.�k��b�D��P���E-{�an���&X�T��*�~,�l�D8�=��`E�eUv��V�)��fT���α>�U$D,�~R�^�� ��\`��Z �A��`�9X��'Ct�L�T�X����O�]�!6͝2�����Gk��!�\l}T���*�;H�2��h��8
�^J�tl����7H�W��I�;�橩 ��T!�fAf����y/�{�6\)�Wޡ7<��(Eu�%fi�>%H�v[cf�}�\S�J!�b���u$c�a����]G������Zq�2Ǝ�	Fb��Le�(7H���s��D�K�/W�q7�-���S�q�,�b�U��r;L�k>z�������m�����ƚ�N����ȱC%͍���P�^������g(����Vt~8�[(��ֱ��Ⱥ��;ޮ INW��Q�1��'�� �;�kf� ���|�`o��]�����Ǣ�%<��9�n����������nSx+|�/��0X�Z�0O�.��{xY���=0{)Fj��kbDص� t�nN�����:�ɝ��<tm��1 MA�(Kf����\�,��(N`���Q"��ah�� Hv��RB�M$�|au�vǻ#l'
ݵ爈�	�ɦG ��TYr_������������s�?_%�^��R��JO�"/z�����.z����*��_j�v�n�seO!�m`��b�S ���řr4��"7�Sf�2� ����x^�O��Q�l$AJ߫� �4MH
�R���'Fn�
:t����`;�����W���=�o�cL����h�<�?Sq_3�@0��OЉ����ؙ��#���bp���;���Bw������}e����tπ��I��Tag�S�^�{�]D��/�B��Y_�K�]��M�O����h!$,�ȕ��K�����*�Nz���͒�8Mj�o�c�R~1U%�%d�K�+�Ƹ�wt4&?M<��
��笮�%�xw��b ���I&���3G&��t-xLR%E��!���n�`�~5>�A���:.4d�z��U��C�m��&��3#c��MWP!��"+��w���ӶN�l��|�5�{A�"�7��F�t!U��-{-�oJwl�ž��`� ����	�`&ͯ-[���7�f�z
�W��{�L�:R5_���>� μ���T������x8��:��9��_D%��3lS+^v����$��|�w����k��XI]��+���T��?,O�M$K�ݙ�����#j�R��9p:+�Y�����D���G��a�!Y]ף>ݐ�����/(V��a߲��o4���]=�Q�u���bH(���x���6� ̀�X�V�b�����mR^�<Ӕ���u�@@��saUfVG�1��8#�G�-<�٫���X��d~Ծ��xt�R�M�r!�8g�\�>B�I��(�����gKƟ�P�:�9��#��2�Ɏ���?J�^Bn��XD2mN վ�V]�0~��Y���x:����+ ���^>*�!Z�o��-��d�0[�{�\6�t�&B_~�8��BW�D����\ڑ�\�s����Ĥ,�&f�������H�I�jd�U:3�y�>l�3��Y�[�(~�<u&+��ɸ��N�N�q�l������5mh��H'w�$����1n׶D�t��h� L�ڠS���u/Q<��t{��@ޠ���uԙ�
	�w��1��`d~��P�ŭy7g�(�C���x�Ј%�pq\�	��hI�KC�i[w4S];�ww=#ݎ�X`lL�;�{IG���m��p���:���M6w4�����♊�;;����T�ʡ�)n!n+`�,%`u�,
N"�֦�����Lk�j�]��z]v3?���8Qi)12�+7���q���JX�Ae��i��}��}�x��	�3WG�A������+��(@�r��j�j.�:d�/������ɵ^� �SVڮ�#��iШ:����LQv���=QJ:\��x���Z�έ�a��2z�H���R"x�`J��7�*s��U�sb
��Z8���롛�B8� �1y�|V`#�x�&�����ڮ/�{�����QA�_���$��.�K��(�� N����IhaqO�܍ۤ��� ������sDc7�c�ǉ�v���R�H<6+�̡C�<a�r��;L�MlL'�� �3�^W���+:]=��0?�	�RJʏ�5�꿿u-HRfOt�����I���](�u��>��f��*fi����u���Y��B����X>�*�<�B���'�zc�C��]��#g���jY�S�ϟu�!�4c;��O�(i�*�0����P?I�f�
�4��Hv�Z���/P2"��1�nQc#�8w)�1+]�K��#�����(?2uq�ۑ���6ί�#�sy�ߴ�>