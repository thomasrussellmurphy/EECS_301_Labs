��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�i��a
Α1S%� �uj?�L�3��TLei-3^5]E�$����u�E�x����[����u�T�"^8�WB�)Q���q��
�N��bۧC��l$�7���r��9%���AO\�Rc�Z�n��5:F�nۖ�ƃ�>�T�	���1�������I������bX^n�=���Ё�dU_��r�6��M;6,4G!�ğ��V���iV���e�I��n���-�հճ����x����S&�q�v��J�����g���(��0�k��q:�T%�5��/zض��C�8��^�lZ���?dˠ���-�gڦJGb��$���4���ơ��M.Q�H�u$Tl�|� ʕu��Ө(�hP�VWD��67C%��{D�Jiy�ݼ��g��x3LJ���+�R�G$���?hbo��y~��(7��\Jt=/��s�h~6iZ�e؏���M��b�f�����|�]�2�����1G������iQ1�D��1U��ǫ����h�T�v*ns�/0�@�F��ZBG��6���	�W:�n?�{Ŗ��Hd��x0�� �j!���p�,��(x�w*�O� >�,-Ugq4&5k!����Y&��U.8�5s����+ �.�瘛,���Yn(7&� �4_�w�}�h����sH��� D<

7���$Sz���֞�����*9��|�؜�g�q��4���5A�)x5b(�D�^;�.���%k >M�2��#�����!�Q
���ji���h�Y��uCp���muW��|o
9^��y���y�Xq�<E��\�*ssX�������w�x��F�)���g���4���9}�7N10��]R��h#�w@YV*ʬZ�:D�jB��z!Io�LN���#�sC�� ��"~k��jW��IM�ȗ����;T1H^O>�6��nfN�շ���yP�&�&o�Ik4i���w�7�\X\R���k��<���ĕhv�f.�2O�L��b����`���Fj.�9��=P�`�o� �N7%�&Dq��sqzps�Ft|a>����8gG�}�C�';��b���g�w�e�]M���;��
�}%<�N���z=D�M����F�oM�LfTA��_���W@�'ci�i%xE���� D� ���[�HML��_(M� 2��������i䃾�h�}������?*^��2A:7�mȈ[b��Ŭ�h�}_:��=�lsS�n7�%���]����f٬[�鬚QY���Ɯ}�-ڈ�P	�z�M�}��;=>,���A�BiQ]��?�����y��C�z�]WA�.�!��ˎ�����`O�2��t7���@'�ۉB��O�6LD��"��B��dkl&퀧��?E<py�#�C��3�Y��fb�7�ڤ\�ג��P�%�ٙ�~e965���j����(dN#c%�d��9���T*�6��:��* �5"l�ޯpd�o/����cp����"�$Ơ��4�+_l@���X�1���`öO�O�<�ǩ��ر*���s2d�SZ�*}m���u@�T�j�凯	���t�f��\3��f���佸����'��H*�+�Ƚ  ala�K�N諉��&���=fj�	*�0��Y&#t�zQ�݅��(R���"n$�B��:��µD~b:��ۅ�iv��B��Z�C�B:�����>�����v�VvY�%���D���͑��rI��<��:���L�Q�F��D&�������0�.B�s56�z�|��=��I�+X����X%Y'�b�DIZ�d�OW��f���H�L�=l�/����Z���Ƕ��a�G&˽4:�-c,˄�]���n����6^��Q��[�"��Ġ�yr��M����(�zj]�b�X���@���/+�%NXz�Ƴ[�Q�ʂ:ٲ���6���:kG�ǝ�E�! ��8&���7�U��ͪ}�:KQd[�z[�ÜpG/��_���t�d�#�$$�����>������I��\!�4�;���_[&6��;�b$1
�$���]���a��n\�q���Lf����� �F��+�Ӹ�PU�Aӈ�<��M%��p����c'.�����W�$�:8��t��Iv	����kQ���k=��zP�(��h��g��\�����i�h��藬��O�#]���Q�c��V���?4&��I�2�K����� �F�"���2�ߗ�,��V}ؑk0�w1���2Sf�[>�*�.�)dGVg4�r2��BN0�^�|7�"���,	��9.JkK��9�A�����z';���v����;:���LqU0b�L�"�˾��CZ��T�gvJ�&��B��q\��Jzy0�Y���(�!)���x���ԯ|-�ĺ�����"�S̍��-Z��F���E:�)��� ���ر��ta`9�,)��iB�QN���HmL���p�ʲT�5�
�|@��Zٱ�d;�pW8{U#�O�h�􂆂�x��P��pc<�� ���\�	���łV� �9����=��v�18�Q�6R
���b)���)̮� q ��&���ֱ�jFbTFP��y�#���k>=�H���b�J+�1�%���tfJ��8#=ė��T5`�xj���|�rI�}kEUkV�.��?�Gsbg�.�����=��������X6Q�̢T���'�`K���P�P孥�_\`����n��C �[��+����LS�j�����
18ԎHc�42��l�P%}� !c|hף������@�9��^x;���f�7A�W�;�?>�Q���;�܁�A��4�Ϗ�-��U�/� �\���J�xy�c�h�s�Z�F
�*USb�N��ۃ�\���G���p�	����Rz�����c��x�_ >�z��Rf�u�AV�`%Fk�
��"$�w���e�U1��X<��cR+`����-�>�lx'����P�!S5�{��=�l;l�+�"�C|������.�E�N.e�8Zy�lQ0T��IhlJ�>�(�a��Y�?�_�9a%{��