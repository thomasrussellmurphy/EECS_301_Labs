��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��We������Bu�k4�)̋���3�2�@�vz&B}�x���0.wExd� e���疨<�(	W4��O>�i��ɒ�b���7�	��ѣ߳��EU0"�vR�I)0���U�ëA�u�������>��E�hKۏ�Nӷb���~�y�"��)DHR����_'җx[9x
!�;����MX'9Wb��w�P�"⽥%��j�F�r���c��.����/?Q0�Ҹ&
�� ��B7y�HY�j��p�0ϩe	���l��P��~" -_����<Ӓ�������$S=*��_�� DB�Ll�gK�y��i��~ei�)攝J׳��S���%����4P��IFM��lU������S�B"g��c���7J�j;P�`\O�X�1L��){_Ir�ń
�����:��i~�0L1��7z,0�&���1��DJ�J;���=1ų���{��u���'b��[�,c	�
lw9�@�$�kl,�f�['A_KSC�|A7w�Xܽcp&���#;��0�+���~��.'������~aD��QY����11�;@�J���8wk~Pr~�׀לh��g�=x2������N� 9q�e�PZVT�O�mP	�]/��]����������|&8�~��=u��a[q���<`�V�6C)�[�<�;�f#�h)�W���7-l�P�N�@��1WF����'0V'�Kj�>��٨�3{�J���v����`��4Q&��.��7� F��<FےU��^�ߙ���*F�g��w�㜥[ u���ˮ�B�
�q)^��W�G�h͗qKۂ�\�$	L�3�%_���d�&̓q�8J6I_��w$�ķ�Q�l��Y�g����Y�):��ި.x�|ߌ.��A��rBYr?
�z8A��򯁇�'�L>�F��@4s/|t�X�ny�x�3m�@��n]�MBp�UT�^��5�R1��8�*
N�4��ED*��6iX�E?|<Rg�Ÿ��s9��@�Ѩ���l��N#Uk�W�6���%�����|C���� �cV��jg���Sb�/��_���~������h���̞�G���l���U����s��@��� �}}�O��0l��� b��b�EX?�'W\���]����n�������F�#9wtY�x�`r�%�҃?�҂l̒Lp��۴����G�6���o,i�v��-c����~�3Q��i��}�`,A� #C����6����������S��{�ǩ�E��8t��'�c?�tl#�]�TQ׿�1�>˯��eyX3�9-'Fc�&�f�����/1�՟/��-g^�bU�
�Mz�0����'\l �����Әb�d��-밊�Q3��ޞO��^b��Geunj2����ln��I�e���W��"�)n� :�i���S1��u��cwM��!&�3ʍi��T�QU��D�OY��	:m{�w7,Z�	)�a�Y����6��qne�LD?!�(�~����֫"F�;�7��(�Y��]�7��b���i���1#=Xw�_����� Q���_�����!*��{�<'{/�����i�xق_d[��VA�\����"��5�M�F��lz����`BL�mJ��_]�'>-;FM�K/e�7�HS�;ZS��)^�S-���Z�����f�E?��d��y��6�s��S����uMv(�8�B,��LE���`� E�oJ��Ν �	WZ�^��8�={�� ^����2n�_"��| 2�z�e�flM -�(L؛���vj���.�H��0u�e6(�6zKH������a;��/��FLA&��S�Qy�kn~�D
E�;M��;C6F#P�ᄛ�� a;���<>����k��1��O��v�/ͮ(��� ��O=��ňI���I�䌩x�u��"�H2��צ"@�*F�z6���������n�c�k�ۇF	U�cC(�S=MEJZ���FG2�T��<�1��Z6�x[�v[�N���!���Ry�q�����D��rk�"´�͑�q�*����0����X�wT��A+�m�8�"	���,�+�hc���&p�@8=ƣ{�`
���"m�o4ٕ ��6��kB�?	#6�|���ןH7��S���Qҝl�eEzl$���RP����kQ�b��|=a&
�ԛƸ��I�٧�v��f����ăp���v���۲��.�5�ލ�19���7�_�F�^��15֩�*��c�l�)�s,���!����� ���/�m)�(��\Y��P�
����}uoI��S7g���W<���B	�H�[/�*+�e��]�����Au���e9��|��F�����h>���ך���`��<�^���4*Dv�=e冑���x �	��M��5���5�'��%"u��db��=�"/Z�ý�;���d>�YE�dA1���-����N���8O�)D%>ѐ�Y��i��v�=�t�Ch�g�f�����'3螼(�& �?�Q4uE����?~�zo%*vm��5��qB�tD����1.
;��8w�h��ѳ���ǚJ�l����� V�f�6��hW�B�j:}M��Y�I֭�K�M����yE�D���O�:�戦�c���ԷS�u����0��M��E�ӛ�]m�S�t�f �S��܇��2_��HO$�	��k�Dԕ�T������)@?�.��g����Ej�-�����x��YJo�1Ш)�I�Q�^�6�ߜ:���9����IE�%KS>�уl��P�= �A����{��pr�ϑ�`�V+}�Ӗub�B� ����@.������ܘ�L#��O[��H��^Hf��Cr	�\og
�c��LSXg���!�����@R`>�و�/��h��]�wZg�T�Y����h\�o�_
,~�y@&,ʏؙ���` ���H�������-���6|-�����S����F�tì�G�z����[��5T�`tUƝ������(�:�ɐ��g�0�#�"]J��ǽ����f*�j��ւ�M��m[FV�L��;�/h5���a���j5��l^��n�;�C�ZT�"� Kg:Ly-+*}�<8����QԮ��=����B��)s]�VH��D!�7�y�d��P���ɳ�����"P]�&�bdY���<�ҭ´�kc�m����3��H��h�P���ɉ����+p司�R岌7Ǫ�*0�]� �8���G��t^&,x ��H#	��a=�,H��L��1�<�ؗ�\
�F��`�2H������n�m��b�Z����h�������y���2Co�i1a|�7^��z�� b���lcr%�>7p��3/���� ��%�=�O?*`�xTr �ڿ�C_��R�R�ş�b�^��g�3�ރN_37�pJ��{�-����|aP�Oo������2P/�~���1p�ыT��4N�JTQPXy���'h<cmR�{2�1`�.�"<K��'z^�.��P�r�����;�4���L>"l�sN/h&� '&���&����_���ma ū���&n�ܟ��{�NǱ, "5S<�R�x�q�K�" 	4о���D�e�t��_�C�&�\hs���4|�`�1j俘����B�t��8�����B���2�I')4:t����ۿ"8�Eh%���
�4ح��Y���G��L��:o�������?F�k���D�yl �N�J�	�§����FT�� -�F���b9����R���W��
�K0$^+�I7=��R�	��h�4��jpr��(P��,??NM��~C�� ��\�B��[�1������*nk�ͷ�0Py�@<b"MZ���R��N_�}�4V0�sA�Ӕ��9�Wh�3��8��~�U�f�L������<:��ō�#H�*��c{�":j_n[�sy�Z;+��x��@�I�l�_\gz�PBjMos%����R�X�>��ZbMj�@J�l!^�Y(�T��v���ASܽ��6)��S�6�3��l�����!��	U����	�( ��h��������(�KU�%4F�~�q��t�moG����o]? jkZ֎�DS�^>U���QM}Di1
@����T���D�����$k�IԢܞ,hGM��3�.� �׋��	�ޓy2�K�h�|Jxw��Lu��- D���4�9���Y�#�|�Ey�#��zn�+k���?����؃�7����(��;a/,h��e3�^\�"L7m7�1�i������J/c/=�U��W�g��ǎ�x��4ٲJ�w��b�a2Ht���d�$��9��MH�e�N�*"�Gے/�b��?YL�&��?L���X��,"|��Ie ���.h��t6�:���d5�4����z���<K��=�}>A$������a�h��o��B�E΀�5ѽ�#�#�ZP��7!��]J�o�u-�~�>S�o�Lq�!R��a���'�:�L!��AD���-׉�W/򢆹���g�9�����Lu�����D}�5`Ŗ�6P���Kǯ�`#+�s/q���})p�@Y�8e���>��|��T&�H�Zq1�W����k!����%c?`�a�-���.�,߁�hG/�������E颪�����4ާϕ����y#�w=�nU�	���l�>���z�}	�x��������3Ν�6V�ؓ�������r��E�V�yÒ�T�+
V&M79�C���n�����H��	m�F�sY,N�i�U�9�@�ig�1��;�t��pﰆe���gׇ���>�~��DX�5wqF{�H��r��?����Sb�s!�݁m�F"T~D�Үc�S3%��C/I�ӳ�g�EU)y�+������2�l��s@��6�	c�1����N��79tE����t/�IQČma�S��cR�F6_z�bه���N��N�����>��o���N���xѶ�}��&��-J&����85�����Y]F6���@�>5��ij܃a�:B֌Gxy���M�j��(^0qkN�̔h_�;]�J��:���&Qy���O��J�f�������j��K*r�8�:F����7+Y���&�z'h(NH��g�I��*6�X:�2y�*U
����@��-��%/�`/������|��k��k�t�No�%�&*���1b<<�ӥ��Ui�M���BZz���pH�67NIj����I�~�3�"_� ����э2�L����ll Č�n�Y.�`�3�'��Z��ও��`S*"u�QdS���]t����^|�k�J���2j�s7cM�Ky=�%(\��_ �F�@������x��H�_h�DDKH[j�Y��P�e�K���]@�_�x��r!v��x��]v6��='8i�R�q����2p���F�֍�DS+56���.!})Q��_4�R+f�Xixh	���v|�0 ���|,B�jrGlw%��$�fBaG�y�U�1���Y�E��	�u�~pN�g��F|ʊ�T|�ב��\�:�P@��^|�f%lU�#-�N^�c�m�)���WL�
8IC���Vu��ha�3���b
�t���?�I�l�^k�x\3Y��]Q� 4���5�e�~��r��H��1X�iT��	���@�/Y�1���&�^ab�F� ,�M��2k�0�4���?�-u���Y�{%"��=�9��I��	O��%H#�M����O8-U�2ޔ��Yѹs��N>�U�����7�(r�ʝ��ȼE2D��s*�3Z�6���;1
�pƓ$jȌ����*ތ��I_��#J��Q�� �*��о��i�n��s]��u�E�>�0jl���`�l{:FSud��T8���<����_@�����.I�j���=����]T�`��Y{T;�{��龕�MQx�:�=`�Gn�$#S��s0 U5�E��})XQC*��)�����4��u)fR��,D�9+��3���tM�#j�BcP��LI�Q�|RuT���$TnZ�u�?�)�,��4w�h7���b5�l��)_k�ne��t�&PN\M;�����ߒ�ց�v%~��Z��(I��^� 9wй�����z,5  �C�4��.3�8�ۓ�;�	8ˎ%�\)F���&��.PD��9�ڱ�Y&Z�������F�����Q�t����e|us�4<��"���58�z���Ɛ�o8��h��[WV���}��i��0��-׈��slH]a�a[�$� ��Y`qϤd�*`�x���T˘������?#T0F�R��=���,:š�(v�>���LR�-,�b��N����K�2m�VYƴ�x�O���k����'��h	26���z)����B�lܧ�	Ͻd�?���]Y3W`�ɋ�z#�2[��f���\�U�(B*��n~�	�<��-�4��f"�+"��,ЯJ��M�[F��vy�2�A40�����/�F���Y��Yy<���f�`)��̃����-����?Rw;Gdƃ�m�9㠊4y#R2��E��4!$�i�7�7'U�ec|�e `�u��y�2aT¥�9ÈF����|������~�V1�8���SʉO�?pґ/���'/�`X��xڰ�KG�\�[�ƚs;���&�.m���0�ž>��E@o%\�������mEm�K��bV�����sH��O��(r'�@�Zb���-&�eesn{e�#�Y�S�lE@�8#%N4��y�ͼ��<;��z1�D�ߝ��,��!tN��y������uY֫��(��	�	C�3�����L��.� �kn*:r�r�����
��_i��������-(�E���D�BZT�},�JVۚvH�}Xd(�v�RsYF��, �:�=��"�1>��o�Z�_;���X�/&��=�t�����\Y�
�3�NV�d��C6r��r⾤��|���"�芡�paA��\��uwY�6�"���!���̸��T]<���Ф$�q��ű�HQ�<��a��=�|J���g���p��`	h��|b�6���%�cpL�AQ���`�s`cH*&vы-p�m%$�3dU�B�wי;e��
&��Z�d>��2��7�΀��M�]�����OOhM���G�"�')b���!��lE+e&�2�\�g�L��PI��~�md<ÿ9j�u4t *
2*��*�<ǭ�[�P����8��%z%�=��D^�%7���F��qx1����!�;��ɥ���`�ۺ��κ&nP�2�Ă�m�F���u�P���,�9(�(�5��^�����[����h�s7¿��\@?��C���
�{;�Y{��T��ф_l�T�[��%�ҢF�N�t�QR$���{�9Y%w�+lr:��@�Q����
Х�����{�٠��c��Y�=�%4�b�N=Ix���,y�{��A�gt*�M�\AF�z������<�X�8����[b35�<�V�;�c�kT8�Z� �R܁}���T�� ����� �^]�XN�*�Ǥ\���Yx�� ;�,[�N���-kdz� �t����Fi'7������%l�^
�'���G�hAO�4Ǔ܋Y���$�89��(�Ϥ�A'�eYd�y��B�|�Q�w���g��N���g��*��Mª8p~j-�����T�����fm5e�U5��:�7�`d��;��W�[�C=Pt.����"�DWW��)4��e�v�=�-���T��v��^ғ�U��Gѹ��1����s�!�E��;�\[�`�'��C�̙٘AzF��8d!6��&��.O6+gj�ʤ��;p���e<SV��`z ģ"��8���~�軰�fJznNҍ������S�#О�������V+�WU?�������Kܳ��cot���_�X4�$H��������`-I�;�F�Έ��7��=�s�
�E�q#���}IĬ�e�P�"���%w��)):�O	L���&���q��#�U��v�p��f]�O1c��Q������LeL���3B��P{O<�s��y=\��|����0�o��]��@3��q�n��9�8����l��X^���,Ete"�����6�}
0o��� ����ISM�� b�A�p8�	=oa�IƖ��X��=�l�?�Υ�U+�h����J{��~���,!�eQ�dv�F�i�Lj7���p!Z�e"�P�����{�`�@���4Qk��읐�%�{U�+����)���P��pp�Ϩ1bp�eMLD�dBT]� �Bv��;m�W�x��YB2
�9S���W��)f�AL4\��槰2U*���K�QF�1|ۧ��O�w�oѓ<�+�w�ߎe��D����9�~�T��p���*�+�*�"oR���1[���">� ��ws��J��~��7�X���@�Z$�6�e ~�Sx���ס���� ׈ Q�5�}� ��hX�w@a{�}���!t�#�~f�$����%ԓ\"�E0��fq#�#>Ġ�m���"��|D�v]��C�W��F�H��L{\Z�_D��=�[�Y	��Ygӽ���8���Җ�*Z)X �Ŗa+ B��)G����wiyT�w`���V���-��i��0�AƯ��He���Mkm�~\%z��_BE�#�y2ka�86spf#�4V�ɉŖ=Ǒ�u-\�_Р �9\.K]����o*)��i�S�$zSRz{d�b9�f�D8O��R�\�N�4�O33(�S͇��ڞ��u�Y��q�?�� �f�dn�/E�NQD�Y}f�W�����m�2�,+&[�#'��i�b�T���߫�N�1da
�k"E_��<�؂.�P����jr[-'2ZK���e�i��`�����=�ݕR�����X���8ywg0����	���$쯽8�U'����x�xk�~�c[N��.[�ȧ�e,̾���n%�li�	�~����)tt�� ��
Û���6'D�(�9fm8�=�y��s�:A2�/M�º�|�Y����@VDSr䶶I�r�c|�ڲ��^�P�R�oe5Pw-��Z
�y!Y?2��4۳|^��6'溞,�Yr����Ha����d�?#R���RGe��G�'{!���"\s�I�D�L�<i�D��]�M�2�<���	M�,�랷�=q}CD�Ff'>���Z'���߈M_���
Kp�����vkީQ����|�[ىw�P��J��-�^l�op�daqH[%�q�Gcm3�:�i޳�ڻ��?[NK3@rh��&%e�sH��C=jEA=`)�ut	D䉿���S5���̧6>���j;z9�V�CI�E�<e�
��Eg�޾%�B8&�_]����cP3�k�|�� ǋW{w!7��l�bIǒ���P�����58��\dھ�Y&�΢۷�CH�kz�- �®��\���U���&��к&�&dO�CYr�Szl.��5f�@���h-�O�#���X��/5����?�6��2�s\�Yc�����jd����@5�p��x��d8@�nuG�]qF]s3��֤3���+2E�{K�v�,g���f���;.�v�+�Y�1�Fs�s�y��͌	��/z,[Ŧ�j�g���� u`j����̓ۆ�@aQDidk�k�^d�PGT��S�\&W�����9��[�5��&�Z�R�y�����S3�������qÈE�ӂ��=���Azh����'�֡^ �[��W����}'JM,�����2�#�a�-������L��gw�ܠŤY�������Tↅ��6j���#�b��Ύp����\�7P~k!y�'��_�O�t8��ݗ5���t�eD	����8�X_�F0`�Ri�]v?P�_[�+�)G��6>��}��%�)��>��!�?N��V?̤X���klV��$���^=�
�i�Naa��i�O��@4����<f�.38�F�*�����$��3?��T� �؎�"��*(�w���r�6d�R�ʔ��WA�w��5ķ�[�fN���2�q!��&�aa�"�2s/�*�FD�C)���
&��8���$�}�T@N�՞�(,8��1S��%�eQT2�r�`b�|�A� <Q��Ǻ�R�Nv���Pj��L���Vro
!�q��uԭ�XR��Ҕ T���ʩYM�G!�ɿ����t�,�ۀ�^�V6���8#a��j.�LΥ�[�V��t`V8���5�V�L*y1��ż'F���m����-����P�DCV����qUL���r~�\xv�R��	�$YUK'@�������-�`:� �-��@��w%7yqs�%��;��Pl�m井e���O�(�Ԑ'	WѰ�����~�������ȱ' "o�V�����|�X��l8��j���z�+a�X4���z�Z��6p����N��TƝ��X+b:����]�/"�4F�8j/� 1w�T����`�Ro��A�B�̕O���V�(�3)�5�2]�7v�05�qD&d�z�o%�������g˰����ȒviԳ���h��8� �J
m��"��5����B�C/Ք�1��W=���
c%��z��F���e_��������쮒~��^���*a�֝k�b����/��d[ݨA�O�� "��U�'[����qv�㐷F@��NM��u�vb���K��\�QaX���#~���{~���܆'��Y�(U��3�V��Q��g:�w'0��Q�1,~��py��t�O�)�e6�^�( ���!�T�c���\j���R7����Z�����t}Փ� ��94�L2%�U���H��2w��!H ,G�@�T񥏽6xR�%<����Y�9*�6<��a/,)�Ҫs�(W�,#�!`5�EӽEe����@��_�w����K�H*���k�));�q�����8��%"4�.QЩ������^S�ҢسԳ�H3Z�v~_$oN�œ�8z�.#q*{N
L�S�{m����Ɇ ��pHR�U�J�3M"�ͮ7��k��b��mB��&a��1(U#�]�W �^�2