��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�i��a
Α1S%� �uj?�L�3��TLei-3^5]E�$�Ԃ�󨀊�l4�JM��\?,���=���}$��?5��^�BUE��jZ�*A#+���0nZ�:I��7���5s��!���:Z�~yW;t4�w���h�4��6Q�9�Յ˵E��?k����٣��)G��EG��Z��*f�1Jd0f�����P�tr]�_A�IE���`s{AZ�0�T�1���Cs����%C����3#c��#�8�7�w�k�dNY��zF�jPE���6Mj�S�{��[	{�Ka��,��,�m�R�$�c������T.��~.s:�ƟR����%Ho+u4�G���������1wKЊ�e~<�ҭ�L�Cq��KY�2�7/�A�t��Ϩ��i�B�5+��"z���N�z�����C�u��0�~w��{�rp���\A��8��t�$�$KJk�|k���k��ϦϽ���;/��̰,eX�iz}����> �$��x��ɭ�妵����ϒL��gd�"v8Oe���(72Hn�O���8��N�����iO`�w�w�%�ǚ�-᷺d����t� H�H�t��	υG��H�������JӁ�M!���qLŪA�������o��?�S�/�� �ٴ��7�n<���y5U ���5��6��{�4��a}~I �S:Ʃ�=|��箹���~��!$4�VL��� ��}VAԘ*#iDb�U�b�:�0O�n����/ZO�`�0�p<��0&��AR��Oo��ț#�sB|����ZI�w�>c��@�Ҽ-�/��c��<�����X�#� �-#^�ԯ��<��#�[e�7�3�+�����)�*�f�h��Hk�7���UG.���n��n;���|bRaZ��5����({'�7������Fd�@,"=_G�4�;���AB�;L5raphf�S�[g�ӆ�����u���]|�Pq۾��)��>��"��%5���|�O���q�1V�Q�3n�s��(+���Ge���D���3��qD.<�I���0��q���8m'�D�,!���_6�hPCm}%/=c���r�j~�k-�x����H�t3��\֌wM�װ��|�#M�ݺ�?�á/�q�<Cl�~�p�?�H�	Q�6��	^��u��
�����o�f���*�KK�����DLO$�����g0 ݯ��`��H�Q]���Nn'%��ݖ��i�ʂ�����ș�~�c[nѴ&B@�]:�uU�!q ��i�)M�� ��� L�̰P:KCI&��*��;>����0i3,��e�Z~�L��P��Nx��L���CZ�UyJ�[@l�F���![t�b�Vֺ
�Y=�&As�����Lz1��T��dx�����l~�����L��A����Z��8+�Ґ	�9�t��:Q�*~] ����*+�aެ�.�^{؈P*�h(�n�C��!���Q�E&UAN��g#Ľ�扢�<^��e~v�b��G&�a��K�q
A%G�7Mۺ���Zt���6AN�)m��ś�����v<lcn��3��yyJOK%}S�ֳ��oB�]=[�Rd6��G'HgPvs��`f��w-�N��a�a>{��k�壏������J�'U.r~�A]�<�����y�H΋�>N�����+�d�+=�Ͻ}ԋLx�����Ї1V�B��z��&�*��B��!'G�U F�x� 0�>ph�Kd�B��M�(s�7_�����jn��^$���M�N~�0���c��C��[�e���r �T	Ux?�U�*./�J�(n[���U1�s�
b0�TO�*7�N~�(s�P@�Q����1W"t �,�G45���stq\����Q����)G��E������kڅ�5�S�ز�V�4�UB�����#���.];Qu��ń�Rv�-E~�D�e� /�~�DrĚ�}��t���_���.����'��B�&�cV�\qٕ�B����w�`B1�5u�,e���кF�P�yV�| ������
y9��ҩU��w�zj��X��x�g��<��Vju�Q��ta7oY�2�8a�(�n�I4k���]���#�_�����^� f�"�ˠu®��y�E�Xh#vI��`_���ڀqt�DYF��Ӽ�:�_�)0����p�F�������m3�#4�ȥI�ά1�ݘx�'K��}̓W>o�#5��[��,�RK�is��&��y(j`���<�2�IG2���Bt��R�|Kd��=���n�[�����/�}�	��a�.�I�+%�`�p1L�%*��Eo��^9�Mz&}u���G��\��
��j
`���*җ����= 7�c�d�����̮1�3̥�䃰����f��X��@���0����A矞����9�ۜ^:��h'�.�{[�0r�h�YD(I�_ �;aզ�C�0=�@@�[F?�i�����,� ;�P�?A�O�'�_4Uݥt�kfs�~AwP�|D�/f�*�{H���+و��o��Vd%���'4h�������
�+4k,
N�g��U�oX��qf��'���59U��";@0)U�3\�^X�?��{�ۙE@bY��^E��Y:v�{Y��_`a���F�E�$���j�7�bK��2զ�C�Y��%Y�
,�� �i�
���Q�oiHG��O���@�j[�r��eێ`�D%%��A�¨���j �l�����DN,< ���X�W�T�I2����
� v�c��X�� ϙ��mm�N�YB�g~=�d��*�L����ig�a{<�1]�+�+��|V�]�ޚϽ83rϙW�Xp7��  ��ǔ���>�D�H�>g���@�1��I5�}��h�U�tIpZ8�8�PC՚�
n�NH�۪�K=�ny�x�֘kӪ�p��yWi�d[�(����T���!�P��nppT)���������nDݭ*��L��*x]�E/����Q_��}n-W���ԧ���˅��\@AZsU�
�K�UF�ȯ�) &�3v9	-Eg60+P�}[� 9���E�s�_��rS&J����H�T��+P;��G���H���V�x�Y�I8���}FW=CsӦ)؃u���!/d��ra���o�d#�9�!2��*�#|���}���^N�?�4��/
��P_�M�[L}o3���]�����R�\-7�I& w�OfU�9�7��*LRٶbR��$-��[3�%\�I��6��>�O��@�PJ��a�c�j���|f�G�NA`�UpI՗́�'~��&�X�s����?����à0�u ��ky�Ji���c��n����!tX����ݧ����"ߋ���:����Yy(�Ĵ�4�����$ݹˮyV�0����z��`z$7��	]�:�l*��\�x$[ �kMF�At���^������� �?��x=�OL�g���q���(���q�4&7��1���X�UN4����H�"IӍ�\a�����²Cl�OG�����R�#.&�2��#~.H��J�#?̌&�Y�;6��E��1Mħl�v	���Ct���<F K�M�x	Fg�j.
|��6�!�ƿ��i�R�q��L ۅ7�^w[kT�?}\�&1]t�䵫.4�@]������=?eUt�1O����]���D���`M�GU�6�h�lQ��oI
q���o���&��o�}H@���#���׊jg�r��m��A2�����Q�
j�CM�@����T�4.^�iZ��6�Mɷ���y|)f��e��l\��Yy"ߨq"�έ]���+Z��+s�|w�E=� �0��~�_[�˞9�����Ab>�@����y���j�Y�e9�Ԛ�$�N�@��gǖ���Ҡ1���9��l�_p��;���ԒrR|A�j�[�� ~o^!�p0���ǖ6�9^���ty&17׎&Ό�b^��F��	���آ�N���u&����<�K�<��y�����w��Cm����p��N�<��[HN	�o���װ$�P�)������ة���A�����h�81&�q@�xO�d�*��� C"��l0��U�w�/�m���I���	�TJ�f6�kw�m)�覚&�T��Xb�O1IY�)}-?�6�l`(R�����젚2��}	��ѭc�D
4�sꁝn��!FcbÂ~V��s�7�mA���W�D*���=Z�L�Px3٬��A�q��$ޙ���|v�~�,M��:��� ���L�3�ٵ"�̨����G��*�M���\m�-�:h�)�Թ��v�����5�ZG>$���3<��\~�1O6bq���Z�ma�9$D�m��9	��S�ga������Pm�0��}�S�IAQ���d/��v���U
�l��,�m-���O�ֱ;��'�7�U>9v�{��U��x�Z�F��T�)��I�'T���|?�q��H�u�5B����0L�~���C�'�G��L������^s���aA�3��ȊvK,��7ࠋ���	ې�SE"��1�ȃ��!�I����Xk�O�xL��a���Cz8���|�"#G�+�t`����J_$�� :���Qƽ�l �M?�l�}��ܧ��0m+$�5!�6��Da�.�K
޸_��J�/m:ML�x���wg0����la�*q'��B�3��X���0�x�ܮ�z|���o��,gQ�jpz�#l��Z���h'[>o�)$����t���=��*L��U��g��ccV����5n�qd������C��S:�ŝ�~�Z�:�O�Z��'�����6����px��%;�v���v��� I~OJ��� �^6k��iaX|���aG�kt��w����Gp�.�֔5�g7���n	np������֟(.�,"`V'��W��D�})94}(^r�ZdU�H��Z���]�q�d�����:q����Ffn��4�/ڼ�a�Z%���cd�G����j�	���a�0��o��'Ã�T���Ѣ�8� D?R�P��ZU�)<t���
<���;)SC��}����
f`p����P��c�;Q
��	E�$̾���	�hPï���o�m}�*C����c:cd(��\��%X�#�e��C��0�&��w0)���c�����	; c\�ݻ~��4����`�{X �"��c�����
-��<��q�Oz@U��bg� ��ٔ�Y��&o��} �+L�R�/�^��fH���|e|"q�3D�.9� �-�Q�����̸��ye�g�Z�v ����1Ʒ����l��=>�u}6������1Tf�g ��y��~�7�p�T�
n�h7c�����^R���(c���ϛ�,�&*�z:Ā�n��D�b<=�Br�����B�#[�a���٧$�A7 �)�a�����_T��h�j�v��8j��o0�d-�co�Õ:�#fF����dY=�
i��5{�6Nk�� n��C;�|ɿn.��5�98�V����턞F��tF6�w�i�y��3�N��<��u\R2�4�X�u���l����
��y	�Oy��)y�=
� ��4�]�o!}8���� ̯����r�3��zҺ8�x�a���:�C 4=��w�M0�i
0Zn�5쒤P��ut���bG�Y.����7ܱo�h�gc\�h� (S{0�ҵ�]*���cA9V����i]YZ��R������\���b�o��t���h����%�<<s'�'7��3��J�����Ƌ{�F�����N#D3�f��;7\s��Zd��x�ef��O��Ҹ��'��a}y]*a��eTdj8�9�a��\�W�#��qؗ�~��]*g���$�#^����m7&��n"#R�m+��h�6�//J���#�B��2h��^�U����lP2����`v1�yp8uU;>.i'_��>�rʲ�ŝ��%���I�Dc�W�` *�jc.�3SfD'�����_��n�3��VZ��x��7�&&�<q����g�j�̕�Ǳ� T��ۃ����?n}��v������S=e:��)����̚�ZJ3�g�)�E) ��Z�\qZ���#�_*|� ULTe��<X�QiV*���
��B��5��G.�R`�#L�^��׵�|M��ةk�N�<�Z�ΰ��@>�|�H\.��0��koZ�ls�>�5��&�