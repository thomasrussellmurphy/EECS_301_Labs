��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\���V�fnvx��ÍG_;�ȅe�~�>���9�>��Y;�0G�J	m�_�0�y,�T�����_�-�V�~���ƊT�g��/�%�:j�7�����o!�	W�g���(�m��e�H��jǐ#�Z�b�c��K��~ͣJ��������~-
��}D�t�ߝZyl��?��1��F�ob���}#"����$�;�� �;�?W�գ�������Y#�͍��u�m�Y��ܶ�Z�-��x�-_�x+�@�G
{8��O*���dz:�f�%D�����њ�B�Y��G���d�՟�J�:�eY�|6{���j�9IԿ��1Q=�p��݇����� P?j��0X�w��"
%L߷���
�.P��1!${�kP���6d.�/KC]K��!V�*:�:�)
�����<j��`>��Q_dfS��#)XP�Lc	��_ك��*��T�����-��j� ����!\N����d-��7��Ĭ��J�u��|q��T�(�'u���txT�zP�N�U����塵��x�.���t����Q$�_�EH�D��Sa���`�;�&��hף:�s!gF�y\�g�X���I�4�48�1<A�n^��_��+���S�vX43MP�Ȅk�R]J����еکj�hkD��e�?����N�LM=g�[���Od٧�+�lT�2G��~�^����+�) � �}��CC�_?v����{K�I�hShs��I�Ӳɸ�e+V3�yw�\�Uo�P����}IaIU�ۦ0W�a�����-��r{�Ƨm���	�K2-$~��>my ���h9�=tM��n!a\��G�-"H��a��"mP@C�`�(q��KgG�u��&t�D9T�;*_8=z!� 4%@4_��b8�J`:L�g]�=�$M�.��v�Гn�y��'��+�>%r۲�O����W�����ѽ��U�bX���ٖ))TӋ}%��ǚ��Kȶ5����F!X�U�IxP�R�;���Q�fi��
-O {e/�Nc� �9K 2:EL��v�l�Ms���BWA)8��ҌO�F��W�k�;M�"�����O�s�|f�G5���*���p[?Ҩ�,j��2.[�՝���U�ZiK���R�U��h��A��q\���r 9&g�-+dm��,!�/L�C5��w3���6ػ��2�>|¨����r�2�<ޣ�-	����{�y�pV��I��Zi(�=c����Y��W�(�i���	_�Ų(�H�0p���o-QW�������Jf͐��
�r����  '�}�N`���u�������r-���vy�0������qQ�B�$�͖[����v�KŮ�̘�S����w�#j乩c�c �ɋa�r���VJ\�ϮK> �R�T#�_g��&�jd��:+���p6Ý{ºj<��*�%�?�o�hJ]�XM�o<�V����[eۿf�Qw����.>Su����5U���[].��z�j)5غC��s:+�� ��)B�{�S�2�b��$�R� ������dhW1����c=:�3 �he�T���v�7ǜ��ͦ*TEb!nA+G݁��4~����g��	k�.Ջ�H�T�i��*)����?���z+����	��2aX2�n�!��j���������m�E�z�V
�OݫY�N]�bb�GCQ �l�Plȶ(�%�[9��t���q=qI��;*�9U_Ϡ��ib����_t)��#v��ǭaH�y�sU0�sx�P=C<�:��s�:,��P,�c��4�S�@������q��C���8�����w��>�ӹ�A�w��U-���47�Vy!�Z1#�i�4�0=��X�(¿V��g���}�L��|*_����O�+^��אE/���%m罤9mL�0��|��-Zoe�В7�A�}m�1����re�AH�ib�A_����c��F)���V�{�;$�΃dk/�
n���Q��XLoIjV�U�� ��<H����ԲhLbV^��\�WxE..�CS��r��l��~�b�f����"8�d(�ݬ�*y�3���K�%��D��B�2�*�Q#~��±��'�w*L�]ˈ#�E5��H�mf�9�?���yи/$C���뷸��L~_=�n��c�7?��̜�`_}U>^�O�M��h�AL$�� �11u�b�O/`�i~�Vr7a�$��f�lZ5|l����Y�@�A�p�-��
0�J7�S�w	&d@�APrf��!<���O�\,�N���Ie��̎m��Çh�xk3������[0uqꄊl謁}4G&9�JUT��kqA�Z����׺FMk	H�iK۷\)xU�X�TR��11����r��of�$MIs#1�O�0%�%q.%���ݗqxk���X��v�X7?�]��}�M��T�Y�xw�5`�u�����СU��諣����c�����hw�+�M����n���k��þ��.��L�<�g���'c {	5�3WZ�^]z<��r���t T͈���~7�e������>"�b NJW�nw�1t�a����% ��(I&��l<p+ ��c�H+�����9�)5T���W|h%г�vG�W�L�O�w��\�F+W�(�D�rb����!�]��ɰ�����+����3Y�]�3^�����F�NpN�g]D��8�vm�F�m������cxSU&���Ω���(PW!ɘ~�3_�4U3f��c�N=%B6B�.��m�����e+ҵ�u�䃹*�E��gLْW���J})�]ؒ��{B��T��U�c'%��xd4�>����7���z��g#N>�����ғF3&OA�)�[�?������˹�"��ݶI-'6ذh��w�Ӯ�E�J�8iz_5J��@�%��!�ώ����MW�@!������v*&���*wn`a,g��UTFu��*i���8�K5�� �Т���+i�11��� �R� 6�-�T�"%�(]��1���{�,���9_NU�1��ĸ6���3���^���:&��,����h9��ϳ}Lv���G�Z�4�3��������3E���*!�4f9���<ʵ_�z�_d�C;�-3�Gꊂ,�Q{/��R��`%2�`��D�B�.��r���\�S�o�OE;Gi�FDP�dD�� �cu4p�f��T�>��<@�a�J|r�bŨ��S0��MGI�wG/���-E��z?MV��w=-k�&�Qy�C�0_���¤�w"n�P��0�0�Wc������5�!���yB��;)c��~��h�Z�F��)s�_�0�$$w�y��&w��0j���(j����W��EO�>��-b��'��a��2�\�`	F��]_X��mIz��౑�jEP0�P�-C�yJt��g�G\ä.��$R]�H#��B<���A�8C*�M��d�K0)lS�x >�<>���D��u��<ƶ#�l�yx�r�h��?��VfBR��:����eƵM�S���m�i ^�Ɉ�)y��Q�Ϲp�>ȋ=h�I;��4D� 7�~ �b�eԼ��FNlxg$������溓X��҆X��=��Z�6e����hj���ӆB�Ɩ]zq�7��yh����\���,���@�5�7M����i�W��O��y���n��8l��8d�+�4�Q�4!����U��@�־�z��XB䑙(t�w����?(y��r�΅�(��(~�yD���`�(j;�d\&�Iš*L�Y����#=H�x�` �l�/E�9O]�KK(
��Q/�'� m����^��j0��j�V���Q��x
�в�cHh���z���= )gd���g�I��?7�9��*�M(Uͼ�x��
�d�Me�%T��FX����7�r!���~s��W}% ��o�ٵ�]8i��j���-���)[%=��cVkW@arg�"��R��s�����o콊���L4�0�%���]yD��B�XZ����k�!EOoC,�B�sl�Ш����Ӱ+�n�)f�T���3�8�n�:�a�3��3���� �|$�����T��ߎ�׮�2�&�F���\�'3Bq@н�#f(�Gx��K-��Q�+I�'^e��gy��9��ʃj$m�G_"������x�"���0R%V*���1��]O��-Q�ήe���,�,-/B��%�ە���i��rw�j��h7���u����Ur�R�βk�r��K�n�M�;4?n2P��f�Ӌ4-�B��L�wߏ��E���@$�����z���@T�R�_��b�^���z l��J�m�/ʯif�G˓�g��� (
�e�%H���D���U{Ϡ�z������n�,�θ�����t��
�&\c�gP�M�~��
�B9��A����/��`�a�@���{�g��zx�)�detv��kDP�x�`6�2���Fa羥����ڳ���Z��
����F fA����IV}X 
9�寐�p�1�q�v�wG5��s�Sݭ��`�������E�c�v���$�!�����3���DM�/�N}��`���p�3(��89��Q[�������X����8À�����U���J==�X;�'E������_F	JV�N^�l~HԔ���	��R_�_x%�b���!r=x��e��@����[ǘ�e�f
��;�|#??��1M�P�5�UR���ߓ�u�* �Ĵ�A�t�-qB�";U#z'�ױX�����$�9�Ǻ	���7�:���F3h����Y��#�7M��CT�eV�9��p���ѤP,3�1�0d��in���@1����xgqN��,�*��lg���=f�i�\QͧV��b
;j�&��t*,��/;�:�ш�2�!ӭ� �?���7��-��������g󫀑�)R��l�gŅ���9�|�F�[7�����j�j�)0�9���P�2�ӯ�T���F�{Y`v`ۿ�v:�!�Ԡ$0b��k�}w�^�2g�59�O������~+�42 IzbU���;~Gv�ULܙy�-�y��������ҙz�+�Z��ppuMF[�����Z��*�gq �q����HA"�s�%�t(��kă�u�#ㅒ�v!�lGD(�`ꜣ·y��Z<[�E+r�'�;#H�伛���"�?���rՒ�{�=\�g�l=��U�Z=5�_Y�S���.|G��=�kڦ"�Π}�^1�X:hX?S?/<e�F��g�ώ��.=�2�?�7H��mJ*v��C0P2�.Ь7X�+�c�[&�c������TϘ�Fa\Lp�����y�S_:~��}W�:�0�U8L@���0�a�ȅ�y�R;Y^%��u�c�۶����/�o�D[m�;�amw�<8��4N�0_ׁ�L�	���D�L�H9�a��XM1._Ҩ;ڵ;VBy�KZ
}df]�HSԻһ�Fnx�QaЕBY�{�6/6�����cn���\VX�cP��7z^�b���>:�8�AG�J���c_��v�C�SL*�3�;��O��m�.��ξ�
#��	m��3���Xʯ@��B�U��[!�E1֪8������ڑ��(x��.�$˸T��L:]�Ǭ���ǂ������xTr2�1��/���<�a;Nl�a)��K��j"ڬE)DS��)/]�Q@D2��ϛ�0�P�VDrۊ]����[U��}䄦�<'/�=(�+�h�H�I�xB�3R� 'D�ݡTB ��L�G�!w�YB$H7ըxN��piT�qt��k_{�k�d�j@�Ku���� ��B9%��/��	Qs+���a
y��x_�P�yR���~�E(n��֟_��*N��T�4WF\9���y6ઃ���6��F�''�RE
'���U�ԟj;z�w���g�ZV��	a�9�S�\f�oḱ^��P>�;`̔�,���غ�*�QV��#h���*OV����2���a�l*5Mm���A���a�)y�/^�q��v�:9?S�y ���~#��d�|!�W3�_uu����*�R8��n$l��nH�g�d���Oh�Ԉk�A�^T�0����{p��jEŌ��Wh~}2� U������x��=+d��C�c�!=y��r�SZ��G��60�M2-{�	�9�����{���}��#�D�&s����8!&��ǽgA�:pJ�{ܷT`E�Vܱi��%����(�Os,�o�$��AݐF�z��H��71�.m4��2�Y[��KG��U��Q�ڒc'dG4�K�Q-��W���I,�2@Vu>�>Y��٢�ִ/u딼�Rp_+�x�����8[��t�@kC����O�ޡQ#�7G��F���He��Yo���m�<s~5�3@�R�9��.�M���{��� �![$u~^�^�맽�&��0݊�����tb�@�;�%�� J:Az�0ACj�zv�v:4�?� �h�	����<��)J����{W��%=�����%�Y���M޻��A�ֆz�i��V�!�
�#L�H�~��3���zb�h��'(��6�1��-��gf��tKv�m����!v���f�{�F6�u12��鐯�̱`&�۸�f��I������9\�1����������ˍzܤI�������E�����>��{��b3�o5��-�7Ƕ9��y�j�c�@Wj�z�^�7h4tp!� yHJ|��J����{�u"�D�S���?Q%9J��*�P�1���gS[<N]���pF�t���Yu��\W�j(���hRY��w�R�8��#R�B������#%gJ�s��w ;�r���i�;=�=��L�;����,�.A�!�K���i�jp����t��d2��3)�K���A�=C�a��Lg_������_�D���м����6`�����[�'[(30¸�	�\k����D-��`�v�Ǖ�XD#��{��.י	�d��)�B��S{����6~:��6@/A��iς���B^�q�U!s`�A��!՜0��*�����QQ���#��.إ%d�uY:C"~H�1�?U�L,(����������ʝU�B�V��NYM3��2[l�\�A�b�T5�� �{Ab|��\�v>A��f��!(�Z��K;��3^�n����;ȩ�:r1�����ܫ^f��/&:�濵pK��4o%J\0>[��@���)���n*�ز���HA�	����d�KH�x_c9F�����(��f"�W�v���8u,��7�W�a�W�R~�k�8����/�2	����\��^�L&О:��)��̈́)	j� AT��p#ꃐ��婏O�%7�N���/�ͩ�C"��V�5���dK�U�P�I
�9�n��P&�k���G[ܾ,�)R�s����s{�d�d�{&HST3�f�*A���Ȳ�
�!�ӐЩj����4A���Z�B�Tr5��N��%G�#	�}�?	�lf���=�bxu3�hv�(�w�����v�%DlW� >%�e���S��:��J6���}+X�mp����z~�谤iD����c��YY���ՓD"٠�5�u�C['8�'���l�v'n�"�������Q<�/��c<�eL�����C�����fa����'!:����zғ@�E�D��I�Q���q�&�dL���뎨���Z��^�I\�Y������,���j��ؐ6F���%X��=��HP�k��?����u�����a��uYK�-�i�:��d$N8�-�=��K�h�jR�݋��7jxml�Z�a�"�����_�R�q_D ^��mT�X/k�Ӿm�p����b�����x�T����3S@���L��5���3864H�R9"�ǐ1����?[[�9Js��o%9�iTV_W4�]�<f�X1�Ci�z����p&�Ҹ���(�X��h��$�8�(A��HfD�*�3��*o��k@O����;ы�;��,�$#�w�ø��3��fK.���
r�Y&/�	���[�Q[~�.�-]�0U�V�����'��k�O~|}P�/��0,m�d������I<
����!�����H�YP����mԙ�R(��|�G �Z���s��5�p�ݜ��W�d�}�K��PΖ���+��t��7j!(���%����Sh�o~���� �	�g�O<�s�-���W}g�5���r��̐��}�
SI�J6�j���������6g�C�򔻥yz��oE�`h,u�Z��w�+�R��Mܚ���g ��9����Y���(������vÛV�^��`����C1��B�z���"!F�kΛ!g�X
�/�D��T�	�0��g[��S�ꖻ�� x%OJ6������H�=��P-�E6�]��K��[�-��qr��pF�@�>
S�d�t ��e(��t25h5�u��N	�M�bT~J�.��#�)���B~��'K���4�=0��s
�|�䗅ŕt���y���HM�Rh|�9<`��=�$�����7U�P3��v�-�����D!����N��1(���:��gs�Zo�������vQ�2�,#hW��O���p�DC�嫘��3IlO�|k�c�_2oX�a^��'fp��Y�c�jܥq�p鏶3��A�X�3�
��j+�,yf��D�u]��P���)!�;l~,d���j�pÞ%�:(aw��X�e`��t�C���G����?���.0�o�.��6I~ʸ;l�ی�&�|Wu�C��u�#�&o0�<A-q3���_z�Տ9��X:n#�����P���\�h�q����%�ЀH��4u�n�O�`1�Wp�E��w���O��v�B���\t�S�9��8 kx����;fǳ 	�zi�S�K��"��\��)�'[���o�{�Vysĸ-��<�,غ�}�"rd��T�z�/�˻�c�[O�
4g$�w}��)� ��ZU˜�-;0a�F_�0FY��O	��+��1-�f���:ʃt2����Dq���ō���V˔GF�ֺ1�XG���qTYh�5@�xjڒ
sH�����ÚIoل�`����#F^}��!��c���%z6_L����W�~ٽ����◒�Bm*�̀��TUs��N���БU�b���X��m׌��Tj����	4��W~�g2�)�OX�ˋ�S9r?�t�48k(���(�V^�S�a��Fg�K���4�Γ��C�Ji���)�MI6�ž:,��-���ޒj�{�7�8Uᚠ�x~���km	w�R|���2�w[�����`,@��97,���H�T�@fS ��f��-�^�cG������jE.{B�%�$�=B�(�mk9�]"��٬��P#JRK���O�⛃G.w�n?D����11��'H�Y�*ңiT��R��?�K�Ѓ�_�R���{o����P����P��.~�P�\E8o�J9gf6��9���4o^�	&����#�̩g&UP�.C�	�J���+�,erSh4�y]6h_�IL���[	�pMoE��HY2R �)�v���3���٢ #�Ĝ���؞C�usT�a	��=A��س�N�+羥��Tp���ٖ�c�t�q?�t��k��h�Z�:9��f�[��I6G�<}�� X�Mu�e��;}��ֺe���U?���H��R{-�"����-��ft�h��9��Nu;SXCn/���X�b}!"�P~��nn(VG���NY�\�����e�g&�/J\��_�JVe��������q35���&��O��䛑l�6	:��ڹ�c� ,�=�A��I�~�3n��P��Xv�~�(#�A���`y��L+AS���t?c�Z�V��H{7���L�F,���Pldם?_񻿾j��vW�e$��O����S�zF���r���d����	�7�)����ox���\:.g�����"'���!�ZV ���R[����l�  �
��ef?l��4�c�>��@u����\�����n�k��97��ᱻI�ܼ�� ��UcB��.�����f(]=��4x��_#.���:�Y�9��V���84�.�H"d�`ai�f�Q�kLTg�P�nx0u~�W������n�㆕�A ��Y�:(�g�?z��	)눁��~�I��?HўTE�l��� ��U.��ReU-�ǀ�!�)��� �������'����0P��`�)(�u!d	ZA�5�ͱ:���cK��0 ���i�Q/����z���,,7fD�6!�\�mzܡ)���^�4�cBDǲ���"S5������	OyI�7�S���{�L���n�Y娜�h��&�����+�D$3	e��`󧏡4�7W�;{vty-��Й:~Q��v���y�\���Gml�z�U��]c<o�F���\6���^h`�����#��T�̈́�8&�/�ݠ�"�\�1M�!b�&$'�5z�S� <yU�f�����[�\"�>nm��"ҟ����}�j:<����d!FtG�І٬�|s=�����;s�.�8j+g��j)	��J˜���Y��8�E�2pFe|ip����H���pI��^.�@Q�u�^�P7>�S��e͒3�A��OI	@�3Xz�����qv�����|���ڽ�Y4i��L��}�G���}�y�Ǟ�sFM��~u��c��뺃��+O�;�tZ`�������)1�Iª��Q�V�&�=)q�qEv�Ѐ���V���h�.N b�+<y�Ы�1.W�賽����Q�Ȥ���K�P�~�����V�dgW���,�����0��U׭m!ח?� �RG�J����^�G?�2R�$2��7�B{����P�U�]��Ԋ35�T$��1���9A�L�ڶ� �9H�����c��Lv�a�h֘��a��q�&ƴV��LY�ݕ��L B̌�#������=��[ӊң���$��9�X}^�`����[�������J�YD<X�鷺I�����ve~�G�E�'�[Ȫ����gٵmp�p��u$�3�}�'_�u�P2Fd`Ν�;%�>�R(�^NJ��En��ͥ�<|�����7�O��{䖫-39&�~����_�x�I]3B�Z��{Q�T"[)[�J7���=� ��w�Յ?�2�l%�5�K�yV䵖(�B��v$���.���T:LmR���9BS(��W��7c(\��
�S��Z���]9��
E�ը��Yfؠ��,q�w���l��Y���ڛ>{�2r�(Պ��g�f��VuD�;B�+�v~��4���O��Q4�7�*�i[L5I��C��b�T�du��Jx�u���0����4w�`��?}I�����(ԏ*�;E�_�VOtǟP�nЈ:�M�L�?Շ[���+�>C[0R@'�v~�c&.5
s���eTL�b�X��z4]@�E$�s�V�2LC51�$2��d"߷��c:6i�h.WI�"��������G"���!��)���v��-���	�6�B���N�V�g�I�f��pԵ:qRqk�?��9,��ctr�tØF��2'�)L:�.�B�mP���>z���^��Q�T���(K�TO:\N�ի3��q �E���RQ�w�A J��y2*;U�2�e���q��Ǧ-��$�[��$����� �O}�;�o �bd���$6�������Z�8X���W4�����Ų��ɢ��zX$Q`��^|�4ޒ�Eݸ��@Wl���� �+�'*P������/x�͛UuK������?�$�q=|��]���'!8DU'�5Oh��g���}娢���N`S�Fc��c+dI�=BpK>�Ǧf��)Z~J]f#W�//��Ԝ~�;2�����(x!�����m?h�X�/��$T����.�֨Cl���fl��M�%�3@2Ɩ{�mj��v#8-d+hG�DYM�~����<d3�y�z�*HT+��i���y���ֻ�輻��N�Hx�`e�ճUH��ˎt.J��k?�G����c7�MV�.uI��g�w���a�F���-8LP��ȭrD�B =Ԉߪ���es����)7/nT�����n��L8cG�����ie'Ǒ*Dz�_Z�Q}d�3&LU��:@��s�.8n_��v503��&l̀�_�+5�l8�h2��$���e�(_��%�=�Gި/H@��d��@>�����4]�f���C#\aZzC�
���_���n��3�ns7( �VL�Ǭ;M��}0@ŸWN.^ެ�n?e>N��D�{�b���H\����9���4�'c�u�Z��?�����}m!y;�$�T�I2.߯a�)�o��D:� �]	�J�u%/�ZSK��ŁZ#���Ymu�p��rkP(	)�p3� �������h���<�h;��Z@��k!�տ����!�׈�;����z@��_�&��,�8�#/gֳ@fx��p�O��<Om(C�V= �wd�	�zd���A����7�a�}WXK���nDGL����Kɳ����*�}L�ga����5�'yKX��;�p-�4$�W� ����5���M[umϑ:�H �\$��t��s�M��ᬳ :�_���˶໋8���ʞ_���]7�'��hV1��r��>�D���&"=[E��o"j|��ї�P��ʓ:����3X�����{k�F��~Q��{�a��+ =3��J�8�i!]�G+���Y?Z��n)�T�ȶ���<����A�f�\��y���_�J���7΅��|����9M�GKV�´X*Yi����nN�����(�C?�ɐ���_���\�]��6�N�Q���FY�-dU���Ld�ԡ7�Y���u��u"�J���pv���>�qa�Ғ4+��1��y��J�Շ�8*�Ҕh�`7�9}��f!��V��9���BF��K
Z(DXsM�* ��%�0F�(`wڭ�pR�U�fAĒ�nͳ�T�w4VؖJWض�ۨ�����d���ľ����<
^Q�A���S[b��>��(i	��P�Z,)&7�U�ȀM�L$�����1�<�[*�W�q��$��c�t]�9I�Ya/���X����$�n�@�^�.:+�ь�sX�P�������Խ@�y(p�e(>�E|٢fʠ:@�g���>;r4��'���wkl�Z!>�Hc��J������d*�f����4�v~D*w@�t�b!�b�o)b<6�Z4|"v���D�jr`E�C�K��2���RC{Y#��#�1�q�'t7/.G�V���zɓ����M�8���-�(J�z��q�0�;�Up�@>g~|���L
�A!�
ٍ�Q~ T����7�:� �����䧀�Fa�	>3�x~�:�;N�����pTh�{��g9��@e�vɝǨ���r���4Z�wa�m��>�V��&ж��7��c'��5b1/��a��D�Jjs���{C#`)AWxg
#�k�t��9����*HRE[�΍9.)��Y�OK/u�|�D����T�b�H����ऍ���>��
�3��T���+�����t�$3w��81�F��$d�b�ը(�챧C�0�X�IZ�U�s���,������z1�r	�z�&��":S|˼&����YT���6wh��2�9���I:I�j��x.&>�`����D��n�������hA���*f��E8@K��˒�-B��@Њ,� ��r��lPC��-&2�� �t���Ԃo� s�������J\�
Ȫ:�Ŏ�d��.�t�7��f�]>
-�Ƀ�v0�&|����W�����#�7��0�=,R^Vٺ�-[Vij��K\Y[����?XF����rf��Nbbw��/��`D\m0����G�d����
���T�tH]�$YU':�l�(Q��R=X���SP�!��;�ۦz��
��Ծ؏&�#���n�UQ�t�F<Զ\1./iWY:|�d#d��
?+�e0�/���\b���rQ�@���ю?���F*ͥ�/f�G-�/�T��J7�
� <f�"(eX+[�\���N2�)$վ/� �yϳ���`���K,������`n���M(�i�杕PE�_R=�������4�Aš�����B��(uB��Su�(�5���"����� ��'Q����{@���Jl����l�m��1�t�L����'�{�݉ .�/BP�-�g�;1�l4�ǅ������;\[����c(/ &�uK���+PF�	!��6�E0��?Qȍ5Q���UL�sz�lDFc��	��a��dB%	���2c¿C�H���yp�a� E���k�����b�٫������Ҹ��.��K�+����*u���ݼ�?0ŉ��0q&
BZ�|�E�@���y?c�|���)<��~v�e�yլV�ja`U�O��� }�烎��qh�d`��/n��'B?�,[����C�c@|'��'[�r�i�&c����m�L���}	j^v"��̵;!8<��bhn=E�nE�7�i��^���51��.=#X�<̟n�[�� z�ͤ1�*��B
��A���4�&ߜb��$o�&B�w�X��/	G.�V�J�DW@|���:q{^�l3���j�͜&m9����=w�ת�������"I�]�x
S$���n�/t�P�,�������7��8��w!��۰_TWh�,��|�O�� 7ޔ��s��hd���>A{��p�V��W4�f�_�Q��� �̸����r�(��B�>�����='���]&N���\�e��i��7g4��F���ƈ)�䗞yDd���l�gb�"�y=tȤ�E���w�f-3�p�a!�� ��ɦ9\�lg��_i��������,8�L :��š0v�X��d���*��J�a5[�]�K�����\�^P���G��{�9N5�5����ʊ
?�Zj�s�������	Ѵ@����;o�}ǌz=��n���nsS����	-4qar:�3�,'Z8/�m?������P��]����-e�%��k��P�q�m@jT�+lR���Ht��ld0��\�#;��S�	4�B�u~���9�xM{�� ����\��om��K��ѿ3��o���T
���\����B��8���ݛA�������ٻ0�h�6�o��Ka�\*���<��6w��o]D���:1�SF�n�O����,�g�'e��`��N�����M���
ܞ�G��H�b�{vO��l�vt��a����9�z2���+�oݬ5
^t���NZ�	�I)��~�|��6q�Kd�������J��?�g�´D7Vp�u�������6&9���VY���x|�է^8pu���]c�G9�TN�,r�\Ü�E���ݚ�*	p����] �p�w�F�b�|Z�[��d	���uyyt��(Z�M蔈0ӵ%M�R`�����nk°�~��Z5!k�'����<$���k�QU��]���a�P��>i@��_�U���_���1�^��,[MR�m��.Ҋ�+B��>`ʦ6C�+*Ʒ۝��L�kL�d�7�βͽ&�2�Ȃ�{�b;|�Gz�J�ȓ6زY�#�#�P��6��|I��>�H��뎎�˟����S'E�8�3?�{ 9*)��Hf C���l�G豚	�Ht"+���s	� �g����yȶ��+�?\I
c��i��H5�X>��ρX9�~9C��-Aʼŧ���蘾�	Y����U�dn#+���oH��hw�&\d\G�&1�2��p,���5d�Ų�VU{�*��n��s���/Pq�N��d5i�� cl��۰ s���1��Q��:��z?��r��Y���o����`;Y?�j�D�P��e�2f[�w'B��o �e\����8���x���8k�t�3Rߐ�)��fI���>�;�"h@�b��o;�M�j6�nF�9��p~IT�v���j�uvrd���	�d0�?�pxs��辷"�`X�ɒj�ߺ��Ϣ�g��� �~�6-�k!i�䉃=�nTm6ѭ_<�Ro|�V�f8:l�~1Hdeսb����Z��TX>�* `�o'����BYz���-w=�V�8����ր�;2��-,�!N���e�'0'C�2�q�צo?*r�lKK�A�T�
9h��'[�����*O,�!)v`�?�5�'��+���s>�:�l�%�L7�i(V�Z>��6@�T�#���8/��w'-�`��k6(|��q�H�ԕk2�7<��n��l��]� �	RJ��lzz զ����d��I)Y�� q�����~���Ⱦ���B�ï��(4��Z�\.vF�w#��]��k�`�X�ۙiʕ�!���� �u>������ە3t1��Mh�]	��G D����t�HH�9�Y���伧ǉ��q�q8o�*��I�/�:�-(���?�	P�m�&���_�I��
afo����i�*��Ƕ�o�+�����C�R��X���|�ڢA���u�&��V����B;���}>�X���v�Ӟ���܏8�2�j�LKv���d��i"i��+�/G&���u ,�A�B�P���t��i�PPW[881�E)�����7'��}*`-?����{�	ͭl|��P���~Ƞ��0p�]��As�̨��''����u�L�%@f�R��L�xn�X��}�.���j�5�� �v�C�m�A�58%����S9^+�X[:�9�=�ـ��<9Z���[����5x��U^�#)ܟ�+�z/���S��!k��y��U`S�E��b�{|,�qA䑡Q��l8@��ү}Q������Y��ﳲ�e�� e��C��#�zu�u&��ϥ��,���;��%/3tȵ��	�aĀl����b��P�~0��{7�֐G�o=t�e^�1Vγ�8���I�mB���ϼ)�W�a���9���PF�Y���P�����$tf}jO8��?h�fX[ g���ܫ#�đCH����R��B�"��b/�Ą�L����S

�^���&w��,��F~#�I�c�F�)	�*^�S���f�;L{����ĉ:Ϋ��1�rdB���= 4���|���ܒ�
PT�������"&JC�G�j�x�_����[[%�{\���-KҒcU��FF%����&�g�d�i����q:o�B��;p�^���ur��|��>M��Yp9�*�%F`�Q\K9���G�|Ha��E�v��iwseo��% �:��F︇Ϻ@�e��n��^��}��y�G~���qjF�\:�M�;hW��T8%�/W^�����:s��7�x0'u�BX��!cJX��db�"�	im�Y�5̵�=���0��#�=G�A�t%A�I�(7�A7+3g�b`H�.s�d�H��ւ�h�Kj�*o�Oa������y�1���fvI���U=����:����=�ȩX��2*GD�D?�[<������u�y��v}�N�|g�Va�r�;���h츖�>i5������f��T��I!gI�������+��M�KJ���dzgY.욖�7j�eڻ�"�0)��,�����9��H��/�\�P!P�fUM/��#�%<ѭO���Bsa)�*�9��o����/�����j�t�Z��V�R�T	������:���e�����q���R�ߥ����9Xj��r2f_���9��{Mܟ���#�wkUp�_��%$�u�_Z�������Z�Y
^2-m/�*��V����V֗�r���N�N�ޥ�ē�;D��(�R)��E�F).���yy�����׃�!�{���}p0GT�ۑ��'37I\+��f��>5sp�xօ�K��w ��@Ws��߱6pgt>H����ٔfx6,�C�xtV-~-N���F	��]ړ�0L��=�٠�֥����t�7�u����Nh��}Yu��e,��f�{Vlc�j�	PH`�'à���^�ϼ;S˛�G�X�U{ BQ����b��f�����*��$���NE�p�\��1�S+�Ю^X�c�f_���ь#�B.��5��@�$O���5�$�e�/�.��L	y���	�!�I�OAA\��[�\~�S���:��3j^���i撘��C�Ƌz�]]r*|n�.�|��z���x]���hDƖ�|�F�����aB"�,W{��Ȓ/pj�K��;L�������_�g�VO�w��+5 �L��M�a؍�<&6�d�;eb�;e���ܔ)L2nUkq������8j��u��*��0)Lף$ ۛ���X��ib.���cO�T	����'�y�R�����ݾ¯��#�� e�=-إtd#w�ߓ�X�����9uea5S���;Y�o~}ll���@J$�n4�u���
 �E�6��0�%j �	����V�S®;�-�������Q_��66Ƈ�U��R΄���/�_�9��ʷp�����yܫ!7,����P�QO�>���:G�]vgѿ��s4ocOb#.�^����n�2��r�K?������PD7�U	j�C�:�x�h���a�I��[���~JY�Q���l��t&P�"�N&ջ �����s!�/����)�������k:L�p��[��^��M�P�u�d
 v<��#F���� �](�����1tqv��(�86nrh5:�MyF���`���}s�p�{� {B� j}��U_-,�3�����K��pR=�7mL�C� �T�G<����a
kd#4x�&w(>`���]H扮�}�A*����2�s薚�����"�q�b�$"���oA><<��w�&��|+zi�7q��Nb����̒���0%�j����ݩ�v��X/�j�_��3FI,��}D��N[��殌@b%�we/��E�Ͼ��Hy�*�7F�b6U���7�9b�U[�~ғ�,]0�+uPYv~�����`S�QUEMvY�s��8����zm�����b��$��<�O��-��a���5n��UW�<K���jS<T�~=�D (�F�iܠ��=�yh����J^;
����W��y6|W��0|\+�Ú���d�ƪ$u�1g���}����s�`�2��TwPBΐ]-��$6D��ܖ��7Nj�xP�Y���:���kkXM�0��(̵:!� ��� j{��,��g/��\�i��}��b3��6�O;.�DT���~�F��8�l/|��O٦H3{QP�īٟ�^�y�z�O�S.���٭Di����a�S�8���b0�7�.�^�֥����C2���R��
a�B����p�Մ!.�V��sb�!�	�����L_��Vc�Bc�*��{���/4�������� �f�����3A����f�8#^�z\<�@�6J<`&f���8z�9�n`���@k���,���$��E�If��~j�ݖ��ny-���n`�<qt��W�����Mm�cAP�#�U(]������b�k��/\��33g]p-��_`MT��UA9�)D2;���
bL�(&E[نd�c-]�矗���b�ȏ�ki.ԯ9<P����M����O�m�W��WD��+��bI�I�]��qߧ�+��<Ă�^�t�m�QM�rd�c�Sw��U�yv2���V�S�K�ր1�L�sb��c<� IT!�H7���a��/�R��`�7Կ9�Lҍ*�1��QZ@`S�<wJ������m� k��Ɇ������	�w�w
v�ǒ�۾�r��"ܓ�z�۟)�G��),m�B��/	�4��ё�>��C��ud�A8՛|��mgiz<�7��~�aA���m�m��ci�S3��n��� ���u�R'N��b��az�zh� :���k,�)XH�Ӊ��h&nw��]uiUQ�P�t	�:�Y��:NPO^�@����vID"���{h֑���:R?.����'�� 3g� ��*/Q
^?���-bc��������<��E{J��Bj��jJ�<W����6�������P��� +�s��Î�ޮ�B�A+���0AD�����>_v
�(�N��{��Tm�5IlM��5/q�� ���ܫE-�ZkO��^*�E�������D��V����\�Lѹ�q[��ZƷ���S&�)�y�+���ޝ��2K��d�����)˔6�R�r��z�;0��ʂ�\�7s���� %�2�آ�E�V
^*�>�[X=Sz�`��7ԫ�xsg�
�����
�V��i9y��(�gX���G��4ELBT���;Y ��,�#�j�6ht�Գ4�ɔ���<6Xc���.��QR+�&�s���LF�KBQ
�ā������:�A;qn������c���J��%?���'��:HVR);�n�Yb?Nh�aۿ�l
Wőn68�5�t4�}z:b��)gP�3������/		^� ��y������F�!��BЀ1�yj@�0qD��Z�m�=D|m#w@A&��a�wCU��\��)����N���5�B:�����'.�P�/��lkM9�Ӭ ��(��3��c0�y4B�C�:j�����	�u;M��d��R�1��o����?a�,�]�d�jf|�B'��g
���} 5����b�(&^�5f�7T��!{!�Ob��K8}��U�ܞ�27l�-��˼��׏N�*vJ�f�^$�DlU�) ܉Kۆ ��C���"Rza��[(4���������)D�©T�?9�?�b1�6�d�_�/|7� �|�tX��&�:*�q�1�t0�o����L"����9!�.��r�µE1w)�	��ēQ ��T����T֖�X���%%�W�05+o��떁A��
�Y�X����Ě�[f��5f�wM^�4���W/�t�A����JiV(�lT@E�Wb� �O�������A��E��'��q�9��O'��u8���9�ԡ%nɚ�O,�#BɅ�5!�4d�<	+X��>[z�(a���� _|`��`��k$j���;�_1�IU&���0UH`���?���o[�2G&/��5�����2m���V�:*�ɴ������,�;v���c��Y�;�-F��` Έ�f�F��n+������(Z��%�+ot���8G��,_��>yy�$[r� |�cƀħv.ಽ< �--�1���(�|�#�;�`z�g���a������쓲j����+� _��1�n��DAc��=Ve�T�d}tj_&�8���@���K�NQ��歀_|M��1�G8�[�9^yz��Da
I�I�@���x�R�
S��t��=He#㡨C����ױN����C�\P-�*���9�eL|�
:��#N�-؞�l�8�F�e,{�w�����6i�_�[1ExFJ��nq�����:�?�8���f�bVV�����K}�S�h?�<w�U*�Pj�U�vB��s�x�V+��V �>w�����S��ܒ�?�$H�@<CXz�k,[Aͽ��EG�q��bӶ�:�	9^�g�� �^��+����~k ����ݛ�]�|�̯�QOb�ܪ&6�k��p�%pv�k�54�g1
B]� �����Aci�b��1BG oPa��vqt����h�o��=/e)��7�jEҬ+�y-GKJҢ�C���Q�wc}�T4�pR,S��?2Mb�"���Zeo�l2�/��|��:�]A��kŋ�����n��Æe}ɶ,���1b�k��;9��T߸2�L�܋���{��� ZZ*��м"ڼ�?1��͏�w������$a>{�|r�6�F ����]S�H�W	��	��uԷ�1��]U�����}�RX /4O5�#�u���!c�h�p�7�iM��X���sy)�6�l�}�.]�O�ս��Uٖ=��1�ZL4_�����Y���{�3�3U�(�ә/4D�	����߷��Hhz�~�!�%7�Ʊ�_pۧ�g���6��J��r�ĬE7�l���q��
��dկ�}��>�+�x��*lvu�i����}�Tj"JE�K;��ը�d�A������
 뫿-���w(�ҁ�]�Z',[y�P\Ϯl�0��P!���rdQN ����+J��UHx�p�L-���aM�6�'�$-�:l����UfwɨQ��#���^�_l#@5dj`�3~Qh��2�tU�~Ʌ���$u�Ȁd���$9f�3��;H+j�Pkj�#.������G���=�@l���O���໕@�C�X�B�D��Ksӹ��@�N�&��*T4QrG����Qg�a��8�*��M+�����$��9�đ.��ܩ�?*�h�C/��V����� qa%b�|-Y����T��������<R>A���PΣ�6�Sb���3��5�� LJ���&�@��cd�.�2��D�h�P�r�W��9B������Z���P��Յy���N�c�6�!<��y�
t�c��4D�s2���7��ÑY-�!�F@^o�����K��a�.M�e g����G1Eև�6q�%����e���,�x���_G��V�Ŏ�2�嫤cV��N_8�0��ް���r~��E��8J�a�0Àղ�����/3��"���r��1�{?}���Q�n��ē47�D��0��3�<q�~ ��k��|h�p~��z�gr\}�S��gd�4���LL�L0���4�V����mS�r���ja*x����������L)S��b�����< b���T	�6>k�E��|7�~��ي��iQ�U���E�@w�Aa�X�%䏫����K��.Z�`HQ�ɺ�B�.(ܦ���h#]W��eOr� ���g�N΁!Ò��׽�W�4czsAp�sT2�k����"#-+.���F6��zl�E���O�,or�Y��A	�)�r~~�3�=Z��E0�	/t�F�ZP�2��5EHv�J�_\i[��g��Lv���S1b�-�����f�u�kE���Y�<pS�w���5�)�r�'Lp	u�B� m�N��ڠ5��ѵŕX4��ۧ+8�p���٭��tЈNw�����(��F�+���ɤuN�D ��M}���ޚ��#�H��`ˮ����d&,<�����:�=�������I�F�2�Lu=>�A��]/�{|�|$<2ڕ�'� #1�L�>l��Zk�k�ma�N�� DQ"�
^#�S>���"����������K}�@�NOQ!����F�r��Ŏ�R�)Y<޻~�V�q�"��c:�¬q�h��
' d��S5uӄ����C0_���>���˔���1Q�����duR\`��o��E���K�a9�Jj��SVH��]!.5xC�i�����NY�o��7I�_��5h�ͬ~�X�7!��I���z�Z��]C]�Cؖ�����%	I��|�/�&M��Ƅ�-S'���Q���� C��*,���z�$L��n#�]ٳ��L�S$Sr�E�+[��B^�(���G�ӭ����]�QRԪc>�P� ��Q�3�N�s���r<Ek����T��d�ݘ��~G8��$!,�639�1���cX�dn��+�#���~��S�ţ�4��g�>����S��i0|�tqߒ�;��/�g������M�NX��Zv���8�mC��͟;�y1��0�C^r�2�������P�_��f�6"[�����.+\
uP�/�:��	�d#��xߦ�{�ǵ-N93�Ƌ�a�(SY��o7���a=��� ��a��=ɰ�i�HA�/V�N�F���0���Ƶ��G�'ov�3�إ�e���E�5�Y����!9����Ů߲:ٶhE��P0��X0"�ּ���*��:�zr�Kf7��h�����M�zR-o��+}}��
���h�n8�r��lN)�C
�/�ْg��o�
�A��n)�/��\3p�/\J�J����g���2+Z��Q�2�Ch���F"X�ze�s�oyn����F���G�f-���ZbFJg�PYb�{�s���XUݑ��#=@)���ZJh<��}�.�}��W�D��W���=� o�}V�5�+:�����jgJ��׎��
*W��
!O��W-B����㧞��D��/v�v��+�LFY�/5�N2�8Z����o�#GN	�q�=��󈋕U���܊U�
Q��}QR��{��E`AJm%����B�#j�\�h�NJ3il2p�i�C �=G���v���ܴv�=��o�CHJRqP��'Ѝo��֏���Fr1b��s,��Ef\�`G���}7�c��i�D@	V��N�-eM�P�S�����DXf��y0�.�=�)�s-���7�0��/���B���|xR�����1eE�@u� ��''�;!r�y���l����Ɠe���&�q�|A�f�cSH��(0��1l|�����[���7��V*X}���|{��se�2Q�p��]0R�Vv����\��ڹU�a��H�1Š�㊨���Χ�p2ON�ܲl�j��Rh&,��{�.U9�>J�[��P��ѷz��� Z�n
	�5�J��0bm81!��+jC@�_�ε� E�qR3���8�@��$,%�.s]'i<c�f�/zo��Mb
n`���[��C>�ȟfse�ɛɵh��ٷӦ[ê7�B_�J�?a�f���vM�w|���Y����q}�<0&P6?y�)��2alN<6͚�5�������-ك�Y���U����|h� dOu�*5�1������n	;2���n^�L�dEe�C�շvF�K��Պ� �.]��%2%���!r����cV�DQ�\��MFNt������@�B���:��^�¤f�,x�=dUأ���M�DF���9l���^m�l�=
���:��s��K��*���+�ٝ@�巺�+�O
9Nؐt�K 1��|-]F����p�B�裝Z�痸6������6���ĒX���{O��f{Oa�ŷ2��/������&�T'�Q~1�����V�^ߩ�ʗH��Ӯ�Q}�Aq>حQ���Xv�.��cVN9�)L(�
N��^�
l�IK���\�e�#8μ}i��!����"��a0����+_�����^SbC
���VaX,�<�,*�q��R�g���,�]l��L�1_}�2����#�L��W�;�ǒ�ǯ�Kǥ݋zC����*���W�4hc�ot��Lkʜ�~?�<�!y��&���S�����Ͼe���`��Ee����U�AJu�Bz)u����'|^ۃ?�^sG�w�&�i����;5��/�������m|�J\7�35�e�-����K�Uf�.�屸Un�N�~��l�ǖ,;�$�i�e��:���ӃGΔo}�4�.J�Jk�	L���-:����>щi�\��f4��'f�N�FλO}`b�IE�!Z���3mA��!?^&���(�[�6P^�UyRc���T*���[`�!��%P|��>ޝuDBc��4DU���|7�])��`Bޣ�`g p_�VH�!dS�&�3��Slr��+��Z�C��;3g�<A\����h�;�q>��lK��i�.N%�JR�A��I�^��..���niJA��i�v��6���I���7��|���:�"��Y��Ԧ!��JN���p�B�N,�<���2��8#uKhl�U�x�)I�I����O��b����H/�6�L5M��\6Ƭ�R�5_$y�3t3N�(��Y@�\<��t����n�V��-V���~�mV�Y<�X!@ƥ\*�U��o�~
�q(����!���;�'"XLI�B����	;w��6�E�r���<��i�]ڕ��kɁ\W���T��ǚo����Г��8��L,p�8ԅ�R�$ q�s��n���x(`���{:��e+��#H��������e˸��x�s���[��pe��?ݝKF�<�&�2xBh[���q���o�D��:,���
x�"�`x��[&N��������f��\�|4e���d�6﹥U)3�5�S�+_��/l����c���fR�k��+�؅oV���Z��_�P���do.t�����q�4Om{�\N������Fy�	j���oV��k�!�����˃xwLi��Ο��N�G���M�SpXpq"@�s�7����(��@�e޲?y�|�
���UTa{���v������h�m�)��c؁����d~B)Ƭ�xVG��D�l�����f⾞�4����s=�ߒm�����Qb A@E�1u���	ͩ�6�u!!�)S�vn�<wm�z|��WТPPM������͗0R�H�7���n$#��/L^�<Dݲ��S�7Mʡ�F�I�J'�Z~�N�XU���=n��`��	�2�W�It�)��ߚ��S
4t#U�QK^���I�-&��K�r=-�t��W�� �I�-�Y�(J2g-m�u,�B�������/�8>ܟ��b
�@���6O�<+�ԁ���d�M�K�c�Ժ6x�C2�Է�����Y�o�%�Lؿ�ڇ-�@-�[V��W���)P>��4�U(wN:'�:�5���`+	�1�>�o|x�rI�_�:9���kG�b��:�&r��R�w'�<�Y� ����%���t4᧍i������%hܺ����	fW۴R�����C	��+
vPU2��vp����d)�C�&� ���P��z2J�s'fN�_����E�~�ʪ�-V���d�ÿ
0�|�CSi�Wz���@P�QKR"/�E�W�݁U�n�_Tc;�	Z�75O3�
H�������@�� �\E�b���Pd�g�0o�z9�iq��[�E�T��`e�1�g>Ǎk�юg�Z��oc~D�;����Lm���C	J��X_��|���W-�	)F�K����$���!�'��<�x����2V� �- 5E�#�2	������$���̜�����X�
K�%�K	��g1s߸��p��p^%��K���5���Sq��:w~c�o����g�ҐfY�I���K�.nWVL|jh߽`0T��^"I��v�&9�܇:�gy�Tq�[�4�q��c�ch\�o�%`f ӗ�7JQ=�_F~�?�]�?�'�c����.a�����b%�)��E�,q=Ge��?��D�>m�S�W�;��s�B�ov ��iK�k��_�	�g��{2�1�0]�A�Y���ai���`%�ʷ0�B���c�����ʣY���F���K�p�ӣxt[P�`f��A-y[��ӽ�sh���+�&�������}�'�2�1%�{
ճet��uj".]�s?������L� 3�4��Б�4J��$�����@�o,q�)���Z��_�z˪<��s쇭Yv�7�$R{|5Q�`��[(bU�4�ȰO�u�]妚�H������g%�1k�a`b�Ik@W!�BR��~��AC`���`\������8�g�T#��p,��>�	ex�B7oE��ʃ-A� P��Ù5�z�E�Y�/�sM9��K���zK��=l̿Z[��Z�>�*�F"3�����5�F��ן�˓j������"�Q��Q���1!֟=��ؼ��Xv��S�Aޔ��7T���S����R)��A~��_%�%�v�$躜�g�$���0�̀��2AA#
z��A�.�ȏR�,�A@i������cg�祦Iv3��B���PHW�����.q�([���!�8NV���۝�].j�1MW��m&�.�������G���Q6�����)�/�࢕�&V��$RV�ލͰj+�o�D&���������T�c���^.�G>�]}���[��s�ݮ*o!��t/2}���@�@�kXyV�%�$� 0,FT�_R�����z�훍u�O�S�*mVMF�s�A���Aa"�<֯[5�H��Eƀ����+Il�q�╌�8��.'ҳ��'Pwl��Ѧ��S.�-��U���Њ�K����@عN�&�\̡�������������������'xy������+aJ�'\�jg"�@���u��B0�K�S��sw�m�i&Aݓ��~4�W|�-�lo&4
�TI Y��dc�Q?� ��e�8�)X#,��GԦ%�'*.�������1iD��-\�l�aU"�
��rqu��#�.��٤L�V)�m���G��8"�$Wl�仹�̃��R� ��ߍ1&�Q���!!�3�UNϑ�,�ޗ�9����b��	h`&���i���85Hk����(s�7�6O����I.�V,e4c�v��f%0��D���"�,�sU}�\���{q��1�0~򶔰4���i�`�S�X3#�5����S^W ��ֵ��<�f& E�"�� ��F0�6���i�f?�'�k�,�m7W��*�p��X��*#�"�\jI(_#���k�>��N��L�!F�0�����Ei�"�	�+G��Y��x�Y�L��CiF��RO�������u,;8��wʺ����_��u�"��6G1-�g'Ql�'�`&:��l��R �0�4i�����Y��v�����!��!.�;��n�t���M�b���>2O�E6*-��bsyqE��c/���"�Z��H�06^�T �5,����������P��0t�{���h�x�ۻZ�#�	x�8��I!�7��o�~���q��-��������CS�F}?�41��>]!���-�������t;�M��%W��;g��M�߿�|�
�]�ʾE�k���E��0H�������lKʰpA����g�ef%;6�bz�k�P��Ν�8�*�f�Q4̂
�J��@%�RM��Dx&#D띉�A���1�":�S�T�s�
�ly��% -�K�~�Y���c�f{U,@�d8U�,���|7Y|&�;-��~'���Yy����-��T�5-6�~�đ�����8Ġ��
{��;�3.���'�0Y�QmVkV5��J��UbW�(ơ5?<��Ҽ�7��b��w[��RX�I�V�]Ǽy��0���r�����e�_m���8�#�KLv�y]�wu+�P�n�e�~ULS���秌�ƌ��HC¡&�6�G7U����R��q���q�EQ!h��͜F�
K�<�^�؜Bpv�7�$0�������:0?������'7��A~2"�+�^�r��k��^B��ln�4����je\J�����)f��[�yP)_�[�$g|J�-�+,�t"��Ӝy�T_��>������E�{N�p�E�g5��J�kە��h?�lͰH��R=���3���c�kB��1D`����p�m��7
+������o��quRՆ�QX�t�@�--,t��o�$��G`���X�{��L�0�>Mb�s�"�;��_�����]v���p2�?ͱ�UB�<lKX����j+�q��!�����\��[�>����Va��*s��U&K^��
�:sB���/}2��l���sZ�&��j�����ȸ�.5���0Z*&�q�U����p��q�,W ���������Dg��܆�� �959ƿ�(�� ���̢����7���I3��d������6]H5���> \��H��KI/�h���Ǎ�b����HT¦�act@�U���L�qu�kI#������y�E�x�팂�H�	�Z�î3�|�s^���([�Y�A�E�d^�˴��@LxyG�tޮ���}O5,RV5���>�?�Ή�OYᅩ�^*#o�H�"�6��+��_��b��|:�Ώ	�m���Sa��H�ֶ�'V��3E|���vȕ��]��<��?��޲�Q��q�2��ڭ�h��F��&�
�������pb���+H�bt'��g�#�W*�2X��vB�y:����1��2�&�«O0����g��|��p�����ۯx��4�U�;VE�����Au�h>����we����n%�Й&0�sJʜ�JH	���Z���vs��Ӈ�����i��8V}�m��(����� ��#j �zy޵lvǍ�[V�o���ڀ(�
.�hc73�M����r�9D��g�i��|u~I	�2�Y��zhm�����\�ڎno��"�{8����L��,�7tYҊyl�a���P����n�j�A�_��ͧ����;�0������_�ߑ-��\���4s�L�����kI`�FY��ək�^_�c�o��8� �H��rC�vm�#��Tի�S�*��>�Ua}	�T߫�~J�L8|b�x�j�fKYU���ؤt���
2ބV���C>�����\Կj��9[����-�!Әq�Sړ�e~�����D��5���.VL/cM���_j�خ]�S��961m�?�C���	�'�rNR7ta��V[�r�r^��.��dƃ��7��Q��e>�țxro�u1��y܅/[+�ԗ�w9�����Eݤ��f)����pѲ`-���S�.�����'P�}�Q]`y�e�rr�eU~�_Z��WPT���3��S8�R��v�r=�jf�8�E����~L�߮Iq|@�6|{�dE�y�3[~e��-B�Ȳv���	��H����I{���]�,1�v�����բE�l�M6Y�7H�A!�y>��S��\�il�kL^R�)�f8<��!�҆Z8x'o�E<xʽI����)��v	W�trj���Ū����FC���}���v�:����0�Mx��v����	.��wz��l���̹mJ�B�B]l�Gw<�u�"-�k�,�+�(r�W�u1"L>�#�?��Ek#��Y�E��8����N��CV�B�r�O��o�%u&�[_}��Ȕt�Ss���$����=<��P�Qʤ��TzF��)�]��cQȾ;-mٴ��@4)
�.�&�>�
�|\nbvC�N:��X�,D��gއ��o����72���E`-��H6��=
5�-]�P$k��A�
��{f ���H��t�ש��.�<	�C���@��n�0�MJO�KiĉsT��1�I�<7x��?�xc/޲F"/�R+��u]�i_6�L��w>`����6rX
��*�*A��<$��9J����S��'������*���K� 5�R��Q�NCT�;�����J�(��)(VR q��	�"4��J���cx5-�l�ڴf�~��>�EY�&ٮ�4�Ȉcx�A��v�n� ����u�!D���ވ�\7��)��g���I���W;��� Ј��0wA�;2�v4��b�ˌ}�ϓ�:S����=؈;]o�=��(�Rkѕ����d��*W���FȐ�
���r����
�Ӯ4���M�}J��ҍ��G���,�|���,�i�w���#����}e7�ۍ�5w>RQ�)0���@X��~%G��l�E@����R�
ib�Y��b��V�+�l�#X��An{��d��� #X��nh�,���t�C�y��^`/�2q���tea��Ó�ɉ\���1P�'m�����n�p� �Ac4���c�R�c��a� ��L~I�Pb��&h2Z����_ r�o�I�R���>;���`�D�~�Y+z���hO�(]̀W��٩�W?^�%�o,P/L��c���eޯC'Wy2�3���H���X���Pu���v�]c%0��|Q��]�2��O�R��JnxtyF7^���5��sS6iAK�W������5�:vZׇ�t�$�JMU�g:q�5�cg�O�aϳՑ6lă�g�k�A��[$���Պ��Y1�M�}
0X�Y��7VE2��pVYoO�Ǚ�~p��F"P��O�x
�:��<z�C��v�5�\V���@��L�f�2(ʱ������!�&)��v)4�߷$D�HiF����&��.k��C1�ǻ�{G��T�B��-ѕ��!��Y�Uۃt�OԜO��֏���?��V=��T��K�r��K�*f�~�*�.9?��`"����H	O4L��k���j���k�����
�0?k~���9����.htrm`�x|���S��O��.���ܗ��)�������KȪ��TCvϴ
P ��4#!�#W��0}9H��[R��vw|�o��Rb�5��|d,�`���<2~��#�A8�TJ&P��07LXGb���h:�	 ���Ti��(\�d��Gu��ő��J��T��_�]�������a9r���q��:���PR-E��O@��v���D����2�X�w˧���[�\�7d֑�u{O}�jKB�Su���CxR�Q�l1��{��b��LYwb?W�|Z��[IS�;eb�qa�WK�4��������ݪ���g�E��Ax$�ns�*/�#�����b�>T����҇=UTቪ��W=ک�н���	��}��=yy�B����z�̂���n	��+��&�C��y���6�{��s��e���gJ�617��ج�Ψ�����RJ�!��t@z�M8�w��c�:Ț�ͨ��
"�`h�2���F�[_	�g,	��LZ������Ό�q�����V�S{�����y��|l�3�ʎ|yʽ!�3_�&��'�--d�����7����9iΑ�A�i�7��>D^�.���_�P=@l>�b��5��'&5�;R��V�.�trq��֊w7Ҽ�o��Z}c�Phn�a���CYk�m��*vl���n���z����,P1����Ĳ�z�m[�4��yF}�<�dJ `�w�)A�3[�dK	�Z4v*䉵���$!L�)��k���G���Ya�ŽM/��wCT�)Z
�B�V5U��P��L�%h��i�9Q��b���u�Zɝ<���o�3B���q�ӳ~Wl�#F�Q>L��f�ngN�8������F`��y���0��f��Cj�8ln_å�_W	�o%�kYd%0ϨЛ�~�l�u�)�Tx��x�/U�($��!�-�՛���V���yL]�vn7�(h��TiS�ֆ�Dk���������K�!_�Wߍڦ��/B�ԍ�B��dmԒI�Z�^́����d�w����/�P��ݐ�x������]4�辏��Ð����N�w6.h�<�Yς�Χ�Փ�v���8��~��;
_=�I��(+�h�~��곃̻M¶o1 ����y�m���E ��(�悅�JW�f�NI�s,ʢҘ��_��Q��-V�s̞xnZ��v9��,q,LJ&.����\ϢR3�nŜc��@s�P��L:y��aL7f�%�t�Z�O7R���r
b�[vFҺ�e����es��wG��bڅ_�|�L�0�	��3�]�~����w.�cT��d�d�:��Q�Q�s�qN����;ն$�7Y
��]bT�6O��L�p��b�Ώ�2X��v�)�f�#�;~��
~��-�G�{�?n�	�+�9e��y�=A�T@�ӏ1����==뙶�6���X��?͸㦏f������ǝK8�Wf���f2S���D������w�Oy�s��^��e�z�X��Ҙ�%iRá��}���g��Zu����Z�*<���ߔ&<-EO5"��>�n^-���ěk-�BW�n2Gtg@�u5�[޿�q�9���{�<G���8��X�1+?��q��^r�8�����A�����y����Xi���L- s����J��Bl�\�O޴4��&
F6V@�r���߱j�O~��"��e���#B��A�}��.��7q_�
�,��d`d^�<W�����U�r�������i\� �xRT"��M��M*��o�	o��7T�*��� o W,�!��-7�o�A��O#��6������P0�x�^EET�v�:�+�j]���=������DKI�34���M+�sShn�;�3p�,��SΖ&����C8�B	?|���7j+�'}L�7R�"��=N��Ͳh�-��C{��BS���9�����PQ�����z���zպK�Ao���g���<�QƇ��'����O�(J��M���JO�T�hB;�	P�0?7�0�L��
�������5���:����^�߾��.��/U1��L7Vn1�u"O���I冱�bvB,Z��x�7�ss�	����<��w/K�viV�-̍Zk���G �0�h����/��z�.�ޢ����� By��4u2��Y�y!��b'g7�`�|�7�����O��k�_l� �����~I��W� c���
��,����_a).K)� ��<����y��-�+��ݻݣ��9������xG��e¸��|�*����@Bm9�0}�#�Y���;���+l���˱�0�ǃ�)��l���
���3=��U�<��+�Ih��?�=�	b��~UaEȢ
8y%��A���@��()ؕ�6���6����4[��J&p9b�M����l��xpcV"�&�2d��#Eki����o{Z�[�D��BK����pt6��es,�6gٗd5���,7����\p��*sC��Nw��Y��� ���|�7���.�r*��⦴넌���Jb�\z������)-�,遊��(� dŤ$7�s�,�?����r��氀0�g(}�Ɗ���lwOW,Jh*���n��i�l���Z�=���%�?On��F!��0�� 0��B�JeS��;�N-״nl��5%����>5E]�p/\kѷ��"AMz;�#��UF�[��a�� ��_���~�-�C�샳�A���ʟ<ַ͓� �r��VB�̦��C\����]\\��E�\m:��C%ɲ���1j�^�	�,�z i�U�#	g���y:2�� ���)�i��y�l�6c�����b�np6�3���s�|������aE�}��ժȿOq���N����kT�k�UK.���f��2����4�M�@+���v\ws�K�8[.�J��!�-��Qh�~z&u�q�������,�����.�!K/]�]�S)fX��p<����#�V�}C���
��𪈫d%���0��EU<�������=�9�@9���`�%hU������)w����f`������6_{��.�#�JH;�� ��k�#�hPy����k4� $�2�S"�k������E�[��!��GT�H+���c��%̙z�M"?O���3V=jv�rO�7y��������gJ��x�(�3q�OR�$;�����X��A�|������},m/�v��2��?�F�l�-*aXBO�(;T.�͗�"Tܱ+�
��G-�9�޶$K}�B�T��y�PC�=n�������(Gq*!��+�<T�t塍�z??��_�v��C��O��{Q���P��'�P�6s�	��O�}gc��"�E;��Lم���Է%+�]�E�M�r5m�F}��I�z��z���94|R�2�n��Bm�= ސ����ƼɭC3�u�j7*���B��c<K<n���9A�����e�Aӣ��+��o�NB����r�P�
�����`���"�;81b�"�������L�*N%�9	���ޙ��{�C���#C��U��<�(`�^K,v���-cM�n��W���� ����R V�$�M�,�����&��;�*GIN���A�������/�{����kd�/�4VG�pW�h���c�dVW#�`�M c@��dT���޶�oBEx?|U!�c�Y����wAYs�*�HG����<������j��u�|��8�q��6���ΞI��;�ƈb�r	*̵�̥���^�ܺ�{��T�yE`�H~1�� ���Tu���ߥ�f� �LkSݠ�������&I��?��ߣ��t	s�B�8k�_szަ������<����T�{K�6cjS��)S#m��{H�#��d����6��ď�++Q!�>�J��iO�4������K��>q4��ɗA���^{ВW�M�l�*��,�7�OK��Uޜ��>J�X�r�RBcɁy3� ����ʥ���!������JL+�۽1?S��T��nu�AOL������RG0�mgL����;�gW�)�c�]���3SG /m�����-gM���RD�����2}�F#�=i��{��\j{�UYh���V�n������6P�ܖ�?���F����~�}&a�aSҊ,�7'��,*z�u�E��^��?f��[k5-�F=��üw盌}'����c}������Etwب��1�J���<䱢�w
�k>�7��mu�����N�\x����p-���3�bzsT�˟츛:�=�DeDP����3F���R�;VS��^#2��[C�͙�au�B4���Fh�� �.���A7S�Y�#js�7��I����d���B��li.���*����/7�}f�Ą��0���82��x*M��N���\q���̌���X�+���U�8Y�u�#&g�|�v�*}��P�x,R�+U�7��a�Ө|{>4����H���t���õ2�%p*>�[e���]YO:B�{��
�(u<�x2�&OSIe/cn<[�R)%ڲޥC2N�Qtq�'pN�
g�*st;�����G��<di�e��w������rŗ�B2������_��Cq�S�B�x��&	��@�T!䰉�uL=��%��ϱ��AUg��������FB�m��3e��.kT��|���nZ�u�~(��E�i�7�_�� }���3 �"�e69�Rl�c�l�c씬0kI 	��������#��i��M���6�L�L|S�Z���s���<�>%4��fb�����]g�H�|�mP�,q�; �鑃�����#<�߆fT��1:��$˨����h��t`鴕�4=q^?�8\�o�w8�A�8t־y��$=���~1	�Ɛ�z�%[Gb�r��QD#.�%�T,C�"��
�w�B��q?�x�Ȉ秊2b�n@^��w	j� ˙��rӊ,ߖN�P���!޹�=�i�]�m���^���V\���E;�����X����@~3��:0�M��\&�a����"/�#����=���iN!��N3�X@}��sPC\/�&q�Z��@zH�iJq�>ޛ�������Mv����h�<��xC^cp�ѕ��%�}��(��r7�`����wj�^.��*'�* �qOJ���S�tGpBe�K���9�b}�)�@�1�$R6�㨱�kd��.�O�Ǯ-�S�,e��Xh��$���6c�آd�~%��1֞3wMd� ����(o���{~24ա6�B'P[V�H!&rŒ�5� P�ұ�G��m+ޚ��&�+�P�d�s
y҇#�_���4�?i὘ֵq����	?�Ad�^�@�m��*C���<�I��$|���R$vE5�Y��� -V�z��r#!��*6�Ք}�)�'ک���x%k�#�+��A�[W/x@M��=h��%:�3��'�E�Oc��@1������7;�VQ��0�Ee?�Pq�}{�m/�z=#��}�����\S��A4�l���i�]�"��O�8kP�OL���>\Hc�	�BJ��싖��&QՇpţ+͖�Ԝ��F�ʮx4��rQ5C`y�m����{$�˕ �����o�'^N�9�����$��kIF=�� �4�@IZ"�=N/��u���H����/Lt=.����P0����`������R��0���C$j��E�	o�����2��!j����x�h�/3�p�?�EW����^����'���7�a��o��)-�������@�g�z����n�$f���\[�qS�ޯ2�nX�!�xpU��V�yE�x�aΏ ����y�(H�������j�ݸ"�)�� ��L{��?�3�>�Z�<Q�cu2��j�N;?_v~��_�gz�M�t�	j�����<7'S�`���R����\4���0xQT3�=�>���g\]�_��l�o07�*���7�;(������L���}l��d-���:��A�X�;,���<#��:Y=��0��e���3�jC�����B�㉡�Ȣ��I�b����|[�s�
�fUY���l���`~��M`<��\OBq@=��o�Þi��{�I	OD�&+E�g���m�L<���ãw��n�>��v*JQ�s �)�D�A�����uH��怡�jVh�;&
$#l��n�g�??�l��'Z����xN����=���N*����E���ͲnK:��t=�'� "v��>�6-���j��Eg�J�-P�l\��z�&wI$���2k�޴Fp��S2d�O�
N*��Ů'*��{�q���(C���BzÀѶT�L~��,��rB2�e��D�4��Ǥ�A{䏫AD�_�0L�zn��(�X`&��[� ���d(5��Hac=����/qEnV�����o�6��&y�:�ݱ`�(?@
 Va^��se�"��,��EאU��^@{����+\SQ�W6���/"�hSZs����h�,r��fK���Ԯ�k��-5b�g�Д�3	s�t�΋��lm�^bK�o,�a��(Nt��	�\o:w���^���\� �&w۬6��8����7���;�F��8Ͻmn��œm���Ơ�C�N��-��z������̢��xI%�s��<���I�?�ɵ�:�+v���?���r:�$�Ȃ>�:�gb4&�9ɼ���z^4R�b�B��֍G�
Zڔ��_Vþv�۹�Y"�f�B�E�|�e�wu��f�)ϠNV��)�X�{.�ֻqp�>�J����0��ք�&!/����N?����T��?��T�&��X%�1GBmn�R�����&�E2��>XrI�+E�~��E>��|�&{L<��V=x�|{yez� @���i��]t����T�g���^隻�2�2�E:�(GP�>N�E�����Y�}�N�[�4C�S9x�8��~OA�$�����U6�6C�P���Ɛ�̮�v��uStm��r�`eI:Z��F�x�:�ݎ[��q�ڨ�N=��x�� ?��1���8?V��fh��0xCR���^��K�b�
K8�&���@2���~G������j}T�Ov D��d�P����y��7�x��,����ؔ�A*gYiH>,u�ň5Y�dH����+7�vz�Pj5��F��q@H�7j�Bg&ו�4��;�0���I��>'����xqI ���
�0s�� ������`����^�ƴ�|�{�a�nВ�	�,s�=C��r�󾏆�c%��Uˁ���V�n@6^6�p9�Nn�H$M�ia��DsGu";�������%�p�r�Uc?�����t�޺�}}6�⍓b=��?D�|�o�o°�*j��$��g��оS��K;���o!�*����9ǽ��N���PJt�]�yRx���O1}mtn����)Pi��̗��|�4��z�� ���7��yu����M-����X�u�#���<��֩�&+�9Jo� �wx�㳱8K|�/��*�l��;�Q:�11_��:
�砼%�(�AY��de�$�d�s
�Q�hEa�hWW��p�_66��j���&̠�$\�_
i(F�Ug��mx4�r���p���AF>ln�協!Z�&��@�q���}p�by��j㣍0�=iJ�!�ˍ/[+,��L��g� m�������i�ύ��V{{����|َ<�h���+V6��y�B��锧���<�0����IPm�O��8���E9��IrH�5Z���/:]�Y������3�����_g���UV���1�;�Q���XV�ԑ��K,�؍3i��DbM���#�8l�j�(c��9sG��=P�f��������R��+ѳֿ0tZ�d�_#�AF��qKG<�A8��i������ZX�trOǺE|a��Du�K�-~��*i���P�brh��̄?��C��QoH�.I���g��E�*($�[�(����1F��G��bEx��Gd�g0�e��I�i�͖��N�Q��|.�\M���J�E��'\�>���O>���`�X����em����vס:H���cF̜���Y�%�����@�I� K;��f�R���Bf� -F�$��E���=��Т���!=�{��ť:xъ,��G$��CA
���ޮ�y����G�x*�DC�ʻ���+���t�3��u[t��^4�ْ���g��<��*����s��L2��:�˂�Wqbw3�&��eLr�&�F�Bv��������U�N�?���)��O�^����
�>��m�g;PG8geXH�����g��׾�B����xQ���j�����pLni�mM�ԋ�(m����U[���撊�gN����}2��^6�g�UP`cʎsP_��(}�#�Nd�+ŭ��;�w��`,4g^}��&.ٍ�Y���z��T�q�Pv�s6K^�y:d��
Š��-E*���\�Z'	��r�"�#�
��;�k�i��g!�to�G�w	�<�n-[.^��t4���3h/�7�-y�a�C<�B��"*n��oxe�����[�9H�O�4&=3�R4]k���(.������4u�8:ҘlB̝{f�͝N��ÈH�Jf���,�k��h�����QAab���?ܠ�W缱�Y>�4�z�_�u
B�~�O'���l���g�V1���� �)웻OQF�������:�����_PR?;�N����^�@����jMw�B��s��$Ѷ�Z&�i��'~�!��11�F��I��k�I����͉Χ����s[\ă�08d�	�΍����?�n�z��	R,�r��6#V}�ێ������?��/���K�%6�0�3b��yė�0�A��b��,��^�ԙ� �^_=�{�jmy{�{?V�y%=:Ȧmvt T�(PY���|�����&���5A�j"�>�u�htRQa��y��x>������z���c��˛ᬟ��"r�� R����6 G�Mi&��׶@
,���lf����-����BS��E�`�/M(�WD�>��xz���U�n?a��.=W�sk:ϴ���윲��Y�Ǆ�+9�2�Q5���)w`����z"�xJ�f0���K������L���O������Iz�<�k��uz�i|X���M���3fA \C���َ�`|�=|�&D�p~`�;��l�y9��"��p�����f^K�j�.Rm����O�fAN�e�]�5��>j�A�2c�ؘ�!!��攏 �٪�8�e��֋>5�2��B��{r����doղ-C�۵��Cw�y%�Y_p��]6[m��;����	�����g�\B�״i3Y4)x�[!q�H�j��fn:�O��� ,�\�2�c�Z��35z|r�̅2�����������T�̓����_y��:�i��wŔJZ���ܜ���%�;Y����C��g0�*�;�؈�����(��<�Z� V"�$��f�����z���z(}+i�6J��?�o����w�����{��/Ë��q�X�쫅�.V(�ߛ�
��/���͈��Ad�u���xS�.�Q!hwO�~����lu��V�Z��9��BrO8kx���a�.�wY��=W)o2��2�X��~���S��WX[�A�}a��3ogVO�>��̎>Q�8�'�li�&SSW7L��k���6�/�B�|n3�%��s�.Z}�;���N�b@V��!)�o�5�Fp�ϾY=snP|e��e��^�2EB�?���0���En��ș�:�""�`Sp(���^����v��Y�	�X}e �`�(� �����ȓ�K��i E!|��ǀ9O��m)P�W|�@����u����$CY��P#�4v�l�ێ���Ap7�%���,��؝�]nڀ�y�0*^6���}owS�����9@$�5�Q	�*�ӓF��@�mk���!�����ˢ?א�x�r0����>u�"�����j
����ڹ��ܚ�u�T�5y�O�+I���6qF��nܻ<V�9�M*yl� �3]E�9ԍS����X�h̩1�А��6t�]�M��nn��oJŵc,b�cy��?�-�^裡Y&�� ϵ�����5��a0����sȾ�5fk��Į'U��uEڱ�v�� �i\F���K=��+.@�NQ���}��J���s$���g� [ǻ�x��߮�\�ۉ��e�[��!]Jj,��K���[�v�&W�ǲ�-���W,�GHvi��*���Ӊk7��kGu�\!�I%��}EFA�u�)��(eQ����Z�&���y9�K��ke�����LZ�t{؁Q�\|��]LA��Pɣ2^�ԎI�M��p���/�������@�# ����*yi��	�bKW5,?��8�=z-m�ͼZ����T��y�GZ�U�9)��]icG�$C���:�䎆*5�\�bm���>E�Kd�
`Is�#o���h���ٷ��4h��ֶ����C�;6�&���& j�G�'h�K�r�)�ub ���� wJඓ<�{����w�	|��S%2�ϖ�82W�_=��m�{7��t��@c����:��-�L��0���6������1��g��%@��6/��5[��랝����|O,���WŔl�F�^5� ��$���	�k��b�Zʨ)k����?"6��Z����Z��� !��Ck���<�S����uI�86>�nf$̠l�	��Psz�?�����7k��ý��ChW�g@��:��a�l�H�sEt��/�-<^Ij�� 0�'2�+��6������5jt��[����I�GG@}�N�>¯��z�B�6�;h��h9>��ۓe휗@z�C9;"��.>������!����n�ުT�O�������"U�M��!�F�@�́�>���P�f?wytF�'��/v	���Q��-��@���&��n@��톲)�ct�}�m��AĪ���c�9jH���[�	g���9�x�r�r�N�fs�Le�z_�Ă%qG�,t��M]K��;��b�I����������$��5�G��qC�D��[���$~�����u)ה�p2&ĿKT�5�,����t���Z�J�u�y�E���kjg�[e��㉎�Xބ΁����)/ �	I�<�~��#F����pĒ��Cq���ֹ�̅΂�R��}��Q�E�引{�G�/ �z�h�����.����[2^I�Z���s��*W6|nz^���g�D�fB+A�B��U�[��U�޹��ve;���˔"�I$�H���S���ܯ�z���ҩ�N�g�-�.��(�T	��m�'�}��?���EWE�m�?�fQW J�\&�~yN(�d�O[|����&P����2fT������kNt>9)�	&LMl�̿RR��&rjU�mL�S�B�� Хi��bϥG���&����3v�s�&p9G������?�x?ȗ���u�,'��@gK���mGz�vj������Ĉ�O�|�gP�t�y�LU��5%u9sgTl�X�Sn2�5�z��)e+Y�U@���5hr��������Ԡ�^�� ¦	�V�r-��t�߹&wݎ	T��,��s�"'0�P�̄�d7V��I����^Z�޳��g�]֌� X��5d��ˠz���"���_��O�Mk�ǁ�v��/+��[GZ����>Dlj����P�w���,
a�l�>��c�x$HG��)�5(�k�L\��+�o�k�O�0�2�ï�7�}|1���u�7��W����W�����E��Ʌ�BC�Pͷ�@��i6�r|���s�����'�ȉ�66 K'z��u�@xl�VJ�u�H�R�Hy:$[�w |�?#�b�n	b�~i����%��L��|�I}l]6iJ���]]SW6J���0�~r��lV��}�k݁EVW(a��cv����֝4��Cl�
�1iH���@���$au�5��7O5
���Gߺ���N'��#���ȃ��X�}V�!�&>Q,���)v[2z��iA�p��c�8��6�ZsM��3�v�Ruk�O.�= /��;.�3偳����CK����E?��b"�P0z����C�㭅�ATӛ�~�6��s�*���gq����U��p�?�ͪ�5�JR1Ⱥ/�U@wk�?��HC�(~ #�p��J�:'Ń�썶�oS�c�V�9��C���ߞ����ϱ� Q*�pA��ңE8?`v�>��A�@��`juaP����k<1So��[EƮo`�@�&_b�$ٛ��U�yfG�"g"�_�Vm���x留���f��	K�ϰ��n�Bt�PYq��h���a�)Gĥ�L�eJm�P��#c-�)k��Ep�����1��j��_��u]�k�!��"0�1�s��Ge�`�������d�t2�	�Wx��a�(l������߹��t��*(nY��fÙ�g���$�,F\A��y3L�b0@�u�sb���_T��'.���7�P�2�#��I�H���,f$����}k}G�NhU�6	́�w���Y�)�8�Ȼ�^�,D��GQ��g�\���5O�_x��2POcc�*gI#b�'�R~������A(Um���@hg��w6/r-�х�yk0J���BF2q��R\h����<q.T�ْ��& �aT�⾀MՉ���Cf�k�z)����9���������2��K�L��:o�{r\�䂶4����;$�@ѝ���8��'9=�XH���"q�~��������\��J��ZЖ5�8<�C���$s�f��a�2M���Q�>�m������|�޾] ��Q�����A�~d�Âb�sd���L�b��w|A?{[`W���^[�bT��;����ͽ�	��h��]:����3��74u����&`����q�����$��`֊�ھ8�u�&N��@��4�=E�T�?�J_O��ǁ��wښz�s�vS^��S�Y5kJJR���fmJ�ӎ%~N�e�T���c�:Vw)�$�ͼ�W��E���d����&�Rk����y�GA�B��#�X"�f����i�r����_�5��7 t���f�_H�x��~��4�"���`v�Oj���l�G��jI��Ũ��IKʒϸq�Kp΋�}I�U�_\`�2�}�fhg�9X���к,֯r�Ƅi)��l��z#g�:����E�W۶Vi��`������wptqX̪�kV�Ҙ�[J��h���rݗZ�I.�Jr9�H&к�_���J�H0�z�,|*�ܻ��\+�#����)%f�\T�Ĉ{K��k���ۚ��#<��&��D#y�o��7��g���x�����B0	i�|�-�.'fOq;�]Lb��v+�&�ˤJ���_�(�V����w��"�U���,{=-�(B��|�5��./��/ ��t�ʂ���d�Hz�VA�0����A7�J&?Zfv�(�rS�NMz���B(9�_�*�0�[v�0b���<ā��T_�I�y\O{�6��{���1�:�@������r�Q�|���6�zw�Z�*}�ׅ�0<*�]7FN��n'����٤rS�B�( ?�Fr��GQ_�ۣ���J�f���y���Ul(�Az���X��$��#D�yJ$,�)ޢ�᏶�N:'o*�wU�F��-m=t��֠�>�d��˶ٵ��f����<���!5^<۽���}8�~=ќ�u����ߔ)���:��Xl/v�TE�� Ђ��@v���\��2�y�=6[���#d.��x�ʭ߱iKJ��wv��^i�5�zT-T�_9zģ�K��κ��{�j���M�Y�(@<�(e��&N�S�-u��o�8�$o&�LN�1��/V�(��ձD70�{R��ث�O�P��{� p$Eܿs�\��9�f�qhH�&����i�5�11xK@�)��v��x��2$��t�9�'���%`k��!� a��SD�y����"��1���A��f��<����MWP�u[�L�c�8�<h������ߔ��5i�8�J~,�Kbt�\�]�a���D���k�a▙�}8�W�g�W�Xy����:x�*����r�]9K���]T����l+}En�A�~4)1�z>ف��jF�|��Kmź�N^�\�r���E���(�e��!��O
���A�-y�Y�E��a�S@7&�B�_����\��e��6s}��e����ￕ�5��4sgT���!�,�<�ȴ �G�1U�������l;Od0�]D�Fڿ̔K���/��>���=������D戎	Խ-2�Щ��_�޿Q*G$�٤y�7��0�F�2�Nv��ۛ�)0�|Ӥwm��8Le����ʔ<�*+kP4�G�ȱ�+�-J�C83p����a�CB�;'[?
��W9�5�=���ݡ����S৩��'ޛ�+���kD�ˉ�P51ɗ������z��Z_�ɠt��0��&�s��W�n�$3#aD�[����o�z.��:ǡ�ψ�yg����^����;�le�Nl�y=F�̡
��,�H3��m�N悕^�]�AV2p�����[���bϡ����X���e���"��N�UQ (o�����x�J�#�Oжr'�����(%�]�ĉa9�c�O`�HS�1��vS�d����ryz��֋+ǚO`;!�A�Q@_p�ܸ+(�[�h6�ǫ�v&�Vh]��,�m*�L���
_� �.�CH�P\���T���imn0����{�3�>�
�����_�~+�Rb8�3��ȿFp,ȖJ.֟��B�~D�e��D�(�.A;��e,���W�9�ә��g��15�k�nUCȊ��"�NaPc������xNh' P��FEyW�� E�'��Zc)�����=�i��rڏ��j�H��fK ��������+��(�|º$��,!��_�V�2�Y�!SCa˅��[%�֊��劶H��m>�/�Z����;fBy��v��s���������UpIRm�.=T���U-6��
����QA����� w��Yl��Px���#	t%��kU,�4�.xUK�҇��L�("�UKy+�8�Kը�P����x�ٶ��z�v�f���/��2��g�X|.�O�s���=�����>&o�����mi-%�S�<��C���+r4d�h����&D��w��7uv'����T����� RȭI��h���.�����nO�G�]o(�/�o�y� �VJ�?h���-!*�Z�V�A���A��*�	�̮�	V3&�}�^*+�@��w��јN6�,�K.�蚕o��.��+�c �&^��Ihh�Oܺ�d�
ӡ^��?g�����1(uf��(�j�WfR<8�:�uC�����.o���I�K'�{H8�6��Ed�R,��3����ߡ1g���C��q+S�J#�Cr펛]A�S�|��zЬ�}x�� ��g�u{��L̉j��Hʩ�*�RK�}�iFf�ے�t�"�\���ce��+�c����i'���g{��U:�\�̅Pn6턉�B4>��8�ޟ]|&��3�����*����Zզ1�o�愤p��>-���s��g��,&��z���5�����!�7�5�؃3qz2t~��LV�5ܤJj� x��R�DGf��	9��kJ�J���ʲ�9{naL�j�Op��w�)u�%��eɹK��� ��O�Q�t2�ѱ��,��.�YZ;� <%��6Ѯ8�%�T[(�*�{֝mV�P��J�G�l˨~��|i��]ʠ�b'�ͮ0��xL>M��bC������#I�N'�R����Ws�@ǂ�r]��-��y�sڨ�7Q�N�f�N�Z�� DS�e��Z��5���5ΐ����+��O��07��X�)~���g��߷���4<�/O���͆ɋ�z"�v�(�E�r|c�95Q"�I��T�P�EFҾ��ۆYa��0v8��s���Hj@:6�C;��C�LǏ��~��^���g�6k����:�K�=���������ē��"2���\Y�����vF�� P
�k�1�8���B8!e�����%N��ҟ.�Fm���"|�d�B�4j�Q9�ӗӯl�#���yVa2b���� 8�'��V���1G�"# "�� �S�xg����
�����q38�U��R����+���G}N5���3)�]�9�b��J�i�"����w�V��Z�@4N:�ؿ���8�V{�v��C��S��g�^x�9b2@8�=�\:��%�@3�|��x�hE��q�ݗ���+�ـ��*�v�>2���cS��uc�?t2����C3�7�4�3���g�NU��*����������k�Q��\�n��_@�ro���z���F�1r:������ok����+�+epj�m����@�d������;�l'�$`���6��lD�[���l穐sSKA"�P9.�$}�RȖ�?J9�����@����<��r���,��\#�t�do��I������ji�{�#��Ҙ��Q�6-�ɡA����"`*����̒W���9�x��a�džW��&��t��*jp@M�V̿vt���<�f�כ�+Q�����ef�K���8���xE_�!�K΍^��Z���Aھ��E����\�O,�q�[w���P����Ɠ��zy�X�d���|��H7o���acZ��F�����Sᵽ���b��?[f�^Y�1���$�H�aiX���ae�܀���b+�m�����Y��ԲOr�c�'�@���X��,��	
vB�����q���x������~�]5������ú>h�(9ĸf}�,&|��!7���Js٦J��w�|��2��u�g�Q<��拯Z�+�G>���7���ښ����hl��|�k\�z72�Io[�۰��`{r�`2.&���' �Л�~��=nh�^��;��G����Ri/v.{����j�v����D.�p\�wj� -t1z��	��o�^xs�ۀ�mؘfu���&H�OC�3D��s����̨�!M�C�ͷ[_��%_��:^0�6\Ia�"�Q� `j�a3�L�6�v��u)��٦�к���T|`��|ד���i�i�r����s�`������I���5|o�A�eCH��8��E��êꂜ��}ܨUȌn��!t��]����ǩ7{�ٲǐjt����Q,��BK%7�7z}�^�u%�h�R��*3p*�Q/:�����#)�����vy����&���1����L����ϥn��TI���/�'nŻ��c�Q�/���i��EkǏ���=Ѐ�o�f�~�*e�r��>��IUތ�z��s�:�k|p�O�/����%�+���;��c�Yo<}���
���6IN�=�E��?������Brd{郐��p��4����Z�B��w��LZ���=H�Ev(d!RX󀑎�+���3Y���{����v%N5�7��^�Gm�x�����1�T�0��	l����݀�<�nzV�y���T$f..��L ��'E�\�r:����ߌ�*0�u�����0�H���4��Jm�yY�0����5`��W;�;ۍ>o��7GE.�NC��.K�7��vCzg�gS�䨂�V����\�=8Ǘ���4Ik�^Ò�{�Ԣ�ppۿ ���!�U�a����?Jr�����s�n�T{�����yy����ؒ��F6��2��4��Q|�_iwg\� �:����T���`x�'R��2x�jEeH�.XWit5���ݳ�(�xv��vr���,(zI�Mъ�L�6h�'��K�ȉ�0*H�b����� {;�wQN�60���da+�{����6)�6 �� |�jM���	���n��Yކ��ۉ���8	ōS�����b�^Q �u�,#K���y�֍C�L@&�G��2o�7���eY����J�3����b&�����(��0DJ��:;�����åFJ�Ҟ�z�/>F�����3�k��˰��FVM&�%�����S�#;#��$Y#D-%�='u�U���ዡ&_`�i�/ɐtv1�­��㽧^H�y�r%��:վn��M��R���U�;���amZn��qM�@7�N����,��Y6r�q�z��כ'���l�����8�9�F���F_!�����Y�c;�탤���A�p+q/Jf�_]�<" ��"��CX�NE��ru��yE+5CJ�[��.J=��G��Č��G��j|0�n��)���׳����.tz��Wk/%��'�$1-~�]���7�1R������D��2�������#���/3U}V,��:��y����<pBh����l��C�D����(�ܟ��r7Ǘ��\�8nI �bL1���2��@E7΍�n��8�������6N��n�e�vU��ݕ<0��s��&�BQg�v#���ۊS��m����z��q��p�QW7�0%U�iGsZ�������_v��`�FB��##j}�7Ҡ�;����Q��=0A�A�V��p�/yiNˡ}�jH�e0M� ���{�c�R	�/I+^��<�8�b>AW� =�!��|n8�&��0��9�T�q���ɍ�6��O�1O��L^m;�c�25��=P��`�^����s;(�����������M�魱����?�4��*��L����G�ؚ��b��E��l��H�o�q�0kn~��6\���$�ȵ�1�Dk���vM�
�ӭ�#:8�3�^�<���ȇL����Rq�R�Fĳ�U���ms�.�P�Ni#�/��-�<{�ͼ�I�R�4��T8��A7����w�:��A$�9�E�pvi%�����C�WH���w�ũb ���3�Ȁ�Ƣ�1沕^�hY�9�\�uc�pZ�TgU@I�>е�Tr^$i�!7֭�?p<[���oWB�R��mI_孠��g?� �2�%K���$E�S�����{�$�����]Zϱ/�o����
���kФ7%dvN4�T�ԉ���%EK���'
^��_�ֈ���|?�\���2(,Β)�qH��}���{�����'��2�s�(����O�,�����]���썰���k�ѵ
7<��+wR3�}���\��G���]Yg�lf�/M�Ih��@�³(���D��7Q�CɈ�f���[����ID�ʷO����̴�»,��y�i����V�q�M��@�l>z9l�T�e��Vg���/�@`{�-4i���(��̬d�iR8-q��%-Hd�nz���+�|T�^BE8wT��)$���HOL+[=�	V.�2б��BN�O���YF	t*�l�XQ��^@���$K���� �T������dTp�=��G�
e����c!z��K��!y�����*߾
W�T'��_����F7��UD���rZ���,Ү17�=�\�h���w�
�ivZ��}j����:���O��w�6;	
,� ~E��RT���6ԭ73�dT6Z���t
�Y��D��4u�c�׊��:�hV�(��J�,��:�+R��L�w�F�i��O����E1+��E0{�ǸJ\��e��jq+�~�'�*��+�ϊ�� n�ኜ��y�'�R�͚�L���o������9&�c��7fP������q�u�4�v�ȼ�lV��k���b݊=V��R���l�(p������b��sڡ���W�cUisCr��ܭ�t8 ަV����
(&X>iL�����r�n�+ʡ�&OZo�8�أbs�3�#[���M*�A�ViGJ硜���^��f�iﯣ|�?b�J:].�V��Q�R�ч֦�	QȠ��!�=J�D`����xG�4��ĉ��p0	-�m����&F�.aT-$~>R�����)�F�[C�5�R��+�a�����
\+Hgn����M�Т���Z�t�F�,�E \�:`(���~��1����B������
R�����'OY���J:;x�:!��[�7�+��̓mx��o��Lw֞���
b��<:�y��0���.gd��E��ID%z�lA6���Q�c�<�n2C�A{��F��a������|W�-G�b-�L�e�������<u��h���LMU�d���.�VRK��>@�W�I��_�x��+��Kn' Θ�/jZn����UX�9<��<�X�\j�|��ؘIg���vۣO�����u����~k�:�k	_{�ne�7���ĿP>o��6�4&3	���!�y���>�w�ԣim�t�&�o�%��2Kω���+������G�]`Q�OhL��@�b|V��U'Q��zI�+8T����u����7�ntfu6�i���@n�q7*O$��Қ,q�}���8̅3ZA�x@��θ>�#�s���V�8��{�y�ڿ�=`M����7���ZX5�ޑ��&�Ij�A��iX��t���O��7�G.#�#��f�8E�յ`f�yu�֜�Շ�?��oe�ԧ��$�����?/�O�w����XR䫘b���R��E��ױ}>��	P���/�$���������C����d�����29#E����]�{�� ����H���ty?D�}A���k�@o�'�@�9�����2�X{��K���$@��@k��ݔHe ˏ�޿����	�H]0�F�l�׀�:��%I��pA��1Tp�/�+����e��ԧٔ:òh\x�K���y��b��é����>��N�ev��rK�%pV	U=�(�mS4�K��?hͮ�q��3���H	���C ���1e�)�Ѷ��Y+�JX�#�&H[���)SIm�)x�������Ǐ,��Fd�ӪF�;�@��s��8&�lJ�c��hU~dY��{X^����ۅ���y��]5%�� 90j1���bv�&�RDP�uC+}d�,&����}) g��`C���(#Ц�u�?��gcu�U�DHc��х\6�����)�)�s2�n`'y����Ɯ�4.J?�}@�ª���#F�����E`f�w�ɦ�v%NxY9�/�H������v��2����l�!Es�󲴓+)�s�~�ˈ��-qu�*V��d�F��=�`�$���7D��P��w��3@��w�X������ǐ�"l���a��:�_P�6B�=�ԑY��� �G��� �R�,���)�tl��Y@�kU~��<JI,q���I��x!!F���*�=�yހ`qT����lf<W\mG�����TՈ����~'�G�7�2�{��8L���N6���F�ʇZ�[�*�m��؂��Nf%fɲ�_r׿���u�����&%̱���u]%-��i���1�F�@a�!�KN�сD�Ƴ!����ᯚIk��[<P�Jߣ��.������|��V���R�΀ȝX���:c��*�@����U`���gIf�5a���s�݉"K�6l�A�Z���`)C���J�+��'q�!�B�f$�!�D�S���AH��z�/� S��&AĆ;�i)&Ж快�L\#W4� �2#��ɬJ�"�qۺ:a��xʵOhu��_�yݶ!Kӝ�Ƕ몱��ܚ�ݺ����ϛd�����D�X^B���<���r=X�p� m��GZ�̒�u8	��c�ţ����!9o���k��!�]RQ�����eE�!�#�(!�)����f���pV��{�������H�F��C�b��6\X7�\���1���dϠ��}0$�߮���(vc�=I%���Y�����!�P?�|��N-@֙�q~�[���LBS1��s�Y��jA�<���Rƀt������dx���R��??U::�w�X�����j=K̭��_ǎ�Xg����B��?�"�`5�;1�y⇹�TZ�B�d5H�ҭ��
�}1}��I����^|�� oή�N4�����R�04��u�t�V�S=]��F�;�������F�H��F��A|L�-i�1�O�HX��Y�l�����$�K���"��[�x�)S�$�Z�?>_�Ԇ�1^P�u��''�S�K;>B�Ļ�b��^�g���_t��z�Z{�g��	;�"��l/ڹ���Nf�SsL�����DeNcYӣ?/PYCD�߸���N�Bф�	�E{����:H��%���#�z��J��dϽ��YMg��; �)[d�2�4	m��n�(!�VX8)s%��0
1�C%�եhpr����w̤�?�r40]zR��z���n�Ԙ���RY�o�������@�ꍤ���>�ԨN��y�B]�WJR�NW�I�٣�k�ЛM���,�j�*@0�S`��a�G���ќ�)W�}ir�06��i����)���&�L���%/������`�, t�-��-Ǉ�q�������)&bWԫ ��7'�a�/��[��HQe�Q�G	C</��#��R�h�]�]��T�-��!���y?7���J(}�ߘ�hK)��/o�?�4�{;��K�Oj6����﷣���F4?�{��j�z����I5.ptq�ps(�?"�w8���9ЀUPl�'O� �<0왟驷��1��5'�E����!���?���{��-\VٝL<��9YG�mVdc�l>;���L�(&>H���]���#�#�mڥcq��(-�B�����Duw��qĆ�l���	9�)�l�#��ol�S��=!O�eLk��
X7����V��n}U9����� ���?P���A����n	g�	V@1=Y��4	?����XT]��++�@�<�CR�~���Xe]$�9�kr�o�|�#ٿ�CԞ��=��X��Ѧ�B�*v�����fd�7�#�uNTn�@|�"L�h?'����{X�N1 �8����"2
������ڏeDmʍ~� ��Au��nZe����5)_h�f��L���ͤ?C�0�3��P��M� m�� �<�GS���������a����{�����y^Qv�v��r��<v�ĥ.�{�+�{�φ�z�fh ��[a�����*��u.�쬦l���92���m��ӊ���yL�*Xг�����E�L��9]a�̖�!��Nz=���;v�b��p�� ʝQYGeӷ�����m����Ch2_B.�r{[���lt�R���t�ؾ���+��!	�$���h�G�d�ej��oy��R#̞`<||Rƣ�T��\FZ����Ȫ�~�Z�q}��^'nK�����Ki���2�ab�>�9dА���m�Ǡ�a��d�%)�v��@��7�wn��;�L%���(�C�N��EIl<�ك�B\���0F�j[@��˖.��{��{!Coya6
�?Y��o���ճ^��|k/�p��7]����;_,���}/��joF�u���e`u�e�d1�}�N{۲��RAAP����p��ƿzI3I�^��e1�jxd��{�F�F�6,&+����m��L��?����qL*ł��2�� G�2=�@��H#H�5�������F����Px�7"�s�UD�Lӽ��Z~p?�Cpb�]R̦_��TĞ���"�ؘ39���ޝ?,�h�x��mP\�(Z�M;*P����j��*������X���%�s1��r�7MU��WD�A��pص�L���t����	5�2� �ԥ<�v��ݩ���@��%��l%��c��}������	�^6�y��K#�g�Sq�:�nR������(ڷ��A����R^�crb�*��ʛ�3L�U�{å_-}�/�"�����ix{ϖ����]]���wB�H!�^E�Z�����a+<s^�ފg�B>�/������W#~�٧wy���uO-RE�M!Ћ�e�]3��]��e�p�� N���	�����~�i���"�u�n���(��Y��xZ�s�6B,���:�B�Hu�x��儦�#b�<�+��%���RT�I�+�/_���+@� �ε7���'7+�K�˳$O�r�T�v_QP�,�3���>�Mj��C�a�N�}����h&��żU�"�c浧����w���]���̻W�����d	������"7��\�Ɗ�io�c��|�4� ���	�f��%N��tw���{̌��|Sp'�m��Ml0���d�,4p�r�؍���H��J��J@}mL^b�c��Aބ�&��j���cë�M�/f�P'~�h�}��6y�PY���yn�����\d$��I9�^��
ﻕ۹��I����1Q���e4{�Gr�ڍ�1��bf�.�$���y؃5=������Խz�;��<.=U�X[O����܎��ې�1>�dLKpV�.�����1ږ���ZԀ~��`��R#�'�/�G �<�*xR��v�?a�=LK�<����5��9"ǹ��O�f��)|2֧}I��B�`t�A1W��-�,��*�eG�����&���Y���Ov�xoYk�=����
���� �E7��"$�ǫ���
�����zB�.[d4p?��/}�{b�w-޴?�a��ƕ;�%�ը�4	⹐�D�+-]�횭��]S

�RT:N5LM�fݟ�I�Ų�LYb����"�B�e�Ɨ�X�;.�i���!�8���1��� �;�,g��s{��U�`Y�DϨB6��L��܎�*<���t�CB� ��Gg�?��ξ�a�7�:�HD9��˼��d�1\(�\��҉1צϜ}��Tl�8p�r���
���ŗԓ����}�Uq�"$��L�W;V3��\�d�(��:bܫ��ƬC�ă�7OQ�bgz|:��YT�[��]~.%��u�]�P ��yQ��ىD	Ca�j���"($�'�p'�Q�M��4{�S��Ue�iBQ�.g_�������T����Ͻ���tM�7����xI�h
�i�Y���s�E��p�j��0(�΀�7��
���Ӽ�o�OG�f+�W����`�(!DQ4�]��#��4;'���a���R�����1y��W;��0K-������(E*~���La�I���bӹѸ[��<(��Ϸ�R���cب1(ϐ��Ś��N�u�c&%v>�Y��.�y0�]C��x�cKS}(8{'�A���h���7�/%1��
p�ڡ��pK:		WK�@�pʦ�h����p*���;�6K ���{}L�-Z���/��6p���;]����{����Γ`�7B��p��_�md~s$�\=�(k�"9�לA���
T������BQ	�u*�kp���/=���A��̰<ݓb�W�&p�j&Kj���A����;��E��i�8��{�~; ����F'��I��Ⓧ��*���,�C��wfh�kT'"<��3�n���w���Z. ��i���'��&�g�1s���Lg�^z��b�V��.4s8g�(���<�HW��E�����ͥ-?�%�a�^�oM's�)P��n0��Sl��{x)��i�{`;��'�Ό��8Z�X|8�k��"}���-} �ͼ[=l���V���f�-_����̍�����/�����)�C6�@��}Ĭ�vS�3k�I5�Ί�F�s~��m�?��C�ɨ��ػ�|g��*���uJ���(?��:���g	
PJ���\@M!�hz���u��/�Ob�1 G�
�ɴ��Y4�ͅB��g�c�3H)�)@��Dg�a�W8~����{2>�/tT�#.R��$�_э� -�v��w�(-��x�4�w4X*�fyU�H��Y��k�YO֝"+��J��sՍ��Y'�<n����W������'�0���>P���U��}��8�n�T�{��2���ݾx�S1��@���7�W�=�D�.7ؕb'e��0�#���㙶;y�(Q��_lۼ��q����L��
�Q�w�ΌG�9�Te�u��)� ��el�K4��� zo.��d����|�A�H]�][jY��bP%Hv��G~�E�ǻ����a�0S}�H���nƜƑoqĝ�3!��6`;���l�Ă�����wiv���S�,��~D�@j�v8�_����`�D����2�&��ڼ��z~�X�o�z�l��8��!���B�&�W�&	�LFK���6�����.2��ЂƭXH�Y��ޓp��se�R�s��5�&���<�9,��:�;No�6n% ��rc��֔�|RQc�[���l �d�?��/y����_D���i�5�<L�.F����=�4��/�8�����"&L1�i���3RZAF�ꖈ�A��n�m�]ѽ�4�hV�-P�2\�G
��bi�n�|�;�t���ݳ�kr��x}��rm��(��W���
�3�ǀ�,eprXz�?�Gl���8�B+&lzfR�
�=f���<��
�`�^ħL{��nY�s����os���=
��~}�M����T�\p5���	�/��at��JxlZD�!�K�[�ɑsy+�5�<���`L���X�H�5�Z��|�V��F�{���Y�N�]I�F�ǡ
�U��L���W�}Ǳ���Mdq�]�o�Ձ%*�
�C�H�V��7�Sy>��꿥�I�A~�+��j�����p���Nc�hN�
�H�hC�Vo ��S�+�I�Uz���Ұ��u[�����af���{�nr^j��&��$�j�xf�{������@��Ai6���g{�l5B�E�ܮAg��XT'��4J%�YX�BZ5+;J}�7�X%��q�Ňn�A�^�Yk���^�*�>���>A�`	2L ��l���ZQ�ʕe��k�,f����l��[]����)!o�86�;��s	p�+p?�c�DQ �e��y6
��,��������w� )+��ۃ��nu��q6/&�>�G�绂���*K�G'�>�r���px`bI*�������1��:C���#m$���iŨ�}�m�m�������P�ߵ����*��Xt��	)��k�E�!�K�g����]2�hU�)�La�)�`�P�=?�gh�5e�jX ��!��lQ�]9e���`r�a��)�Ak�D㖠8����oY!\)XH�$�����S��N�C�8�F����Ҿ���8��;T�	SŹW������!}4��pkSf�_�GCY^�k��ĥ��#�7$F�	���54�EuT�ܽ���$M�VHb�K�N�6dW=&�즨N��m��N��6ٙ��p,� � ^�C�,S+Q�H��)�dK�f��w��} �i������=ᜱ_~-ٟv��}�W-��Eۤ�D9@�Xr_X}ZW�������΀�y�E2̓��Ely�㯃�R�%�y5��/�Ɯ�VI�=$#�����r�L�뀾�{�^f�Vn`�2}jMK��n�v��=��]E����z'��x�$|�E	��8(QB���h���-��+�R"1������T��.1��g��C��'�P|�ˀ�?[
ăRF�U��s�:~���<v���D���c��	�͆$�c�ME"-i��Ӑ��ƍ9;sҋ�#/��u�g"�V(�g�C�g�#�S���|�O�}�17A��!���u!�n�nk'�r���F�
u��~c����)�>LU�,=��#�=Ն02
�� �?�Ri�wo@�Ӥ�I[Udi�x�t`U꙳�=M �۟=��Y��<'� �=(�(�p�Ё	onm��H�'�'�v��f$�͓�� N���6�cʧZ6��Ȍ��vd���6+������0I^�x%խn����m)���L�S���/�t���b��_E��!��]3��QMZ�r;����3(�f	����Q_�ܭZ�m��姛0h����y���xl�c6δ��e5E���	>�s{���P�L��F�����n}�˖��Bv�
j&f�a�a/@�{�IÔ~/6�%z��&�!E�s5T�Ҳ
=�Y��J܋��5�*Y�X�1XQj!�#:�0z چ�(�o�"�èS[��y]�u�|������7�Э�l��X��~) ���������O�Huw �h���d�q�"�/gqto��s��*���f���Z#]�?U6�JD�O��-�	��U�c!k���Qk�5�H�f<A��i.�� !�_|�:G�fG� �1�P\��zgS��^���n7}�-a��!+����4.|�^p;�������+��+Y��c����� �,ς���b���0����#��˚��G,@�:�e��1�8��h� ��Ap�k����4{0�Rv���L�M���Ni���?a?݆�����8~fǝ�Q�a�����sU9v��������qSx��ot�T��|Í
��~�qM�����XU
[a�cp��D��j���f����5ʗ@���F 3�x#H�=H֐iO_Pu�k�[XXJo`�� �"����#�q�*��І�	c��HH�/@�콎㏃kl! ����3!fc-;�IS���!l�+�XI�g����ʧCU������ va<�n�n�zq�C�E""stQ"��&����!�5���{7�N�^�9��OT�0Έ�.$߹eOV�Ĵ&9���p���bQd�#�T������r��)jMH�b�����SIZ��}JCh��fpӽ�PG{��}�Uߨ�>�Kf
�_�~f��Nz�1�˚^���D�[���s�6��Pc��KF���,?::�s3�(�,��*�S*k�/����܎��k�˭	:q��&�����J^>�x�'�$�����x���v��zհR��y�zJ����P��RƻrZK��>/�h�pSq�-���!9�u[�\��|�u�}�u��:�Vɜ�i����߁k�"z/ݪR{�nXn�y�hI�����u%oU���4�#�3`��L��aJ�$.wۈk[�y�3�����Κ�놷)�L��
����޴G�0Զ3��a�~ͷ/�B6rvr��u|yn���cF�8�{6�h��e8��/#*ҍ�.�+`���@s�*��@W1���-/H����e1�$%8F��1P@ꨄ�}���:
�a��3���p���T1���Y�C�Ot�a(��s9�o���e=p���h��XEEz5[0o1b �J~��������H�;�Rܪ�#wUq$-�U����;1�|��3��ԵZ
�њ���3!���v�T��Z_j�HPb�^T�BwG����UA�H��cs��S�{�8�� �Y��[!��{�� �0�:K.Ay���/�QbA�y?�l��G����J�~��zP����q����5�3N�T�l:+q'��R�\,g�PK�[�7db��&�);j]���Ϻ4��`7�ŊP/�t軓�vI˭� �c�{g���DRn]сRx���خ��~e)������Pޅ�5��s �=)���y���pR;3=�s`Vj���5��#���#~lӁ?6�0���t��f�4Sx��:���Ⱥ�F�_B�/C���}���Q�b��	�i/�5;���6.Ϡ>	���X9��j�R5 Μ��.k�!(���ЕB��.�F�Q�2�<�fx0����fi�s�t8W����{�"��|���&^��=��	��Kj���1�W���2����\B(L�h?��B4ݵ)��o=��`�� �4_c�3l������<��wj��jP�6[�hO6�!���V�k��Զ���Ϧu��*>����~U��/g��Pܫ ��U�%B {�N�7%Fr�N�)�٥�ug�\��V��%�����w��r��!:����Bu�����5����<`X�|�-����8���׫¶VWE9p�F�7�kn�Qq��|���8*Q�Z�D�^I�fQV?S���k�[E`�V��8�� ub�v�a���Y�y>s�{M�����)`��-���ͩ��N�!t�_��c��-az�f�Cty�~2��tЄ��;H�h���lf�}��zk-��m������*�W/�_���N��~�D��W%����ےG[��XftO�.En{,s}
��y.d%��*��69L��|���QA��N:y8��D�O�y�(������mY�7����Ӫg��[I[1�|q�6m�	��/�3�Ge�,ںʜ_�֨��#�ndK�@}��P�a��m�d��%��E�+}�޴ܔ0����W.h�Ч��6�~��z`��NLt�����x]�}�m�q�h.�
�P.�)հ�+�fbVȾ�����_ϗ퍠<ov)�O�2B5�}���ds�`v̔th5��_�I�֢������	�_�h�Ei�6�� ����W,��Q������G+WA�ۆ�-k
�|���>�R�|���l#|=R59��,�sv�2���	kC�m)<A��V��"e�|aE��[P�Q>�X�c�P`�Ɇ��!:�أ�FUߙ��a8�_1g�#�P�j��<*$�}�M�l���#P(jO�N`�z�8,��������DL��R�-�RF�z���p9�߭^�h��-+����- �ry���mM�gYR';��P�OY�Z��׸��	!=J�����8�ݠxʁ��G<u �EEb�`Z�h�e�l X3&6H�8�&��N|�ի�kb�M�!�Φ�r�;�� @��i��Z{�b����c�`�R����^��F�s:��
6Y#����{(�3�P���,o}h��7| �ԅ��gm(^-�Z�����v�z�f�!�(y����r~��%r��	S�����q>��*���M��k�Ż�)�JO�ڢ,��y��*T�C?(e�D�;�?��8 h�aF�j/�6^�[���,/�#,��BM 8؈.4F����@�	��/V\�a[l�]v������޵��wK%�p��������IH��i���A�ѥ�K"��x�a|$\�j�+�W�lo���!X%P���y����˻�-#��![Q��N��
l�u�*̅A��0�z_�}�r�$|�`�K��9�I�B� ��}�A�9�<S�v����Y"}'��z0�TT�%�JyS�Eq�^�d�3�I(W���[cxR%��dcD��Q�R�C'ݿ��zXh8}�:�F�|�/c�y���'���5q(�y�s �F�.���}�M�@d���F�u�HPO���m��S��z��°�� ��X���9��Z�U~*��s�X��}�=��൴'Eik<��,2������9�[�Z��k�jp����4~�wg?�7� 
-!���@�V��� O��7���	J����}#.ZP��;�&�T���Z[���z��rHzj(�R�����6	s�p����S��
�h��8��"H��=����	V2iH�Z�'�>��U�FT�"2�)0�R��~Ss��j�|������q�Z�̎V
f�E��� ��ı��@FU5�V1>B��?�*Xր����d���n��.�E:�QLo��kԘbV���T؏%�ڱ�,���FAEօ����2v����
��������a�KS��J����`�|һ��;�Pz�yq^ƕe�������¢�覨�þY�e��w-Kml������'�1�ۈ�8!�IA$a�ץ؄��L�ɧ+�T 2p�P�q=ޯ�a��Rn	n�bj��٦/p�Y��9��gM�)�C���(U]S����W͑Rs@;��离!�he�4�ZU$��f��3�T�T�i>r�I���AP	�����y���0!&����a�fΖyd䏏1�p�e(��P���F"�:W
���^������G���hbQ�ם����
�hv���c�cN�*G/�h�,j.Xz���c��'�Y�J�P���A
��4��)�k�:�c�K��)��O9�YG�=[�N������v,9�(9\�M�F��QT�~��&��
�
�ݭDh溯�>l��J��[6���öti���; DI����7K���,��/��H��Հ)��L�Ӎ��c&���#�-���q�������_�	0��d�Q��8U�� �)���ڇ��{V�rh�R�!����#�M|輟���P&bJ�.�(�ͬ٠��ћt�.�0��lѫf������8F׮�1���G�O:��V@2^�0T�a����F=kN]������\l�܆@�a��"G�y.S��m����������8��s`� ��QٽdH�7���2��zwF9��*v[�QM�5� ��6p`�k?�'W-�r�1m
����|��s�	���HҒ��4^f��V���R�Y>tx����I���G�N��7�_����(S��)i~\{����7I2���L{b��^�aL\w`����z멪�������*M8xdgW��D�τM��ɳ�$_�eM�,a@�hv���V�$�d��Y�T�s A<�o�|�&�ω�t���*��u����PɅ,�gP���lL0X�)�J��\O�!�r0?�f3�:�g��{�+kx��h���~�?:C�3��'��7����Tu��D�mS� 0���}!����E�o׽��m�:z�q�C�)�|Y	�N�r�(&����G`�l�j�D����A=x�"�N�����R�	��#���ЛDo�Y���˃`��xo/�+c�ru_1��͔^O�M$`���6>(m�O�V�KM�I�kYGtw8��̗��KJH��:h	�����Uj��ӷ���w\��3�0A8�_�@`���X:ywA�f�'�ڴ��e-�l�����M�������0� L;�RL'h�e�7��~l!Y����9M���]��p����h&� �)��)����0��\��-���P�W;�H#Uo�O�8V?�+7�M�����0ɚj�x?q;�Lb5
:��4���%3�"'0A�w�܇�V�d	�1h���S%���)Mʭ�u(ϻ�/h=�H%9�`��ף��#�,e ��7�$�����
$�:�S�y`��|�⼷]Ȩ��zBQ�Er���*A�;� ��FjT��1�:EQ�����Ã�����X~6+@m��_�L~�If�m���\�*�4���R�2IyQD��O�=7�� `yX,��.M&S�.�����rL��"��I�iC��5H:e~�Ef�	8s�����=i�젔�fO	�A�Q3qM3��C��z�����"r@p���6������i��L�3��/�/,��M���~����vʵ���-�Gn"s�>�a���ăk��ul�C�ɒ��	{��H�Z�
�C�G:|K1h�ϫ�{���!�Wi�>�JCf}jz����~�T���3|?o�>]�z�!����7�#x��l�`{�L~%,U�o�?Ts��[oM�s�䰋�O���l��ߊr�h �
�\���P+��$T�����p����
�f�dw��@;�0)Ui@M���g�	���\��������E(i�6�l�O*�ꐊ#�X��NAO�SkWB�+�(��pɪ�t�V�`�R�g:�+	��U�Xa��Z���F�y/��y̶Ƶ�]x�����������ݩN2ˉ� ���!��򕊉�R�U��e$\��m��$&+�kS�.�w�����D�b�I�YҸ�.=#�F��e�s��Ű�^�!�i̤9���@*���vr6�b���E�Q�z(�� ��G�%]!$Z</>���3���o��� cc����C���~�̤��먅� �����o	��2�P��J��I(}ܾ��s?���NЌ�m�>[��0!ǰ°�V�ۧ��m�>�=P��i��kPЗذuE��d4��/Me�O����uӆ>]��Md`�ľ���=5��6r=w*/k�,���� �?F���I�ϣ#i�ת��K�sJ�������k9`ڎlMJ��n$;[i��V\������R�Ŝr�}���	�8YLT���_��
` $�Z�t���O����_k��WvZ�6_��̔�*+�vh�'���˖��k�n�U�љ���������TQ_�{UQ�p���)�}`jU
4 �JYp%�!�j�4DCk���W�m���AM������<]V�*��c������Dgm�H	*�^s��q�����~���=iw�L~��u���M���X��mQ���9�7u����Į��S�j��ܮӞ�}�a�@�y�3\��W�o��Wsj"Qk-����]��A($b!��Z��j;�.S�N�s����:��y���8M:
���x��A�7�9N*-UJ���'�[G�2a�G���2+��'!��w�����6�@�[Gڼ1��k��Ku �4	'�v��f������	�jq��0k�o$��}ؔAz�nājn���,��H?Xg�|	K⾡���+�3��:ڪ���?�g�W���1�����QZ�E�i��^��7|X��^��nlO(I|=����[��|c����� :ɻx�B��Ut^%�+^���Gj�B@o����첩��@q&aZq֡�`�M�@2n���!���**�t&�L�q;�v�o�T?��]�����:Z:��ҥh{ݚ��nw��p���$�r�C*]r�����C�1�ѻ��Lk�L:�YKW�o:�.�O$Y���֥���D\��O��M����A�y���'(�$��r�Ձ�/M�i����_M�Cib���������a\0a�{�z�PEV9���K�W��(-���A @�
������6vɥD���)/�K��Ѳ�D�aQ���� ]�A?fM �����8�#�>��`�A����*Qs�N9�xp������R+j�%�ZF����j���Gi ���;f��C���I��TAh3B<2����c�M�$cP�)������~�k5��?��Q*L�=>j���A�H'b�!����U,�*�:�|��P&����=��{<!����̢4�T1���v�-��B٠��EV��������V����D)+p@�S���@�hJ�w�& sw���)q�Ti�&��mOax��Q�L���TL������W��Cׅ��/?�n�)��a��D��~�ƒُ��-�ч��*�I�v�lz����w.`I��|4�-�!�g�nX�,@���5Сb�3�T$���I��7� #�J\I,����,����rH�%��tq2ȩqϙG[�.{Ù������u��@����g������﨎1��
��_n~{�j|�ǎ��&�>�σ��	�&�e"��$�L9[]&c)'��\�~C71�'I9��$8�e�(lbyw��!/�u��꬙&e��Y�̴���?��L����;|j�Z�0<�oH�u��WL��bNn+���#�y+_@�R���wQ��#�yvm�Hv���K=5cp���A�`�O�d�%Ed���B��$6��q���-g�e1�aB��(�ʡ�a0����-���>���U�q| Cj�KIEV�J�uY���q�QNW|�p�r)��]�NFKkq���u̶Ώߊ���7%���<��74g��|�\��n�K���$�W�Z�5l��3�x����,�G���n��s�5��p)��,���f|�k�A�,��D�'���Mz�0_�p�~��}�@�!�%K&�=Zz�������s�n���{]����M� ��r#�b@J��!�F���lz]tJ��D�i)׌"�����y��:"7������֌7��m����xS�����X�mN�� q!�������3�/}5X*������ϗ��B�B�W瘈�X�`H���+^�g��c~�)F t��u�G�3�c��}y��Eϻ�dq�]uEV�j����e]<P4�b�Ͽ���g��m�a��<�0��c��ԍ�� 8��&�aX��+/��m�fFT�Yz]��zC�}�DN�w��TV~H�ej[� ����N�D��sM�t5�$(c\�|� �F���s2�r�6+F Mč�ud����RU���;XE@����B��Gy��Z��M��Rî���X��e/��\˟���шkj��Y3^nB:I�W�!�߾��ة�<�;��ѿ��^�g�9[���h�B����(���o^����cn�d�'x�#��B��]��lO��D+.^�ՏP*k
®�9@�# �"�B��ܣd[И���dn)VTz��D
�[#OJ�Te�އ~^x�MrY�<,��H�B�`�*�gg�{�y����k"�n���$�X����`5�L�����N��8�����}O�6R~�i��w!v�z*����~�E��h�x�Ի�dT%�tC@�ƺl��`r�^��g���/��#�^ee����ٗ�Jn�L��z<��q��`C�yWm�uf
bq�V����=��� �p
&Jbd�q$@��T��Ҭ��6	{�ɶ P/Kܻ=��!�� "&qe��/�f�X�)�����QȬ�ؖ���?B�e�0z^�7iLHM�v�H����Դ�db-:*x��ni���i=,ۖό��V���1S8�Ŧ
?�+���D2�=�Ѣ7��U�N<V�?m)_�P���v�������+p�*P��e^!3�?P�X�A�c`WW��h}�C��o��+^��VY.�� �\Hך������Á	�� �*B�0b�ΥIQ�=�!Ih<�}%'�Qm=�w��PM�n��nN
j�33�����:9j ��DIS�̅��(���֣�0I~I��Y�j�ԍ:l�f#V>�P�"�:b.������I�E������ø�<���χ�/��b)���ö�K]��Z���هIMCq���qݧy��5'�s�9:��Q��Ơh��7�z!#hS�w��e��D��q6��>&�ё�W��,˿���oO"�
�Tg�a9���\ _}J�Z�>��K�
�
Q�*�Oј�m�`\c�J,�-�s�g1����_��
*�`�ܴj�b"��X� ��'0��wq÷��⭮v��W���`���޽[q�A�[Q�a�.�y%��[�uw1Q�b� �)�x��I��� lذ�ӎ��P颫���UM,+����l��]�Z�IDQڋ�3x�k!1��M���2���r֍�e�Ն�b��)����~X�@gə|)�O��;
�nѓ)Ok\\�g�Ϙ�P�Z,'���|����4^�� �йih�́ϯϸf�;/����K�T��=�j%�E�(�Fi_�l*�c�[�,�pg^Ô�[��daў:�ґ����zR6�J+����pS�Ԟ���{�ڛ��e�ˉ���Z!As{�۩bM����%�s����C��S����)+O���O"���Y�*]��������x��
�=�� sW�j�QU7���"�KE�Sx7iz�W�AM#�ڟ�B���'�K���J�!�-	��<������5l�F��TG��:�'j�	��E����(�j7�d�I�_>���J�0LtO�e*�1P!�ݚ?-D�0+�%�����o;�Ga�Q�\�F&/_��1V���ue�0�	AOs�.�'"N���RZ[�"J;��ӎ�����b`�x�(�DFq��W�\ֈ�jW�[L�&As��`���f'	.�^�$S�a��AFy�v燂�ɵG�'�\`�*��k�|�Y�D����	:wB� �쬚�� �^'�w�Ss'�t~�y�}�����|;o�����.�a|�"E'�!~g6����wo��F�˶ ��`Nz���)�K!��֐h���0^�8XTԵ���aQ�z�^h�/S������t�$O3u�l�$�{9Ψ�El>Na�=�q�H��0j�ȴ���7��I(.!>08q:%CΫ�zB�KN�+�e�#��u]@+pp#����������B�8��,=��>�뻐�C���5���@[��6�=��1Xa�@&�
c!�Pޢ\G�*=��\��<�a)<r_lsf��y68��Oe6,��AI���j��'P9C48�L5���k*��|����S��N�Sp��I��s2^R(n��w�A�&\���Gp�S�l�Wg��'-p���vK����U���U����4Lb%���G�q0�n1�h�?�M�~9��9'A*VXњ°[��`2-[N��!X��(�.$��p��(��5�<×����gk3Kx��no�_��*�YN��K�̸�2j�&��p?��	���a`���\�I�BW�x�d�)G�@�;f���7v��L����,�=l0�O��:��x.�<��RLV2l���x�f�6(.kڪ�!��?�>�ө'd3�nׯ)G�n����j� ������.R��y�}9�GDe=�p֋a�1�X�Uf
�nҽT*j�һN�8�֥N�P�E���C;��?�4�l��9�Mb~��X�>��%a�<5�����&`,N���7��Usj��qt�	>,��f�x�'釻�9� ��[� 1��=y�_Kb#��|y�C#�9f��kv�,�E�!o.p�l�qR�e'�O=t>�6�'�=�;��ʕM�;XQ���~�������-���3v���eָ�nI��aZ-(\[9S\s��=���1h��tOŧMg�Ctc(��q�����P��}���-�ʬu/��nA��T�qi��_kB��v��{��$X��S��b�zg��~�P�$@�����z�0�ˤ���	]�<~ڒv{��/��I[UQ\4o�7��(���[��"z��!�y!Llٕ=߳��_uD���h/o	�u��PT�0,I�"�XY��e���8�ظ�޹�ó#�����oɝ��t����«�L\��t�4IIGA������huz�|�2���������c�G�����I%�����>S2F�T��oӂ���zD���K��G0	�G�����c<������������}��>�nIe+e��o9�(Q_�K�׿���]�F{[Z��p�4���1�6�n�Ub�/l;������g�֗�����k?�&�&���8) ���o�F�Y�.A�4Z:o3_�L��zw�����9L�ɻ�WM���L,+�Y�)4An��娋�ܡd'�K�=�䚈��@�ǎhl� dbqE���	^��ܤ�Y�W�%���ݬ#=��`�y��ڮK����q��q�fM�""E�7lUh�ir�B�M&�q���a�[��H)e<B;!P��Y%���y�+���$k��M��C
�3�'�̾�!�P+<���lX�v@����4!�w1?&�\y]�u$}a�<��z���i�F�Ajf���S���9�;N��e�8�~I�cgI�Oj���'�
�#t�&}^�?��04`-�O�v���&ɝj���OU�)���\gQV1W�U:_��X����н��T�^�"�ܢ�ɮH����db�8�}
a�A��wP�Cs��Y|�G��|M�8P��K����R���qw�����x!#
7Y��]�6N��GyXB�úR7�k׭ߟmqv֕T��p@*|��c������G�<K?ȍm����<{���$i��s��\��Vq���4&�>G���k�0`�w����*����h��W���"Kà
(fѡ�DͿt�h�� SQ��t@_���xE�hI����a^��/�1��T�%ju���5W��B�t$ף�I�X���t7l
6�^f_�UV6������~�e���T��&�Bph��C��Uw�x:���J\B�o�pb�c�}�?�MM��
�%� .��'v�5���:}��4N�t�T�r7�u~O���g�ߌrŋn�al�!��!�\�!ϥ���Љ�sOM̺���?pC�T~��vs����±tA���-!����lͺ-L���}�K =�_������s|�8��re(�t�	c���OL��Ŵ�t���L�v�}�DKĂx>ԟމ����UiN�<�&��[B�N��ĺ���I�PS"G�<��~���s�#���e��}���&t��I�q(���)�NP�Ƿ�h$�R9���N�x�����R�. G��I�^�қr�֢���ίo4/��[6P�� �u�^A�[l���8�!���B�ܵ�JE�̀t�fx�W�5��LY����_��0
Gď_�Γ��=XF�~��N��*��o��?1��\�.zy��G�#FѦ�Wd���T�󜘧s��W\����t��+>�(l}3����R_G�A���*̕dtd��Cl-�֙�Ƹȧ�2�{S����j��պ�D���i(&���S��aMޥ�!�'�D�RPl+��'���)|�f�X���#8]VAr=.kx��%}��A������[�}ۼC���Z�����!
��+8u���������o���%�!e�bRL��A�w���n��_��5��Tπ��TW�M��m?/b�T�Y�����z���L)�)K�xn SBN���G��3��ۯ+������������q�q��d(Z�������>���Md�ξ,4�?} ��`r�
[����`}G��,��m��?¸+��V��,��AfL1?���)lw�e�����7����Q�\zCc��T'ID����+r��ʪ�P�}am�QGt��5�G0[����(}�A�;�y��p��f��E���Lg��#�8�#�΢����c�3���E9Ll�L�{��L���"��p�?a�F;�����v���9<�<P��{����d�T�|���n�]@�7\��7텴S4
G��A*.��M'�����������1b�)��]9�Cy!�������((�)�`�Uqxg�|�@>�M)E# �B�ӈ�!]�}ҎS�{��.�:��׻|/��z�ཬC�z�q���~� �~���[�3&L,�\������n]��e*L�Vwv��]��:j�aԒ�䞋��+�\x�R���ge�ݚ��z�Bv�3��O���~��fG���o�%bB�Lg9ۤ9����ܨ%��3|1�C?*T�r�Lj�V7	)�H�/�-7K�M�R'��7�l_����F���>�Ӛi/M��Ѫ�%*��aG�)�έ�6������hR�����*-������1�3���]��$�L!G0�iKZ�F��@�E��z�G1;�ىа=�~!��S���x���. (!��$ݨ>� �<���@��]�3}��/D��&婙�3_G��CDO|�Zx��y-�3M�\/	�>��C��p#�@$���f'ebR�X<����B��!��cALq�0�4{n"Jh%��r�#�ŕ:�"҆-8��ǁ�� ��}���F(�.���U� �.B9���9�������z��W�:8�֏���ǆ��Ik��!�=���y��&'�����দ����}r�m�MY;8j�![�,�p=F}~�=_�B�]g��F[P�Q`pI�|SD-&�����SX̰��:���?�ӳj�?��C�u��߭���S��0�X���=ᐫ�NC���9��͗��K`5M�틗�u��S����<k���'D��t����`M�N��d<������O%+��MU��e��?B!Sb�
c�W#�D��`�e[T�=OН�q���8c>������B�5�P�Jʷ��=��h:�!���f�ѢO�upv�������E>��g�_XD�2��P)}k,0����xMc������*TN,N��H�Y"h7�9�Oa*.��0xI���>��;����
�6�DױcZ;-_&4�B](4x/)�Y�"rkR����J[%���{��_�v�4s/Z�0~4k��ռ�n��v�	-���߸�넣9竖u�E@g:$�}	�~��ԗ,�x7a��EW'����������h�h�-�>��)�#]��F�{�V_��ei! a0�z�B�⛕p���h�y"hSop���o�l��⦪:���*��Z^
� F��@�)��ʳ�/R����#l|���œ�Mxw]��%���B�!S�H���LV֪���Qw|���rr�.��|>�����D5�:��(i���I��ݖ3鋅)�9��۪^p����}���o�)M4�}�rH�l3��5$���E��_mH�qA83����� C���:��Y����	�o�ʩ��
O�-����m�!�n�\9���$Od5���S�{��
��/Ayq��	��6N����2��姆DK�%Nu������$�-�٨�F�kEۘ@	���;��L�����=W&A���1!iS��F������}N{��ԍgi�dyZ'��m���N��~�*��NVX��{ŉ)�|~��7�";~p��H�5��KdʛK�R=�S��Ԓ�Ί��n��o��m.�pȔ;��1x���������H��8⒍]�%�2�tf���P�ʬ߰N$k�]:�'se�{�L�G�w�<���J8�vT���!6�^��&���rg~3T���w�d�ܬ���ז������|�U�2,��Э\��c��{������&D.��"p���~I*u*6-<C���(��Z5I�V�Fܺ#1�XLؚ��ۑv��w/�F;j�6piS�B�ٕ0�*�P;���!�5��?�^\P+9B-�6bU*z��\� �xqS�RΙ����WĹ!�35�-�y�롈�R�>��H?{c�{#�;D�1���dgvp�"&ğ�T�y�LB̓��ˣ�V�<?SM��4�b!�6;�8&�%J:��H�n	i[��?����F�����I���_�S5��L]ի�{���B$�QR[�-�u����V:ӹ ?���YxP�N��=��7��)��9�a�W�"nˑQ���d���_�v�+��y�7WI��#m����[is��M^���	a��z�|�7z�q\O�T%��M��K�
�B��S~��e�7<�����������Ώ�P��+���b�H�-?8�!}M�* Å�6�Zɭ�;�l�$�)�ޚ�Zs�h����HS3��KPdZO	t�d�ҿ��F�c,G�tċN_Q�A�7r�]I�c[����1��?�=�󁗄�V>
��]��x��r!H�I>�q��]h�)8\����C�8d+]���k�˓��;�$I�X�_�Y��t�ؿ�^�:�߅@t0���X�t���]1��J��=�\�hxh�@p߀�;,s��ĿX�0�������t5�;n��8k53�i�	�gz�r*��
/Rg ��Xd6�w͕��E"(�5�Y��]>7���Χ�Or|A<*�#U=&x"�4% 4Ny�k^��s�ĵǫ�Z�r� N;5�3�b���%�v�´�c5IxlB\%�B���0�B�;��P����s�G�䁾Ft�'7��xW|G*��+��y��.�ػA�vR8����q0�t"�sC�j�ʶ���܈��ц�i�<#&�b��,)�RXQ�Q������*�fn+y$
�#���K��'Y��OHЌ����U�ݤ��"�Ƞ���Fj&���|��W?��'R53��yNV֟�\g.���-�^�غ�<��ú0@QOIi=P�+�ށ���{(���@��zģ��`5�J�2d����C������H�M��}�a,����tv:�j�؝~���ve��y�pCyy��%����D��ĩI�n����WC�����͢�<��C�Ya|�Ck�������$C�W�Z����M.pt�+�l��vC�ؾ�8���6�I�T�{�Vp�>�Gx�c#p�$=�X�����`R���R<�w>�+<�<ziVP%S�FU	e�����.d��uZ�G�v�$=�E�\�t&Q�=
7����
Jo5eT��O�7�>ŜA[��UnіN;�5{q�l�x6�P>�'���&�C3��a1TZݏ��nG7_;Gx�؎��mi���E�FʉJ�BƗ��LY�����d5�0?ժ�w��X���Q���^�x2bohA��#AC\��pm���3�Ry�AjoxR���O�+�ߘ��^�~yàڔgK�\kS��BH5����ѓ(�"+���Z}�Yc���մ9�ؽL��
�}G�,=Q��u\�D�������r6M�2�<D��Y$H�|�B�F/(rͦ2<+�O�5���H��?ap��߮�8iDLϕ��gC�C0)'���A2'J��~��h]8��&����t�<��6����@��x��ݲ�.(z݌"�JF��f���[F��UUY���ܥ�m�F��Fu���Ȧ��%K��z"�֭_�����j��>|{�(L��KUa��nl4��9��|� �h��L�v��__Qג�&XQ~FH[|�;
0�zvRp��!o�J�Glw8�Cl�lQ�*'>��d�~{3����`f�:�ټ�a��M�����m&>��ux�,.�D�N�ȊD�94�u��`��h����'c��E=@��_C
{�+7r���H��K)~.��'�E��(c�ُ��1�$d��ͰH�!_���^�
��T+|Q3�-���X�O�3'�����8��;�k�I2;No�^�avG	MfA*���̝���5& ƹ�A��F�Hc��*磸�Vm��rXQ7���;8)+�T�Dp���h��-H�f�dA��3�؄�V�r��]�ֲ�3��[��*<�LT�� _�J�A�4���Lؐ/Dno�������A�����J�#�#G�D��{���R� �y�6��i����YH{ V�����}�<�/g��
]���_�A �*��g�	�dN���*C8��9'����dR/۳�*�l���cR��-��\�.O��>np/�=�!z3�1950��qXΜo��9�kZ(�]t�!'�l�憔�y��'����)��p�5�h2��等�:)��~-q�#�Ș֓&lqCJOߚ�>8�NJ��?��|f坾��MWD��|�:���@�ᆟ�ּ�\�E���c�gkp��Sx_�eZ*^H9��k"��瘽	@��9���^w;�K���z�>I�E^p�V� 4�D���/�8Mf���H[���ϻ���pW�p����#DWtNfY���EuM<�g�?:����S��RO�K�I�s�����Y.�<������6B�����\x�˰�m�� =����Q}����/v"_Xȿ�2����Y��7�(?���Eby��CPW䐳�P�Ј!�-��3T��)�yi��
,�Θ�.��}y��>v}�)vV�$0uD��x0h�SÄ�`�sd>,�:�A�77�c�$P���ŢN_)�������m�F��}�'�S�tW<�LV#�k7�n�\&�9�W�/����֩J��Ȓ4�
	���4�q�z���KA#�"�i9���Y��L)'��������Y&��"��j�i_�K�״�NQ�z{�tA37
�}��p���Սݕn~g��/����1X�~�u#� �R����	�nJ�E9]�Tw��H��-H�s-T���{�_�Ef����6�:�`���&�hݚ8�r�5��<p��/����B_�y7�.��� _�0��Q��	���z�XoN��#3��zC�n-t�� �,�j�g��Ǚ���HB�c!{�Y���=_�͇�f͠w%��F�//v��_��.��d����8����J��H�`r|�Ui1k*�)�|a&�յ2®� n�?�ׁ��Y��2Q@E������O&[��o��N��4_H�����qa0[�L`OD��t{ò��F��Ѷy9b���O�����Sf�)��1޾�X@�/f�jJ�2�A}f<���sr�CXN�O,�p��>8��|K��}}�e�e+^���ɹ�I�
zI�K��w��.��|$<��!�?�������tw��І5;��l�d[?��wk/�8j�[m����i�kۣ�����\�gD-���q_��]�6[JMǤ�hF�š4���]�ٲ8%��|�=O�Ũ��i��sq�ͭ�YZHb�x���:���& ����v�-_�L�h����!��z&,-�b:l��-Գ�����hK���p�,Nq���3�ii�!�����c�ѯ���>"��t��5��{]j�,�h���	�X���B��$_ԤI��NZ2���ƍe���Iz3ŕ��C�.BT�
0)xi�������cf~�����Z.h�r����l�;2�6��4�N
�2P��G��Wb&A��nH�I:3��3�X�֋��cYF���ˉ��������t0���^�, Y̰���G�����}�fTF�ǐ�5�H�H�?���js�sI.��r���e8�:�K>B��J�����V�q���{�ov�\��pEћ��á�G��!I�	N������T��ֵ��$�˄�΅�bQ�;��f�3�b� rrf��=�_�j���.���"Y��!���G�G�i�{���Ӄ[�E��C"��[�b8K�JN ;gE,%���daGڿI|f&�)Z={$�0���7���J����i�\����wM����L�?D�N�����nO�n�X�2.,�ϙB���c@�m��$&���q9��n,�N�b�?b�����w�u�|�]%�q�>{�S�i0�� ��XssI���6Fޓr5!�#�gLg-���$�v�ض��A���'˼o��k��'����7Y\��F8�3���rf�FJ��p��q����ķ������3x�AT�.ayI�w^mI�����dS�c�r��."�������;�r���h#iH����_l�%@�V����9D�8��ea�:~��'9�?�3)hH�Yy�����2K�p�4C������5�|E׉&1t�y���\B7T*%�.+��!*eR�3�z+������3��{�/�X7���p��"�ǂ����ĳ����#(R�b�E:B�0t2<[��\�ґua�k"�/7w���H�;\�U�Qy��$�;�o?����]�ˣ���B�?Kx#���E{�kK��
ǫ��[�|�����遺}�#�u��ӓT��*J;�09��y����ċ��ݦ�(���	��ܻ�������[=޿u3�b�?�Otš�.F���
bO8'��H;ȥ���6vM�m���E��_�|��z��B����* �`r�����mcè>�wR�g�8m�A�!#8?p',#�W� !�PP�CȂ7�51h��}�Xg3�����2"��d�0�����5��q�l����s*�=�J���W�x`VcI��`����a5+�g��Ȳ�s=>���������e� ����aÞ�Y��	u�������-M��Fw���ƶ-r�4�i��lF$������l� �"UE��3ײ�w��γ7�x�g�j�W��]TM�S���r��&�lv]����n(AE8ϲ���?'"�B�m��9�*m �M���"�;1ht�+��zx9�O��V_@���{��zGN?]��A�g.�n�]F��ƌ�?
��������1"�|FZo�0"��k�;�:Rc��X2+CU63�1_ʳ�
 ���M�v�g��%�h����2΍�a.��˲%b�|�˙ث��8�̃i*{}�wF|�u�mI���U����������"t7��'B>n�#���4����a=dVHV�cU���k_�ݍt�
`�w~��-�q+��
�ɒ�Y��Rb�$�)���S�ZE�����ln�Y�h
�wbj��GM��*���H�%=���q�*9��u�VO�L.�=���<��I�z�J� ��)�^.@z�jl۪HI8��{i�R?������=�4��j�z�F��e��+�d̂�Y��:/�} P��ɍ�@������m���#,����^/|�_&D� ��8�\t�9�Y?iӈ�{��
;�*<�֟%�	�U���H�m
|���A	��c�F�v?w�&��Vq
���j���4�����o��Sp�0(6ʨ=V+&~
W�vP-\j��"0�+���ꈺ�^`S �'�z�֧8�ڕsU-1
��c�I+��Fꀒz��՞ RG	2���3*�0H\�]�<4,�.`E�{�o���}�vn���
��1��������,�Ғ�����7�p�(�D�gݍU��!�\:��oQ�{D���|a,3Ӽ�c�MibƜ����T_��9��H�:�*}E��&�������7,���T�|��^�R�d��_�ا�G���/������;)�����QN��G	�8a����I���XӬ�G��c5�+^z
��ʊ7�� ��U����b��PP㿿���Uh�ɼ+��+�3��}� ���U��W}�~�	)�ȁ�>��054x���Y��W{�IB�c٩�<ԪA��x>���;�k�B�z7�H���R�9=1�$�ⓕ[�J�i�����.-�������S�EN�������pCd�/A
՜ӈ��
��<]Ԩ��|�S�1��Ț%��1�J�B^1Np�
H��D�� 8<���V'w;o��"��@���.�k��I�����D�����ӟ�� ��=�Htp����o� K�rJ��dλ�֛t�c�#�	m�d�Ɩ[��u�I1�~�iQY��U�T�ixۯ��u�aE����M}��I˭a��Z�js��`��}� �>�5v:�Id���3G`2z�D�&�z�`!kt�R��d�r�^���:�Y�sC��o#nt/8��U�/P�-��@�~C��?pǲ�*��o������f���Wz���1O�댑�#K�?5���'�YWzV�ѧ�-�k |��
�Y�4'����k{�l��8�`z���Jh��(�$���~Ä)(�xw'�vg���d
�9k��.��*�����j�&q8稰y!c�Մ�x$��v���m�I�ШNS�(|n�s�eP
�U���2o��B���O� _���	x��(Q��?���؈MbWX�|ϩy�xdN0������>��;w��UV,1�q�ۋ>���:0���s�4�Wy�#Bp�Y�&�֩"���F�qL�3���A�G�d)�!���y��zC��Vy¢��`�J�Q<��^��K���ӑ�2��@Nj�t�:*�^�W@|��:��*�g�H	�8?N���%R�n��d�D�q5��;�g�!_g�h5mg���ڋB�b;���+���P/���5HG�<��5D���ͽ[{#$�l2�H�W��ǩ"w�c�o�Ǝ�"�A���Z�V���$i�:���٧�������0�_��4+}�x�a8;�z"�v��F�rl��G
��R����������(�;��~x�'�3� �m����UL��V�� �Ro?a��ws��e����`]c��7�M�>����ê���}����%.B�|��`et=��a���F�q��*d��T?����{�}0樂p����y�XFI�lr[[��07T�JeX��'lH�xf�2:�ޮAAQ�%$�d;r��\�����Y�mhMrװi�]� �'��B���v�PK}��>�v�},U���UC��r���^\˰Í�[�f�ye�r{��{MA���g��M�w���R�:Ɏכv+al��Tnڰ�"8{���c��}�8�hP\�9n�0E���c�Ǟ�>�
*ߵ��#r�����=�r^%��[hY�#�ǳ�H6c�:{#�M��}��a�=�
���ƣ�Z����CzU�����tHmB�|*fk[0OGi�G����9ᴊ��xK����{�I���$�AבdE��XX�=�C���YF^�}�R��4+����w�6�=���L��Y�#�5x_�������	�zZ�c�	q w��p8�j��n��{ �Ԯjދ׍%���e��P�2��vZh�*'Tb�{� [(U;�=<�!ى?C"�c�6�S�=^$|*�z���`���/��[�)� ����1*�����2����8m��\���Z������gJSa)I�0&�A���J�H�������u%k�~�>F߅A��\�-h��?��Vz����֭�b�Ò� � ��U���dPĐ~����d{>�3G�w��Zo��v�sSN�N��>
�l��5$�X��8���L8��R���!�/ea4C��L��*k�uS��6L0���k����������" �����^\�����egV1AO���aSd�� W��n�-��Q"But|l�)
")����-w*1{�lN���-+���*^g��N����u���؋*RI�S��(�Fm���~��fid��"��k�q'����_\�h�Ӏ�X\�g83�oC��>R�y�����'}�OIq��{Ba���axC��~��'Sa�O�F��{�H8ԓh�0� ե��m!R�O�w����jV�w�D�����I�]�*AdHe�/�T�Q O��R��_��1��k����+%��79��R�4[�ɹDS�������:�k9G����������sk+%mWdO���\��ﲈ�˶�k���x����MVw���UQN�)�dE>�����H�N������ݔ@���==`�D �L���NI)��
L�2�N���Җ�ꏭbei5���v��i�O�8d�7�ͧ>�
��^�}/%��Ђ`F�Y������]���Y�\�oYi!n������F9��yXYفרUb�,.�0��<��'D����%e����I������d�$C2�q 2%N�ṙ������~G4��3K0)y���M�&|D?�!j��πEvq
�|L`�v���|@��4�ߤ1���j����` m�/8� ��s�����hs�~;zk?���}�G��Q��N2肈C��C��/*<� ��(�>�s�Գ���h���ӏ!O"B*t![�jɑ��𞌍~�Q�zQ���]�0�I��d	���p�h]��Ԃ�)��V�!��5�������*��5b��!OBL1�T����M&�}�Fď����,�g���O xÓ�@��qt��-�#�^���o�`�Q�m5l���A3�9=���8�Z��2>dyt\y*(�u����V>o^�Ϳ,j��>K��Y�TާӤ"Qȳ~/Ҽ�>�X�\1;k�����Ȫ�|���1��t|f2��-�C�8�Ǌn3G�B�IW���FV��!�
�|8�:�c��u˲P��]Yskf��������*����{�������~Z�dW磵�N����g�|��S�0��Dӎ�ĩ�Uwt�.�[���� ��1�1� `��_AFY3�Ydi��,=�;%��'e5�� O)�Rr6���Q_�'a���'8&�H�.ͫ�4��j�>�ob�� ��q��О;B��Z�ΘbM���^��e,.�MY^���kN���=�˹�[���ѓ!�姑2��Fx7�R�¤��A��i�šj���ܰ�ߴ����|���t��}b���{L��k���;��`���}��i��������st���sc,���\��̚H�.�q���\���a�Hc���|.�UKé~ ������Է���.�Iܾ	F�PEΈ�����($r���� �Z�hRr�U�zXg��bĽ���);�{�ƞ
�l9�� k��(��=<�&�����b�V<о�Z�Ъ~�X�S6��zo���_J�I��/_�9�$�+����8P?��l	�S����}B���x��:�x5��n��sB�Sp�ilٔNf	n)~�@�n{�}O��NT���CZ��1VY��ܯ���1�"����)����g#�%)��(uc��ș�������v)w��
�~����Ҁ2�y��@���ƽLj�=��6����J�v���='��&���������e���Hׅ;�0�N+�:.�`{Ehd��!�S�ڙ3[Mz�[ڹ�liU\�K� �	��H#�b��{m�ܤ!�~�'�n�$��܃�15�yT#Pudu���+���<�����/c���G��.��/�+��C�G.ӘSh�)�D7[����v���ݧR�Ǹ�B�p���Q���А���8h�������%���:���U�Z"��Ȃ ��oc��B��S-���HN���$���N|��:P0P��p�|�R��e-��Xզ��5}گ�벫#�M�\��G�]o�A��O��
A7,�l�u�<l�sF��m�y<�bϤ����?]�]��e͆��Z���v��I[�R���	����4Z���� �|-�T�P�G��ڻ��>�����5��N�Nj�$�ϓԻ��p� �'�r�فR[f.8���|�Ű�˟I1������E�H��>���+J�;U?���'Xߨ��\�#_}�,�p��H�O^@��"�o��5�Y�G�?���K1��6.��6�e��O��|��H�uӍ�ݪ�����Ґ���0�>�ʜ������
�(��o��߻���T}-��n�m����1yP��^$����T��p�9��E�cr���L���b�! �v�V�8��햤���C�j�.ֶ·Z;���cH���\ �g�ݰ��UN�b���__I���B+tpBTtRf�|�hzK�<�n���l�s�Պ�tW��v�#�f�c���q�[���uPtސ'�]���AUe2[�x�A
��Ҕ?���<��׃�9�h.V���޽��{(z3�( ���\R��b}F{�sY��+-��D����F�C5�Xѫ	�?Hk�a��#�*c����6`9�ɠ3�פ���u5��/l�%�	����h�I F%�s��Xr�¿��:���1�����������L�`8�R��پ��5�{M�u1�	����<�C��d9���w���l��aH�u�"�#E;P(��A~��w����	F0|�bb��vw�?/�a^�3ͿF��f�� jY��D�V�,�7���{\K���Wg#,�mq�}I��L�(N��~�-��Gl��2��'{XmR��[�TOe��HH��ۢ�!JB$P�a�4V$V�GFcg���zw�Nӻ�wa4X���(�z`*!�7�4}pM~���.
���cL}���<3*�|�O�c6-{:o�@�����$��X�gߩ�o̪O����ƞ{QY�8��/�tZ��!�q�A��ػ��_��TȮ�4[�m
��9� ��������(���ko
* ��@���x��ا�;ҳ"�-Ϸ���b7���>$�Jb��-!^����-:�/�g��B��E�'Z;-.:�)^;���&:#|d����SO"zz�^M�Um��Hyz`p���<�ϙGN�#��5MHj��9>"p��U<������"�p���T�b�K�o�U�ȘWK�4�����UiI`����I�ܻ��:@2��:�������������TJC�a�k��Vx,[/�P`W.Wl7[nò�A��1}�w�L��yY�R�_�]Ip9�9~A�09B��� ��.亄���I�׉;��h�/��
�؈_|�9���^;��D�f���p��C6��a��"�@��;��#��P��c��en�u.�����Џ�
��gb��Ծ����2�}�]߬Fp¿s��#R��I�H�m�ˈl�=�~%��;��!�������(i'���,��Ƒ%Aa����0�g畀���]5�h�f���:V�c����AW����o�S�M�d�sN��	���Y1H�����f����槹W��@��;ʢ��>x��*3U��4!�_V��{�������o���["/ PUa<c,���8�*]d��7�q�rޘ�\o{A�@C���uG�'�n@+(�.�Z���B�]�	�2�w�4���۹���߅|��J�3�q_v��P�IɃJ�����
���i�r�k�@�^�� ���oh�FI=+�lm��c��邍@�͠ش̸�\	�D�g�a~�jܦ�d($(ΨtL�w8d��j��X�AK���<��$l����a����bCP�o�4+��L��BT�{��y_ݘ߃7Pu�W�R�����O�w3����S��~�9ױ(�wb������{��2���z��mҕ��:N��{^��&7}rcb�F��X-35�g�!zPC��Qtd+5�-���!Y�������M�ckL�f�:�b2e�����B��(��#��c�؈
�m�d��ȟ�o�W�q*�a.iF�X����''�N�H���l�2	zE<�`��U����#L���$io��\a����ې�O���Z��/���hv/z������+�?uJA�R3�N���όN�:��J�iWk#��4l=�#�K&&��ԋ�=�v�<���zMb��ٙ����c#B��s�tv����q��uS��)�U��M(��;�|��g�O�)��X=x��)vc�8Ւ�y&��rX���>�EԱPP�Ad��T�`Q�}c6Y�\o|��=Vq����C�S��Oª�)N��7�r ����P�[�
�
2iz�A����v�q��\�^� �;qܜGǁ�H����^���Uəm�H�8t"�MX��?Dcby{���qZǻ�5_1�Od��H��~�O)��	��C�hWM�`�n$D��N�- �Ĺ4�;E���m�ٻu��Q��2D��M�Z����2C��x>X)��e��/�!��(t��N��r�ϸg'�F݀�~jE�J.�����ge�KN�����<r�F@e�R(������5B���?d����Cm4L�>���4�D�v[���t���L7�&�`�,��&|�f��=p��CKH}ļV�Z/�Љ�����/=�=i'M`��
Zs�6D�f�H��(���Ôn���1�J�|���崠q&�G"ȇtK#;��]'֢�qY8�v�f@l<�79���a�?;Y���᫒ik,~]�
�N&�2G���n�;է84cTm˛�ޕ��n.Z�r����/�����F"��|�� ��P��`��\H����� �B��q��R�;*�1]�����8���@P���X ��������];Z�ީ���4r<H5dY�֔U��t������YM�Z1�뺂��җ�'7�Yt�jn5t3B�� �P���! E��$�Z��$�*���C�&LC#𐰘��B<�(��
%���#f_��abP�Z�eȘ�8�6ݷ�l�(i�K�dAJ�)��eK�kS���!�J!�\��:;�~��zys]�5�d;���ʀN�:&���H�\�{ؖj��TE�|����Ӯ��A>���[g~H#�#su�w&�L{��A�����m��G� �)���
��P7�ɑ�Z��W�H��V��}7e ex������gX���NJ��2����q�ɚ5I�e#Y�/ɡ&���x��Yi�o?���) �zp��YfFI�f�Ĺ ���釤b�y��*O�z]��+Zg�����iZf)�(�X	��}��̘:ͪÌ�� ͺ��fW��o��k�vN]��:8"���N{��e�ɋ���?#Ŋ�u1H5B��C�_W�6*r��q$�ַ����H��Pa.�>Y�'�s\p��a7���U��,��5�����}��oc��xTj5@��ؐ����S��ɥk�~&�jG�3�i���8L�8�I���sgz)���[�,�.��Q+�	b��&��M�]1c����;�G��;P��! ��`O5{�`�uK(ԍ~x.�)~t��o쯰�2[�X_��c0�R��Ϻ�{�L��מo�2�~v�xY�-xe���h���r	��h/���cS�qR�xP�T���D�|�ഴ��g��ٓ)y��m_�U�	LΘ=� �gLW��O�j@��  �
a�G̳�F��O.�2e��0�Lw1H�����_��/!����j+Nk��%�n:�6����b�X~���=�D��̨O��������愌�7�蕛��)��ČS��ur?�x��u1U<4��[6�"������7�K���x�����K�		��^\�+FT_�rm�^�ĝl�c���v[�� �m!Ne�A'�o1���k>W;�vD�$�/�3�f_ɁaI'1�W�����z�Ƨ��Ҋ�!�o:\CV��,�!���� �T�+qO�B����0�};T܈�pt��|����ّh�<3h�H^3�2DzË�)���1O(�_Mp5�>�8�ZE�A��k���+A�	ن�$��|o�\��>i�W��/O�g�~o�ذ�&�n�PK`k�HzmdaD �3�0��Nqj�"��LEAg�������5��?�i�@�=�mj��,>���_0�#��؋*I�Q�6�(P�5s�^/��P�>Ck�SDɡ�kwz`C�`�s�T@kz!���o���O�{����;���"��U ~���ʐa�B��:����B�r�m�R��A�ݣF���X������܍\(�R;kۖ���KE���z�8�jK�?��v�O�y<��N����%]b��ʙ�e����qړs�x6�M~|��<p�я{���$IR�q�*�60�9�Iv���xnwq2��F���.�(�T(�#��Ô~�O���I��-����J��:؁��W��S�B�wG!�l_�{��K�����Jx<�N���*�|�_rh�U���׻�W�"�jP+�,e�HT�^h�&�wb�F��|tN��]D�ix�ȥ�T��}iz���G����C�jc����`��`dL�Vl5FQm�gF�o��s������o ެ	�]������p�*!�aʩ��ZN��!���n.�.���䲓��t{'�Uww�٧� M�<�ߠ��ܧ�Z�C!pf��R_S#�(���l�~��b}8Jf�T=+�"���Cv��z���O��c͜�L�Փ)��8 ��²
��z#����! �g�y����ޥՇ�ޙ#Nc�h� 4r`Uw�`/�x,���]�Q96���kն=���! "I�Pv��3P�����`��G����?/�מ:�k�'����[�d�SУ̎4��l_M��.�� uDρnh��<��sc���e�7�}��տ����s�����8Y���@X��̲g3� ��;�^�E-/��&E�>���[S���Ѯ�R�@-���;/y���]�m����4�ф���s��ʓ5ߏ!f��
�3�������ps����Sܤ��j���ӊx�CC���n,�׀�þ�?](�x�}��^���y<K OKT��5{
(�%9c��[��Ф7���qM�6�������n�О�X!з�tu��)D�0��+�C9�zo��h~��w�=��>њ@(�[ZV�v���3t�5����������w��e���NY?m������>)�Cn�G1M<c` y`�Ɠ�]�.� 5�w �����%�@�i�ʔ@ViL�iF�w}yD�H^��_��ny���Gh��;��`d�`&������O�Ĭ��ת���ҙ,��e��o�Y��ϣ�4�nQe��*?M��[ᡀ��chv�Vi��ZŰl��!G����d
���\��W��m����[p�dm�G�JF��/6�+��=�ҕtgH��{7V揯�
7�XV6�@��^]���vL�U�ؕ�3�\lq�mZ�S�ͮO���z��@�k�ZX�Q���x,���Y&4��xq�n7X�\`u�t�
�1����)��|f��6C�m���hR�BYa"91�D�mge�&�r�w�%���tkU�eZ(���P�x?�Wf�^Z�7�����h��병�cʾ3r�ܦ�N	]<:d�I�ܹ�T6�B�KQ�~%L��j��i�kbeҔd}���YV2V"Ե�`�}�+��x� e����^L�2J\9^����\��1�Q�B��A�ݗ�m����CHGGj.#~��f��$���߂�X�@N�
����a�]��/(P�w���ڍ�����^O�(�wL~T���!)V�.���Cs���9��I�)�8�'�V���G{j�����`Y�n���/R��"ɢèo`s�3Ź@���y]g�����	�.��9��η�,�
o:�P�D�a6���sp���A����M��)t9u��k�:d��<�o���e�iŒ�9q��v�m�7j$��������ȁc��� �o�lBg�08$���@NZ}]Z�sM��� ��_��J��mCj�t��Mň��%�2\�5u�`����KwJ�k���6hU��N���6��%��KBrl�l?�k|܄Tc:�irðq ��4?a�.�e�/:Q���^eXfV��D��C#_���v}*]U_P�*[����_�6AZ��e]Sq���|\��3
L �I��"b�����ڨ���#�xN��h2��۪^�s鴲�;�U�Fo�b�lբ��(�#:���7/��*����۴�@E�IFG�j��,3J��jk��y�c�3��7�DM���W��܏�[�'�fpY��u����Y�i S�ؼ DZ֔��Q�7�~����K���>��J��9�����)���.����ă���z��5��`:N�6�}ɟ|B�n�<	z��L��+p:��ֶ�n3�XM����;(`�.�0u��6��!���}0�~d�Xp������:�����̤W
�/��4J��lm��5.\ğy�Ҡ%L���6���Dc�xy}�k,�<�[���Ӭ  �;�4��>n���#c�V=�%�PbѨ�\��!Ϡw�/��ꟙEÿ�;�\�	��k��>�?�!��~T��N�R7%��%P#'�)@�j閷���Q�eCe���_��G�\���^u�����Z+��o.�o͖l�Yӝl��A� ��_�J����PS�nT_��	OTlr���0!� _ *��. ��&kj")��(#�v�=$O�<@���/���}�L�}��I�8rƲ�C|����Pp����A4�臼���ɢ�9�O��ŒI����<椲&s��(o$�D2|��X�kS����KR�?��k����$?�+\���=�+��G$iG7jжi$t��Q!�^�W������@��X�W�8��B�~*����ߩ���B`N�gU�;"���W��i�c<GL��i�������S�-�aX`Ύ{IqD�AȲ���M��ۅ}jĜֺ��n�ya�
՞6�����2�?�PK��G��)��$�Z�[�QC��M%�`�mm���P�;��F<Aږ��op^*N��⿸��θ�9��?�ۙ�E��3�%a��J���
��fj�6�%t_ڬ��
�5O�қ`��e]n�F��B�kf���;!��2�u��0�<c\Ա:脀\�B�,�]�h�>�=� R�jalw��h�G�����%�=�L���
�W���������`# �r�%�h�/?���.Kn1"ѻ�	��VBB��g�ݐzv�
悌,X�^㻻{�\��.��Bp:��<���X��Vs��^���֥�L�JGj.��6!�Ő�g}�Hu#��&�Z�&�G4,���M����Z��ڢ���Q��3���ǚ����"B�X��h���} ���Y��:�r���O��zA@��K���'��[*���6M�t�Я�t���X�r��I}Bs���)lA���E6t)��N�v��\N�ޡ�5�k�����|�}x�߼��p��	:f.����'T+٫���@�]
��/��,<!��PX��V��x4-G��J��6�$��6�h����A�^ױ?vc����C%1й��&��}+\��A�Ѝ�P
ı:�FǤ�$H���6�ǣ6)s���0�L�6�hQY�L}�{����W���)m��v\v�棟B��s(���\���"*�o `5l��F6�T���a���M�,�n6>n�o�܌B3�$2�Ǵ�,��H�l`_.E��;��[�i��q�~�e-��P[��"t����#�����h�:0{3?���.��<%�[�T�k���*MR*��[Xr���f�>*n1�=�g՗�Z��8m�;�N&v���$�X�Tl`�g�l�	����_0�),���q]!�b�{�c
�)eA�� h�fv�g�����֟ZAՅ�3a��E��#�����K?����6�x�x����Ԇ�h�I�=��`��BAYI�������"J��:^�x��39H�d��x[REe�<��F�N�f4��;+z�|����nsG\������c*S9��!�0�/�B�~S���n��8����|���ú�L	;r�/\��+b�<	R�I2���iiy���$��
��d�L�7:�(�	^iJ�μ:�4��'&��F=	�/�5�������	�Y�ǐ��$�O��@\yB2�ZPR��#��d;��pX�
�v�Щ+���x�b��~D�B�o5KZ.#�;J��V9�^-ȉq�6��k,���9�-\qf���:���]'W����T殉���C��3-��D3�|��o���w��\:�މe�P��d���e�Z&�D��2�Q�Kj��_�}�쒬��m�umJv��r����P��j*H�yN���0��\kڪ��_\�S,���!��e���~��YaoÔ|��á�� M��mO�1�x�.��A���0\������9����O�5~� VI�{O�Ms0|�뿠��K��瑊�XM;w
�b"[����.I�Қ4�Q����kh&��\��͞�k����,Է�>k��)��)5�����/����W4��.�,��&��� ��-�F��R�s��L��sQP�P���k�ٻ&e��~m��R��hK(�y\�7�O��`&.=1{������[�~͏r��
E�
�;������H�7L(��7�=��Dy>K����>�cֻN�ǥ���u����B�N�*�ؚ(T<�c��v!���������4���a�qU6��YE�'�6������xq]ֻ�U}
qF�l��#�֓;"E�ݥ.i�pj�aR 7��J�T�P����ǂ�~r'��j��E6^�P�(���?�I��vf:`k;h�_��{�ɤ�������quWP"�#�UB������G��8ՙy?�)��Հ6�h7�����Rƾٖa(�������.
��O5�Y�Q���k��K"�DL�I ��:Φ>�X9�Od�[�e�f�;��b�qΥ)�2/��#���Yۖ'�,8���?��T5�ξ�vd�ĝ�X܂�,��.�a�r3.'��ȡe�u��.��.�f̸�q�#w���
JS�j>�W|Y	&$�P{h"��H0��i�A_=Z!E9���	}�X��a���S�t:SZ��Xm�Li"�m1��^_s��.�`$�C?���k�J8��>N_n��[�����*e�Peu�c���l�����m% gz�J���CyVe\�j�O})R�r��$/�;���g���En��yJ�cRm1y���`��R�gb�Q�,'�4�j�a�tt�6���w@�v��'�1P�+j��C��r)��>i��&6�f�ۚ�SA١kS=tC�8�[���1f������2�!2L]�Ҝ\8��qVe��Nb\�`�;}c�� ���`*d��|��~����Z����u5zW�-3�+��#���`��+o���;1�i4���eAf�P�D/�t%0��ɍ��J����Z����h������^4Ă����yU��Wl�Xg�mϾ���9���;L��^U��VXTk�`>�X�ͳ����|a�Z{yv�����W�&	�f�����:�>y�z�]d�[�w'��?�	�|Mv����I�Px��nQ7Cò2�-�JFO��堉f�hX�"��� *�E͍�n��~ȼ�%�G3h�Ҵpt�����I�>\EW|��tv��֒�Ӓ�f�f�V�º3XA�������ȯc���k�P!9�c���3/��Ы��7����AD�S�=+������B��P>qQ�IK�p=և�j���?�s���y|B)���d����u��OK�=�7�"k��!h��~�Ҹ��U2'�H���s�C��oh��R�?��R���N���M�U��������_�~0�$�P��U� ��� �5���̆��28�	����㺈N>N&�ba��gNxZ����mDO�� c�(�c��^(�b&T��f���eDi�v.������Q|GK��8�:�
|bnv�N�������6�u_��F����uX���+Q'��.��σ\L��3|]���x~oy_��Z��|���_�*�F�Z��GW�Gs޻�Jj��"��ѩ^�0ct,�V��G=%Hp��Z�Х���J+�[�N��@��6*&sq�V��7���:4hAX+j��
����j�u�O`�Ú	F]�J�I�"Φ����8:�x²|�ct�RYϾ�MX&��6�يk��Tk�r(m�<��=����Ƹ��2�x"aO���L�f��1v��N�~q�.��G\;�>�霛��ޟ `���d*�e�����������-,��?
KZ��o�p����������,�N��06Z�����1� ��{���� @�K9�}	�q����
�X�ّn��(���j��uղ>up��Q�9L�F�����<��a\�;\�x役أ�&]�<���&zg�ը���9m����K��!�ivBB��:E\k��*8��gڻ+mN���xZY�Ʊ�S��t�߈�&}%�$����`t�r�\f�xd�M��Q�X�:�����κ;k���d���&��b�%?���	����=Hh�0\2�/;�Y'w�m��cK�����6��
n8���`�;�ƨ���wa�����zL����K=��d��?�9���<1F��߳�ŉ�L����\ϝ�%���"��,� wm�U����
�˶����A{����rȎ7)�����_+�x���at;w���u���Ԝ��I^�靑�X��TI[�C)����uln��2nM𱁌W+Ch�'iLO�jO�
���
�}�Dh��Q�*��s�M��[��+Y��Y������M���r5�7�Ad�i���s�2-̇��FȨ���3r�:���D�O'�v;���}n<�Os��Zm+�4CP�#��݂0%�*-4�D��`�@��khL~KIq����!<���Bu9�#M��G�#�-�L�D漛fs�vVlm���_�u�)Q�L�l��$��!���P�����#y�^��!�Fζ7��Ӊ�=>
��E��$N��9
��5 �B��K�h�-����$1��tMw��'}ҋ*)ױ�S��m���L�����v\�7����{[��^�s����{�c	ˬ=���"�����\��Y}�u�:D�	���:f(��Gěӏ`]�yü��
=�	 ����v��9���&�i�mZ�܅��PD2+E�~֜sP�4�'���cn�h�3z��geE������?�l���iS)�w��&�V }����ϫ���}+�>@�$4{���V�-i� �N��6w`�=��qnh�A�q��il~H_�W>�S*M*!�a����e�u��VX�����V]3���7�I�R�_���$E��A?1ߵ�����~�?��5�o/��D7l�c8����f^!�t?�,ANnv�'�oI�
�]�� �ef��ʨ��f[��^�S�(X�In�`j�k罥5��C����T�rI�/q%x�Wv��3rCP�]��O�qZ��H"B\ؖ�608?��� c�vۜ��P���\�^kF��t�Yu�-�Z����
J���%t���Q������[�ֆ`0'�}���}0W ���6�1��н���t\@��.�8ao�����(���$A�xӵ/z
���"��h�n�R���G�͇����k�c�<V��ٸ���"�Y�}O%���Y=�2z���|svNc�MND�7\����형�A�@�$�fv��7b9��H&��o�N��tK'�0ϏCɁK�/9+ਜ}Aw���(�Xah�{��t��d&F��b���	��S�7HO,M���O�.�^���1Q��9 _CB�S���@���v��@hoC�,�a�d��]�	�yw��]��5����1���9�]-�a[w�UtBN������+=�b���έ��4�t����H� ꒦�	���^�%�h_,�V���#�+\�Ƿ�r�[o�f��[�p��+)��>t�G�tLt=~f����R_���� Z���zrU�Vh��(K���N��gs��j��O`����s��s穸G�fRV-n\��ȁ��c��_�5�JL�
�T�b��[`���n$_q^����5��qg	 ?;�r��t�|�cQ[k�'���ARE�>%�uӽ���e-T#N5	� ��sI�	�D";�f���;�N$2\�^�I��ާp�2�|�[���+��[����t,�O��<�<�3GI?k�-��@����d�6g�0)۷��	ߣ�B�2W=,���Wu�"B��6v��Al���+}T3Y��+P�L�}�.,�R���=+9�Ɠ%�t���o-���^p��"�|��oB��P0��P-QYI��'��zrX�j��@�sM_{O{��e�G�]F�n.s��tH���s��sR, ��Oc����'|<�O�^2ߘ�)��6��'b{��i�f��������
�,�P��]�"EX�lݗP�M�g���q�=i*�MC/�ZA�W����H�M`�;)��e+���rO�#���{�I���R�pJ���h��EC1rI�i���A��:��,B�	�J�ԧȝ̵�����|�Y^!�kc168��6wGC�O�'l1ĺS�î�)�
s��k�������0~����˿�?7U	y̙m�\��?Fq:�8�H��b��>o}��p�ԝb���f�T������v4�c_FȀ�v�Ԭ@ yС|j�1�X�%9o�1(���b���:ځ֊maf��r\�T�ـ{�x�U��܈I]�n�I�9YZq�F~�
�$S�16���"��ȃ�� �S��h�8������7~����tZfK�=��-KW�,k r�t��{q�G-���W�b#,�*��3�R�77���c��ul�AvJu�V����I�����4��$��+y��C�UL�p9I�Pd%�7qT��!Mvb��뾙�I2�Ke_�ҙ2az���q�@��a��'~�Wu?�fҤ�mL�HLE[M��L���A���N��j��H/�M��V�ƾ8�������qC��^���c�}��Y���ؑ����:�ڏ����g�W�E�T����-��f�4�A9H�������ϫv��/���voH��k�)0�������U�2Ӎ~�}V�z?.hn����c1���|��ڌL�O��n����}ˤ
<�=���tl�����B��xY��_1�?��\񯣳U�N]Ш)�G�.�̭���Y���@�D3��7ޘ#�!3ܔrk�6��R���P�������1+�L�,)�᳗dW�UQ�3�S�r���py><v�fk���Z��%�����ʈLξ#�Fn��D�z�zO���o��;����և�>J8�K�Y1��kB�~V��%�[�n���i��8��0���&I��/v���+��QF�n=0,o��6�ڰ��{LE�"U�K #��p���}[�_L �靄;J�����򞭹;p(��>.������2�킵0O�^-�L�C��|�*"�c4��%�A$����.�GC�ј7ڙY3*��Li(�l/ [<�3�)�f�(O;]����(���\�5Y��w�\m�<V+��|��e� �=�hU�(~�=^A�t#�G����q���WY��5 9���p�L��XK��&]P�	pp�0.
}d��j[)�:M��9^晻*I蘒H{WY=�*߱��wˬ�!������I���6A��׌2u�.Sv�i�����^^ �c�B�sl�9(v�1�E�76W�O�Q�0��M�Vه�ȧ3��{<i^��څ(�kQZ��}88��1���Q���-.��"����d��Е��ӫI�����I�1�X�U~���x�xYN��{��*:�����,#N��2��>+y��p����`9ͽ�nಲ
��uÈ\0��x�D�}���&�@yc�u'-iAWk> A�m%xc��~J��Zɐ�KDQ��(ϒ��֓(O^:�PG�y���V�Z�Y��R���ީ��.�ƒ�{Կo{�B�B�c�嬺4�u��F+ˬ3z!{E�&9�N���4����5����6���N����f=�z�{�N��f��\�$��
H߼"T�����:��.^���}�a�j��n�L9�f�� ���/�[���@ʛoBצ9~p��x`���W�ɤ�e���k����4R
0ۻp5�5(ă�&���m"]<�&u7kQַ�p�-�[%e_v!���u�L��������&�ަ�N:��;�k�Q��z�j5�с�o�e>�b���4�+5M��:{��"�Dw 5��<��(�B��s�6BC��A�Ĕ!�K��@ bZ�N��]}	�� ��r�����(���"3�v�*W�F˯��U��S1)×)v�̪3���@C'RhQ4�y|f�� �e?3�Mv��N+���(��kf 9{6�t:�k�xã�(+������|ͽ̎��H�B�����u�&e
ac
/�q�xӻ�bk*�U~��0�D��i��mu֭�Y�"�-'�ԈY��M0��X_5 O �� Ǩ�Ȗ��d~ �]F���D�7���e��{���2װtZ��������*NW�H��qNM"�x︢ SI�Ap�z�,P��>.���Ί����YJ�A.
Y�˴�6�8A�1N��^���6��6��Eܞf��N�.|��u;�:����a�*S��~��=0}�c�BMMAa��a+K�ɎzY�C��	�?��YT���9�im�S�U�0,��%-��I� �.0��v'�°o1,�F���ô[[�z_i�j� u������+��M_��t�#Ym���p�Pq}+լ|���r��m��O��x�K2��Ŕ�܍�F�F���+/��Fg\O�	���Ai>��a#�eaĠ��O�������@�p�YF�R�:g<����d�3�+�M���z�?v��٥^��iw�H5h�:��㞫��)�k�Bs�����~�E�d��-N_l�[����y�X��^gW(G�qx����p�����Z����t�]s�_��p�ie&�<"��8?��le��j�� EygQa�c%�.�Q�'Ua��}����)��RZ���B���F���*�fs���/���/��@���&�{�8����ӭ��e`s�~�g�~p��G��YD�s�� >-����N�(sE�_�o��=ɳG{�Zvbb��q�e��� �_�%Z�p�5,������c�W�Dd�#µ���ɖ�d�|���T�Q�u��x��{K@i�T�"r��
%�Vg��3�x/���w��n�S2B�LJ^��,�4�EDw5W;[PP����6� ?\=�80�t\pn��ՠΙ���\h\ɗ2�S����������K3��z�h��?�R��"�V�;��)�!_�&���p8�a_�t���mKwa=Ĥ5�4�hZQ��U�Ʃ��ɧnW�Q�=��Vu,�%L�fv5�<BZ��#�h������?�z�q���5��8U��T��E9`�/�=@ƛcN��i(xjg>8��d����M�MA%���M�l]4eZ�e�����r��m����UA�yz���m�#�"��n��;�Ya<!�0X9R�شp�	fUZ�rp�q�L�_�ꅵC��NUei�xt����5�#z�a�k��V�+�)�*��Q���w��jz8��`�-�IIc+��ة.oP��f�Qg��G�j��O\wB��~C}gds�1o,�\�O��O�d��@�	��<�V[2Y_��2\��*��F�<�@���q)��Y���+`)�<�8^k�;� ]
���B�.�2p�2o�r�r�\B}B[Rj�9�<ßB����V��-&�ʞ���9���hg)����!�!������\TI6Y��d�@�J׎��!Q��Ml�w� ]?��������yi+uq|�j��G�zd�6����f�q����Q/w�Z���z?�R
<���%�<e{V$�(q���gt��da!�D$6-&�P+�5خ|#�����a�=��3\���id�:�A=ʇ�+`��$����p��;����a;P$���l�����g���k&�i���&�o��Dr- '�\C�h���~#W�/�)���<6A ��}��X3�r(u?���%gx��mh��B�ma�_��m\���wIO������;�FU<elw�(g�~�U��2�#�Y��l|��j\!^�~ƠDcP��7?�h��h3�r����W����L��/�&������3cx����V��9\f!nz %��Yrݗ1��I��o&�U|ҝ�+n��S5�6�ؼ����jCYR;O�|�v|Β�qWZT[:�"�Q�}�|�lZ�=%��=�|!��G=�Q�rC1�J�"?������b��M��y��E6]��6�Z�G���@�;��Tn5KG���">���ɢ���Wx�O���T2�ٝ��9��Sׯ��ő��T�|>i�.��b"��1���ְ	D�~��G-��ɢ�d$�?��'V��&�?��m�q\�n��Ӓ����`�)�BI�\g���*Ex+>Ums�Ou�M�9�T�:�>F�_JjQ>f�gz��M��,u��⇎mB$C?�i1��M���� Gg���
�V%�y��G.UZ�aw�饽�-r��B�D`1��$��X�u��Z�O7+D�`���W=�^�:bp+Q��B���9 ��qҀ	� &��TJܙ��MwsC0���C
!�{%ܞ=��d�va�g�(�k�Y�{k�Q�H��b�%�F�8���FA�Pjy�����N��̛���j����"^��K!k��2��NJ
�QHN�M�.����� �m��X���m����Ɍo�q��5�휫P�NJ�!��p�����KrC׹-`mC�+I�6!ޅy�h�Q'�Y:ټ�E�������<m������Y���H�D
���G���8��f��<���I�����P��nd���$=���]������S�~��ϗ5(��p�V��g6�M��n�U�{����-�G�-�D�30ݬI�{��AŹ���x�wH���r����`^Q!{�3�9���ѹy����V��܅���m)ǥ"n�ަ�N;�b����G0=a/iEħJ!X$7"X_��`(1���4߉/��E����Y	��$���3WM���9$e��R�l����u�@�|����7��Y��z��t:%����� �Q�01	&
KǮ��$p�LvN��q��A�|�1�� �����<'��8�^�ʼ"yV'q�B�c��b^��'qT&2�5��k%R��+7��|��G����Jؤ������l�L�l��{yI3Hf����#�JμUd蹧/���)W��������j�0&����=�3aDD_ٱ�7~�He �r�r����1u��~p�)������Ņ�������=�ڷk���k7J����s88Ŭ����gܚ-&�D�@�<]��g����a�׍p^)ќ�ų�\j�p�����B[R�@$��h�b�����P���+yp��{]Hnr"��K4�Źm6hr�z���b��)�������6����a��� h�e$��F�	~�������S����gtBҶB�%ī� F�X�0��87,D;����Y�Ȣ���V��F2)$�D;e~r�Z��Q0-�(`�#��r��fE���m�3F'&1RlK�b�>s\T}���́��5.�<��d��V	�{'G�2�4P�\�=gz��o"��CM�ִΔ��Bj�ϒ*&�-�@��{�g����5��cǐ��p���oj�\i�W���5S����\l��V�I����������yX��2�[Z���M�3S�?o���������UЗ��b�����^@ l���Н˴����@ǈ}(�=�38>E�L�l!���#"�Kɐ��'�K9��\��ex�Ԃ�!���_������]��s�؛$R!�վt�S���Z����Һ�r���r��¾�=��J�Uq�+L3,*��ޯ26��Ů*^�[Ǹ��'I�lU�W�TBf86:�9����,��W##z.���8��T�&kRH�N˄�P!���Bk�[��қ !%=Щfuv�=2��޻u��@��e$�ƞ�gnP�r,���x/��I�z�A�ܽ��	���XAH�5��2��c�E�V�
�4����μc�GgAׇQEM�3�YU%s��P/�w=(�aY���oMs`��V�V�Y�1��/�k���oW��kjh����`���G������GÐ�=���n��lq��-��"E���R�	c�� H�w٬����m�z�]j����8$�ś����X�a�!�&�o�Byjg��ۅ����j��O��Y��gY�oQ5<� 	"Q[u���Yc�D��Z��ѿ�6��-����.�X�'�L�yː���<��,O~|���XE&�
1�3t��W�iF��{0����G*���5�ld��O�"��#DjFD�{
@K�L�w i� �����ke+�
�;�)�aҾ��k���#���IksY���N|�xqJ�|��5�ݸ�<�R	�ì�g� �+�����9����X�8�{[���I���N��)��{N��sG��n�8x����0������Jo>ջ�����5�\�[�3�G#`�A`d�Y~� ���V���X�y!@�f�k`5��6��Ȇ7Ώ2J�!�� $
M��j>¤�^��L7���i��lj�k��3�W�	D��v� ����Z�b�a:,1�b���IK>np��ܜ˖gn��;��О��>�'oB���!V�s|�ܓ"���ʽ��8І/=H�P`G�N�����P;��p8�Y�5|!���f��J'o�户��S��C26�ˡt5E"�v�@��-�$���yv����_Z�]��t�A��ȇ����
�Ҍ�No�s�E\<75��Al�����<�P����~��O�I$�>���χ�Yڢ��Ӛ�:��FGrJ�'��A	ܔݱs%�V'|��N�#6����	ZW���G��ݠ}׼B���@tb,2�Zt}3Z��sd�	�;<�i=�V�0�9A�L���><b�!|�ˀ|��cC��SPs�!�6��9eK%���j�a{������83����s��^�]���$�;=�`s��.�Yj'8k9>��h-����v�D/�CY�NW����>	r�3��wG�����5匎1#�(�h��5z���;	��qhc|�3<}��*�(��>�a��#��e�i���j���n��b�R������?6Ǭ(.�^��^�\�Z�)����s�����e����Bgw~o���d�HC��Ye<�:��(��0�L��kT��u{������O�p��`ܩ�����ݳ����ʠ	b:>=emEm�b1�Uh�r�fy��<���W��9��Q6���i��x׀��zʾ^�V΂];ݗ��T�giw�L�Z�����0���^F�W�ͮ�I����\I�v1{��վv��U��Ͻ��Afd;�"�\��@�ȍ>)��j��6=�nT���'��*f\	\q0&/#���:�.=��	4-��\�]��K�R�B��]���pa鳸������¨��!��kR�_y�!�"�F#Z��T�6�%���~aN�`��zrs� P '˕����5�st�����C��c4P���v(Op�=7����2X�.����#IY���3�f,$g��x��?��$*�w.�+�Mh �7t�]�����*{�\m9m_Pdrc1�ݾ�M�ri{�*�$ڪN����g�K�" �C[Z5� w��a����ٮaXEf��Oe�i�w�����;�_��Ȅ�GM�,a�������L���"q`�T���M�����$ik�Ռ��rq�v3�+jT86Q�w/1��|%�>7w��iR;^��"t"�`���I�v;��w,�T���������@�i��*d?<2�����v�(A}/K?�#������[O�
Q����4��z���������t�?ʀK�d�}W���+EN:�D��\������H��2/ZȪV��� �����E(��h��)/���=��ٵ�;������pT8s���������L4U�
��U�P	ć���.9j9Va��xj=�nu�̌��U��΀�X�-������	a�/��7�9	u��a?yE�9���K��ߪbx8�����:Z����_K��K�_43%���m�-��c�Τ���p�X���Kz��~n�ݒ��H]c����VuE�N���D�8K��j�t�e� �C*~dw���U���~�`�Ǯ�e�m�E������i��a��&�k��y�)���#_�i�	������f���"H�<Ld:E90���I[�;��.���p�����K]^�\�>?bXj���d�w��/���D�N�af
�_
w���ѿ.�2L�8Ի���r��UP���6�r1c�H~Y1#�`]�whI�.Xs18�,L9e�a9��-6 �����P8+�Im�m���܍�6r��7d��9�wl�E^1�G�/�k|{wn�}9
a��ۍ�tX��<�����2�AN�U�^L�H�tHQH��_\2��Z��2`�d, .P-D�E�� s��/sQ�Y��c�j��v��x96��qkO����e�N�-?��� ~(p�� ?ȳ��F��(<�>�܂{�D��/� 6VZ��% ��'V���D��U���{�=�Z4K_�����=�S��^3*3�����;�X�f��$�0/#g�Mƪh���ڢ�y���� �)�(�L2,LE�ee��a���6!_w̺K���d�$���
�#AQ���n����n���(��O�q~&5(��qI̏�G�_�+|�"؄8Y�G��Y�HA��֐pښ�B�B����%֮_k�sE��nmO��do��=�b�B5�ZzJan��ӆ�E�
{�	�d;WJbXp~zg��y%`A�� ���B��e�v�Qֿ^D;Q��A������j_����'����lj�_!����x��nVyи�������f��<=�z�,=�x���X����= \����%up�:����GmE�A2��G��n�-4�[���;����~9)��>a�)�N�"����{A4���ӈ$������u|��W�^ �!���O��x�xM�̬��/go}��W�sHt�V���?Ya�@��r1����!(!����F-�VG㝦���b3�@
�u��m�W����B��lw�$��)� ��@�q�W=p��~����~_��u�O��0�T[���<�N�4�1�&�Tc4�m8z���Ą�̘Nߙ��׫hT��[�3�����$&�6��XVF����*���>=��O��+Nˮ�˹D͸R��v�DO�<�1�)0$�
�T���Z��	��<��Ȇ!Ua5�H��,H
�հ�)��g,��k�^�����Q`퐋�m�E�Urcn."��w�ihꤪ��l*ʖ��4p�
w�9�k�w�O-�6�m��@�o������w��>9v��������'��u��S����c�h��]�#��.�׷���#�=ޜ��2�18$��&��0"!��n�c]����_���Hґ?�z�"4�W���9�m�:J��ZZ�N�˹u��q��M�&��A�:��5�8j�u_�&��?��=�$�7N��S��Ӈ3n�b$�g�!+B%H��j7L������4��̷��?�G�;�%�I��W�n�>��WDs���<��9�o�5�������{�{���qT]��d*Ư0��8��φj�������
��N>B�W��;��L��>yəq���6ӬS&@Ƶ���<�O�[z�[� �x!^���
[��*|׎M����<�1����P8u��'P��1�SS��X�w�s*D�iNk�a���T�Z(12sk�qG�ߦt_�%�#"���tD�M�n�өet[�-���{�NU�"1fϪ"�m�2x
��T������9/v�ћ�Z=�j]��kZ~#h�h����H۝�x\���\�A�~5ON �-7��FWR^1Y��[�"1hG��L{%�@�$MɐU�u!r��t�̰ �z�a�j�D��ܒ`	xCq�RCX�@D:�c5�����;�ةJ�rX�r� z��pm�� ��Qj��.�i�!�Ӊ���S�.����K��� '=�z�%�z$F�eOw�z܅��yQ4�8�2Ite�P?]�Z�!� Z������d7Fc�8���Y�B�0K������H���S��΢U��������A�*n:"-����A��>"�U�ς۸���}#��^
��j��Ycג�E)��g���1}6(�_�N����
��f��,1��R��E�Ku}����H�v]����ߤ�rOPT�ɻ��VE?�l��&��}�u�|�-�m���ÙdtH�M��Rb5�},Go&���Ҩƛ��&��e���|})Ji�~β=��e���XL�0�!�0�;�"*��ָ��h����T-V)�Ƴ��ؠX7���M�ޢ@Y��"�� èe8�k��	/�x����n�����[�O� ��f2<�t����#	j��҃�P�dK�ٹ�i?�ހ2K���(ne��i���7^=b��9���|����w�-jnjL�R3f�R栔,]�@q�O�x���7<�׷�"D�M���w����Y�5�F���[���T�:�,�իPk2��K�e4/^M�l���P�į�j�;u��b�{/��� a-u�����Z��JL�Ufܲl����^�b�+��}���&{,�r���r���7�%_�Β�Awb�)��8eEV��}8���țe��-�/�js=�so~�㻼� �_�CvB��[߇>t=b�ŸlO���l���i��c!�������Q��ڼr��ӫ�Atxx_�Çe�E�k��J�0�-�!�L5��.�To�C5�*�DIe��A��僋i�C��D��bd �C8��9$`�$�����v45_ZXjp���!��m���$&ϟ=�P�ۤ��ӟ|�)x68g�R!{����@'��h���XL��[��i��g��� �$��{�P��h�z���ǔ�,m��<�ns�C~־/A�,���8���AR�r
ԟ#o��b0�8A���z�M��ٙ��[�&D��-�8,�����O��������*�=���Kw���!�0�"Y�Z��y��z �*�oM�'EG� ���j��z����	2�<7�.�s��C"\��vߟ�z��%b�=Z�,o	A�����\�t�j�Y����.��^Tډ��!���:�J�ܖCHϗ����%�^��g���.X�>{E*kH�Svb�`��{!��P�l�@�����uc^&s�j�qqn�$�`�����M��@
Osol�L��W���sYjN`� ���ƙ黤=��{t����6��3t�fd{��&S/�zo�" i�[���g���G�u9"1���z�/�����)@�XcW��I���GqfR�c���ƻ�(�>0�%�r��6����:=$8c�+�~se�o��IM���A6HT�T`���@�S���\�6�C.HXO�g�����H��~-�&���o�5R�~������`�ö�@��&;ƐO#"?����֋* �4^9���S�A�U��u����C�W�Cs�X?���*юn��"�S��;�o3����ĎS)���R��k������zMܟW�m2cdin���R"���	y�Թ��~��^@���0�9��q�u��;T:��W�>V�{Ѥ�`瘾�!&�\F2�[�/V�<�~�@M�����9u�jEI�/��� ����}�t@ै���r�Y�D������N����c�hO��?�b�7� ��IP��)���\��*5���!ә-�	�|P��|I�c������(����,7X�����;�Y�h'�a��-Μ)b_;��'�g����CKF��A��_	6/Q.�o���>�M-H@P�fa�nl���2���JZ��u���L�p���QȬO���)_�Pԁ��Ͳ�ہ^*ٟiIX�g�-P�����0p��`�~�&*��"�ݶ�YPLW��T-����a�;�o|x���ߴ��M����b����.��Dr�K�\���+�t19��
ɝ�dl�\6㼮c��X���/���נ�Y�?�+'޴�dMA��Z!4z�s�U�;�,3��oL;/+\H�8P�S��_��[���{�*^'Â!Y�����Ĭw��U}���a�Q��e�8���>F���獓V�P�)���HSl�.��#����;�%��a�F�c�Y���G�?Y�������6��:}V����Ү��k�	�ENLWY�a�yI�ٴ��Kw�&�o��z��oB��[B��h�ژ�L �=��k�Wbo���=㈗b�!��5����^&�{P��+=���?�'�$�
���qE��7ir�E�����	��_�+�J�T���R�NKg3�cz8�w-�����j�S�?u�:���
̢���H�-K�&�&�-�����)�#��D:��������p_��#,z�&\nG(��/���W���������%Bp��'��� �j5��4����L�w�t����,"��e|����%�O�M�F�g;?w��*��f�"����ȧ�¥n�7�@+]2�z�]$e�i�T�9.��a'�4"-��Z�i�b���u��FVg��Y9�ӟ� T@�4{^O��]�>�T<Ի���{4���(���4aY��Onl�|��q��
�0�1#bH��[7hG�oo�:��F{Ώ�I�x����3����&B*s8Nl}v���Rqfu�:��6�W����::|�	�b��|[����L�����`����`*���H$\�?��@�\�� Q͍�����R�Mܘގ1�5���>6�Ϡj��kS��KЪ�k�a�1��G�3�UV�v�ZP:M	�n�y���.r��vPƛ�F0~�#�fR�����򵱈-�8��RੑBy�^Xc0���lFv��n����ӛ7Q�H��ֶr����S�M��y�����Ʌ�J�{�}�9g���h�̮vC7�%46+H�
���*��_#�
0�QC����!vZ��CL	�JP��Q:O�]�I�(�w�v�d-W[��U:��Mi�L��<P�˝Du�*�mG�h*�^߅�Q+ps���A �?��Q�zI�)u��9�#������My��O9C�(��j���	�TE�k0�c �2B���Ql��薑+���έ���5lF������-xLXL؄o��r�z�3��Xy	��Z��o�4�>F|*�j��|�
m��r�x$Fmy��Z��gp�o�����}������gO� ��S�4�WV����џ�̚*?��Xp7��#ᡤs��zs��}����9}F^xX���7���o+�D��q�-��t�*ǿgX
��k��u���`;~�"�#�
��t�!�햣 �
���񉵡��0�+4\�t�v�g.���>��� �Vs�A�)&�v ҉唅_����n9Z`�� �3!"�@�.9���c��e�}�0�5I&7����*�� �Pܐ�zכp] ��:ȉ��������}{�u��\m��}��y��_^��繡[�"�Vv�����ݿ�����!yy$:�ն�x�����Bb��NM$��������.|{@8��YR٠�V�	�%ZO�+^?c}���Tj�J��=��ч��h�w�Zn�ʳ�Y�]�1����n�k3$[���L@E��&����� �u[h�>5\��F�pm�6B�?�Q�륨�DnX!�ގZ�[��c��8P9�#�2>�7�*#ш�mx)-'��Xj��+��:Y4Oe��������NȱK��u����"�����c?ˍR��x��p�Q���Qߦ�5�:`F������Z��!���/�ެ-�[���4"j.=U�}��l: ���x�Uª�i�+9Y��'X��w"���Z��=��Ncx�?����h��Ƒ�t�'�<�)���9-��Y@	8�Yic���%m�\��CR�mM�ZJF݁�4�|�rt���gw+/(�*�\�7�g���o��*��P��ͷ��Fc�&�X�!��9k�ƴ�x����hn�4'�m�8\屿��žW��$B w�
�{^u�tR���"$�/ا7����RF��r�~�},Ǯh��}�sD��򲖦���h2f�J���qc�\:�C��o�/ui[�i�����f��g��e�ΨG�*��+�F��\ބhѣ�m����kfhn��.�z�q-��e`j��#���@�����\�t}��!n��1��o�5��#�Z�Td�z�˴�P�>�]�x4��#�2a�ۨ�� Q
4'�5�E)F"�CiG�4Ew��ӈf:��>��4֎�&{���v��=��9Pk�%Vas����$?*;�}t'�%}��p��8���@�{�z5�w/��E
�7u��W�b,�����r���>>oZq���0
G���xh>lw��V����c�X�k����o�q�>C�F�ܭHpK���:Ƥ�s�3�V����m��ۗ����܋E�2G���S�Ys7 �9��hz ��B!�_��U���<�s�|���}]�<�fx���i?���o�<@ɔZHCk����c;�����ݟ6&=U��;|�p|��H��0<��h��y;��H���.!N�r 6S��du�2{�I`��->f:FԜB�AZ�'�Rnrn��V��怗�K~̈D�9���/S)>/q��g�|/ֻ-�y���yJ�t�f��Ck���[chc]'� M�[:�ב�.�䚱�'匳�E�tʯ�l߁o�?1�y'��ԁr?q�Đ�2��-DmG I*x�dk�Ҵ@�jUZ���e��Z���%����'�3�ѭ��|��ym
��q�K�1�|N]�`t�A?����6�!��~����u>i6�~����{�	}�[��4�r��9���mE��=@�v_�	�(��Sc�Y�-�q��˹s��\&�vb���jZ���.0-j~\�Rx���8li��J�5��
�)>��@�Ϣ���p?�!�-�ݍ07�G"�����Z�x:��
�DȮ��DN�+a##�V�K��FՋ���6!ug���4ڦ]e��s�ou Q��$�yc�T��r�÷�>Ԍ� 9�3t��ћ��ְ�v]�qo`Y��k���/�e��?8���;�#\��#�6
���� �:�<'&�Y)�=F��b��5���!T񌱤/��!�M}'m��Z����ñ��̂3�m�̈́=�حO��Q>��b�kA��Q�29\�@;�uwXտ�ar0�/~z�h��?K@H�\���E�p_�AB����4���U���ajbH�k0&��ƃ�\Cw�>*F�y�
�_�(�a�����a�O`����:�&��k{�p�5lQWʐ��^���wәth�j�������}ʵh���IE��4B�J�� �e!��{c#��"HAӺv1��+������Y@F8��E�-n�`�+nwCjD�/���Ԛu����y\��Md���O� ���'r���8�0n1#GI ��<���0"��K^��t���1�&	|1Z 'W�R���r+bЌq���S�*r��Y-���~�s������Ӊկ���U1���{�\\�X)��d�OR�c��@�uy C'�j�����+R�2F�[��Y��M�ڄ��z nt�F����M
��R])W�׽�Ɠ����u	��@��C5�Kϧ8��N{�� /C�m�E@Df)�(#~�
{���T��TXA�.�Y��Τ-=M�L%_�=���m���PH��m{2�9����ְ��}��I��^��=����aT��p�d�9�~;4�ȁ���M�q������ ��k����ct�J�r.�	��Ck���4���;�kO0�=D��;x	�
�n_ �d�4S�V���2�%w����>]J8��������ߜ�� .��'2�!�))��@�	��w�uY!
��@��� %�\b�V��qr�%�-&��X�쿘,t䄃��*X�=�w�����)�P,�8Z��^�)͗���@"L�9�}밒�L~=�W<:7h͂^�I�	�p�~����f��^�k��W�a<9�OL�Vif�(�NK�J/��k{�UA���t�|j�:*��`�N�@��=M�!���_wU-Q��آ�����Wcy��i�qN�݆/L��(�ʸ�3���4br5�))���`�cs���݀�cId6��n�p��p �,K�ӵp�R&^@�Y�E�1�+����jS��l�����0Αn)~�@H0����t����h"\���M;>�z�<��C�wp7�u�7y<��G��Fryȓ;��B�}�Ēs���{���BZ�M�ѷFd
����|�2����(�>#%���o�����ʿ����E���^�ɪWB�e�T��st�y�?���t�NI��C�|J�����*�W�)�f�B@�e��0�69!%X9�S	y�-�+����w~�t��Xqq�I��ݩ�pЇ��h�{�'Bϵ�A/��*JT��#�J��te�n
$�W7\�c�rG����&�`2�*G&�Ǯ^Z�5�;Qq��0n���z�Շ(�0��7��S,�$o)w�e@-~҃Q+����.
�2.M�!���}�?�OX
7?�1 �Y��1 (����:(mWA5��R�,u�c��-�q�m�&)2r�gg_ޥx�&�!N�Ȣ^�A�v�N��^ ��7������d��d�<��dHix�V��l�`fUyv��ژ\�Kw�� ���� T�M`�/����\�V�k��˛Y �Q��!�7y�Z#LDMk*�>��. ,�N�,		�T8��`"Z���;��1[| Pt2�*�(���I��O_����2��nڰ`��.�_������d̼K�w�{D��.�?Cl�$��obI5�@�h�©���&#��:����LtXw#ѵ�Y��Zu��<�a l��k����Q1}$U1��ln�M+�F�*d>w�҉[u[si�"�"��5��`�Aw�1�� ����V_�b���؉�b*Ni}	إ�T:lO����Y�( �8y!�z.�]�[�{���ס�a#��0D��&9>&�QTl���#����A�r��Y� �UY��^�|1F*SYg�:��I8�qro#�H]+���Q;3E�?�/��z��4�Z���ֿ��Ј p��r�s.���3���;ϵp#*���x?����9�VȪ�+[@;�X$h���c�@��(������mj��t�q�EcOf��_ڌ���'.�h�GK�k���_(��ɢc�EƊIț��Q� 9f!��_���W����SW���h���|8��hN'�H�LvYVt�o�c�Xo*��s=T��aHO���6��i���-Y��j��Z�.��� h��z��M�I��\ˬLj�9�Nuq�"��B(n��Z�<=��s�1��c"֡n�E��6R�x�_�4���1��R$}ٴ�z��6��&���o�e{�{�,9t�2�x�_q� T�LZi���*i�>�L�^�5YT	19?)�-�{a$Śk8��C0�Dr�g��|M̜���.0��"�2��AWfcP��T�(.#��eR�`$^~�2ا��^�G�W��O{�R�s�g��f�h�������f�Y��0<!�V���R}�6��h�U6�W}L��?�4��C��<!���]{ 3��`�#�se�K5�~u,.7*7����T�x��z��B�(Z��	��	z�������-�`Et��ݍ�{�?����&���`��qA�fh&h����d���6�\�[����o�(�V�*��O^u.t�US����"g�]��w�C���h<���|�E"�~��"�Jd (;x�xO�C�.j_M�(��$�t�,b�S����7�[�d��!�]�]-3Wn�<�A~(9KX�t6ӏ\���s���8�I��T�4��f�{+�7s)��kw5�
���!]��s��o��X���.��'��q�����q�u��� Q(�FEĽ/���7b1~�9�V��x���y'�{0���r����I�l�ӊ�$\�8�̧�1����fy�1��%�
����1�R"*�=9F����pGO
u�yXI�b��r3��S���C��I��'�m�O���	F6Ƒ��=� ���!>� d����]ύQ�E�-�W�_©�T����OZK�;�4�6;���ؗ~H���ѠB�zl�(�_�o�I��� %���X��<N��`�x�S7�݃ΘAA����.��%���i蓛R����E�sw\	�m�.%�j�Е���S+�U�q�+���o8Yj����p��kw/��
����H��f��˜�9�5���s�g�*�t�A��S�3��+D�Y
)�P��$(ЙD�P��R�t�Ýc(x�����	�I�T>?+ǅa~5��S.�TDX�i8������Z��=�/�����pn��U���jH����B��p��S�6�����pt{�j�㊁[3�Mm���$�{F�FH�E������/���6D�Q�+�/���H���vo>���O�2aSζ˶�,�A]1k��*_��]�j0?�7��D@�lvʍ�x�oz�`�����S^.ώf�X����0���_�b1a-Q_vv12]z��98����x�+ӲEW��2�m�����?��m^� o|z=<T+y��������$aǦ��o[V��U��|�����e-!���og�)�a�vsޒ�L���Mr�#�
��p�Sg�M�@�5��?I3�K.@�#����>]��9�{�Ͼ{�S+I	]s����12v�WC[���O>�������$��9���K�~���U���ɰ��Kg���iD.BJ�AY�@�G@(
wC�lCY3g��̏�=E�A��E[�{�XM���G�nq���OG��8�.yg�#̖RN�WTW�iym^��D��S��y�"G\���
�%�7��M����ly~apfm|��$�zT�0��@���,&g�{��;I��m�����'���\ƶ(�Zgf�͠�[U˃n�3E�H�{�,�՞u��z�ߐ�ώ���9�)X8P�5�>�?���� ��;�Wa5��,0
c��^]%�[�?�y��8�2幍2�KpA��F������d53�;ߪ�$ȭ����[q��<�0Kmư�Q�����9J�(���M�Q�8&P<_�[�M/���cT��J��|����^�z݄���먬�F�8ud"%�ɝa5��j'�	8���n�]k!�Z�*� �N��C��7�����.��������n�[�e�Y��J4��]����E�C�=�Ue�!�eϔ߰�)��m���S8����{<{)xq��
Е� ���x;_����^��+z�ɦ�x{��q��֛^�1��/w=�.�`���J�d�M}�*�v����h\�*ը)d�^Wؕ0�CD��PP{H�E/ �w,m���xԵ�Ʊ+��qG���י���U��G�<�}�uqoI?��$h�Mɋs.��%��Ћ@�	��ɴUa���[L`U'j�tE���-�fV�ۢ`7G߀(>�̮�����K�f�ksyHB�Ӆ�)�"�@�~S�\y7�
��+?�S�x�"0�u(+Mi�R5@B:oeB=�{s _���~��L��x���a�]�:����jƯ*�.�g�0��j,ň�Q,lu�B�3k6��\�&S���LD�/$?,x��Gjv��B���xT��ց�oq\�C�T[��^GV��]֟DuO�P}2 �w��'�`�d^-����n��D0��e'f��J��������"�l+�2�vF2��6��(��ҥ��3��bV_�8���c�LG���8�j3
�ה睋)��:��I�tvX�+�8��V�[&��;��I5Vq>p(Rd���y6�dJQ�k�f�/��]���ޤ�fYϞ �L���5%�zx�?><`�0�,�A�Z:O���f�d6:ї��CT���QǞ�(�_r��Q�X����n���!�]2U�Q�оC?H���3��Xc�5h4X���Ë�,�7S���A�C���¹�oΗ��� ӡD��H{��q�ذs�g�F�'k�mF��F�d�ę�ﱚ¸�p�6�=?��v֖���?F�Y�}�yq��$���&`G�<��3�'5�5���}�Mj�J���OP�7��ϒ�8�g�Y�L��sU6FL���x������������ؕa��W����4Q�i{��hfVFmt���4�
�S��ݞr�@ *`>�6�Enw�<�c����x����EO�7xk��T�K%Ū��i�"���ku���1��!�Rܲ�CU=94���*H��'7Q��$BV��F���-�ʲMC|����bR���"~�%О����>r�XOAys�QT(� ���yL�vOK�F�,�!`��X��Y�0M��ϫ�um�p���٩*�))%�Xh�K�!��d��Ŝ`!�*#	�����Q�%A��Q��kG^�m�b`6�l�����"��������&�t�c��t�k�E`a����l�7���Й���¡Q�t�^A ��7x���"X.�E��qLx��߆�3E�;���@�
N�Vc�[37�x ��G�����?I�&s'�Sfw��95����<U�o����h��r��3����Ŝ��>Vƹ3T�V�U��g�t<�$�J2@ǳk�m1K�PU��ܩ�}��|����4ёC%��mpt봐C5լE��9�B��S�@�C	�9ЭB�fܡ���@�R v����=��ȳ� ������@�a�i^�B��H�0�^)2j��{+��0�Aoۓ���n��^$ڍ$�C��0���:�6_�J���ZN��f��9��~�#m�P���Ɍ��H�\%��l�REK��pJ��6Ǫ�G)�?�G+*�K�T�^xː(b[�� [o��j|Z����]L��4�0˽����?��X/wOD� ��ݩ�η�kT�^E�v�j�=��j�������\�&�G��J��u6jA!3:�CL��X�T�E�}�M���� p�m�� �WlQ�%|�r���V��!	H%�|�˽�?��N�,�|�<Z���QUkA
;bⵀ����v���(}�����?���W/���C��� ����Y�;�u �w�Τ!Q�.�;�ӰG1��W����\���w��R[�Ĕw��p���+�7�zU�1�I��O����9|�XP���FdT��	��m�L�Fb&g�z`�7��t,�+�3�T��wb$�|��~��L0R�|4�0�]��M��řj����O(�B�d��Ըs�̑Q)��]v�T#��kG�#C�<�̝�$����� .��>�Y�*��>���~<b�IԳ�=N��X�~����ިX�-Ԛ���BF���9Ҷ�!��dR��.y_�����'T��YSd�y�0@����X��F5O�����U�0��qa*U��������
t�	��pC��P7z/|�W�g�f�C�T�\���)�Tq?���<��OF��q'"��wb�6���\��s����յ�#	<�,�����u@"cY�Hѭ���DY�]�._��0�v��w������	+�������b2s!���[��D�.�2C�T�����'�ҿ�ka���xt���u�Ɍ���VҲ�]O�m~Z�I���o����@\zTr-�r�>�T�Zng~vm�r�?���i|[���&5,3iRŽ��&�\oy��{7ÎRb�L��L��pT�1Dd��m)=?˷��k��������*^U�{��!\���w�66U;�D��6�.���P?�bLQ��=X�Vvȗ�1L���^�Hr�����p*s���)���wZ�| ��]��0��%P#}2�@\7݇�2�����Y�"�o4l=x\A��|�������L ;e/nFk�H�.��}pt,c���l?(�|v>j���kE�:�
N�<��2Ao���Z�
��[H ��$Tg�ڄR0+,��'�>;�?,�mnNY6mΩ��\6�R�t��<Ґki&�e��:�\#"�1O� NʘZ�����g�݇T��qj���Z���@�5#��8.�p�L$�08��^�f�;
��_�_��ݮ32���N$R_�! ���$�:�?t_[Da��������5F�fC����F揍W��ڔRZץ�_p��)���/��~	�o7E?��]l�e�����ۿ��8�v�:��Fs%J����7�t��.K*9��O���a���$Ww��>My-]�w��*4���ɚaȟ��xzڧ��Xk�h�7?>h��4�!��s��z���2DC�Sv%�%C�98W�Sj�?�z�v�7��ǅ+�^�l��E��ړ�� [�\;x����xf���$�L�ɽ�2N|��X�2R�{����h�AL�d�:���fi��{	��n= -��κ��Ӌt��ng�&�:'��Ǉ�H�=��LyǖJ�
AB��@{�1\��\Z���L�)�5��������c&IY�bSqd޶4�����8&2�4���R��'��[�`�Q��-��[B�h:)z���7�2kI���I��lDfN������a�g���Bz�ϒ.~(��A������>�<��d�[�0��aOX�\I3I%��.�6�UGoi�A�A>&S��D��ԭ����:�-C����$j���eC��xϵ�l���:N.�5�{�3#���D���J����o� ��T�32*�&�O*G9I�Z�(gۖ�%�O�A���)p ��!w�G�;��.�`�.�h��o��a����d�#�m�ٚ�u�%۳ɸx���Td#�iw*IΡ�R��\�=~���gO���9����T��c���u䊖�C���� ���O����?x�v�"��\���Շ����LB�� �)%8!�sc]�Q��X�+����Z�x���S��ߒ�T(�9"��7�`�\x�s��P�Z2��!�&b��x�Oz�Z�\el	/m��I�8]���LH�x��_o��G��zW��2�B�V�@�7IU�T��X����j�qu������'�Eyt��3c���_ O�~y[XU�J���$���҅
x�o�xn먷�{��,,�>IJ���hAϒ��1�E��m ��Ћ9�W=E���ZMd�-c�/��a�����Z7a�~O�曆�bGh��dp0o��2`��VD1Aq/eY�*�_y,v�l�F�tR��پc) ��<ּM��Ɲ\�}�C[ـ�X�l�^�������Q�3����d�х�W=:X��k>��-��!�V�@P 2p�eO�٢'ɤ�}Rά�X�*���F����1c*7i��,�n�w͎�X'S�����˘��w�Zث�iY���]&��˔]��a�@�%�F����T�<���g?>�m��﹕���[��O��O(%���5.M��t"m��;�d�#�`�
�9��}�Ƕ�W8��Q��60*�t�\J_Ud&��a/_�OS�3��^gE��F;Z�+�!\�|d)�W��p���@�X}�/fj�;��  ���H�Y�hVT���b_k�vd���/�g���=���%��������&�q{c蜲ld����M���MB���3�ƌ�Ŗ7f��ш8Ǵ� ���A���n�!�����d���sbu���9��Mf�=o]"��m�p�Q��>HX嶉s`k;S}�J� f��� ��8�����B����IM�R3���!���98?���eF��'�U���w�Y���KC">�ؑ����Z�Q=)q3o��P44$�$r/7oQ�̼��.�#�D����e���U�E)X���9����Jlf9KJ�[�#d9�_����b��!������S��B�Qv@�;�
xH�X��?/�Kd���������<0+"�|:fF�]����w)�:jO�CNӟF��n��
���� �0� �?�N\}��'I3�O��Ɉob��u/�������;qA�J��f��|Ep��q�3����_-�-�-�da&�Z{EDJ�x������1�Nq��J+�ұE;|
yh��9�����8w�JR��R��Q�������nc�Y�T��X@pm�W�&�?EivK�Roh��}W�z�&����2W�>��M��*���_���K����	_&��nOH��V.6��!X��S��q�jd�¯��z�Z(��}�#�Ydߌ�����;���=������6OS'¼�2t�/���]�M�C�\�%����}8^�!ׂ��������N�����$����ٶ?���i*!��m��qM�1��1��Q�3;pN0�D«��!�&�էP�$}
�\�p���f�����F
k�\��?T�Q"P�7�&dvu3��=\ւu�"��&���lq�z"�=��'��mX��,#Ց"?s4_&��t!EiG�^|X��&�Z�?�opi�ܝj$��61��3����%B�v���)F��/hJim��|֊+���O&9��z��Кۈ���T
Dԍ��=�Iw��W���Q�cm�d�`�wR��*>Ą[��H�[���F8�����y)h/:E�,�v��`��C�9���g�"����a´�o�9h`�v
�>{��\�2�9!;���3Kh�)����P���<#��5?g!/��PLJ�y�,Kw�������$*�pd�'=8"i��S��z~�5��a1�q�Kc�2 JAd���݉����3����ԅ��y7�ܜ���+����o�_ُ/CZ�I�b�np��l��[����`��8���<��~w,?`�h=&O�S����{_�a�H�B��؂��WO��GM_��1���|eą�5��Il�Eήu�����uyb�>�*�34L�5FbݖZ��KWA�Ӆ�9��gKB�u���,F	h�!�?�q�ЌN2e�*��9�)Ht�bb�m��'��)�s���������W`�M�Y�����]s5��i;x��D�xT�B����	�l�t͔^o����>�A,h���G�O�z<��A��\n�-��ټ/��X���Z�̣ȱ�w6-#W�C�ʓ;�"D��&�)�V6�〉��:L
��#@&Gk�����s}�ϣ��]���7d���d����C�<����Q���^�#v�k�Y෾"x;/�W�)��eΛL���5�zx��!in�
s6TG�)\7M�%�V�V9XK.>] 
���t�`J�Gy�n�3f�@5�MO���y���m��0���>��fR���w �[���O��޽��(-2��sW���2M!ͭ���H�žU���	S��
s��Z-�V0 3�]���"��@���)E&P7���Ͻ��q��7h�I�o�o�ge�Ch��m�I��SO]r�1M0K�c����b�bֳ�fi�(��i���ˀ��᥻1�I;��k��w���q������P`g�Mk��l"ݿ�zQ���]8v�w��c?��U�����ޣ�
\��V(n�aiHPW�-i����%hD(ť�g�\C3pܲ�&�vkR� �<÷�V���%K��E�p0���">����2c�2��&We������Og6	&�v(]�s����r�J��z��������@�����<��1��3��!4�۹�Yu����B�<�sXUl����ҳ�S���9j����e�@.�Ĵp��N��_t"�/r�!�^�U<_0{�B��ԯKy�ۙobc�@�a��6�xЋIzS^J���g��q��$E4�#�9 �`#�[emN]h�g��5?斴V��NA�6�0H�7�a�CV�45�Mq](K̤�hؚ�_sԒ��
�7���K۟���&�1�X'qP|���6ʘ�@���������f=;�쉮��en�D��4'�����Vط\$�	���![U��|\H�Nk�} E9b�6�Y,�LWĈXew?�����{US���AzҴ�z�2��	$ֹe�~����33���6)H2�yW��ĊB�	@|}QS�BF�ɵ��W��W��5}v�V�hӔ�<�ސ�a;ˀ3��cm�3�ؿ�SHq� bu���u�<�;�(��w�Xy����3q��?�K��w���ۨ�T��)������q��U�I��C�!�^	���6�|�7饦���&@_]�!jB).@�'N���c�u�����rhBye8.s]5�W9��]4XMģ�J�Sy$��w�w�Q&��"aE<��:�%�����)'�Y�-xDd$d,3'��B�h��A2s��8δ	�������D���Δ���v��^�_&Gn��(�l���+3���n����OغȆ�Ѩ4�˃��?�"���NM�?�[��LgVp6W5�P�XXE�]|v�ɩ�!D�G��E��B,�N��D^P�jQg�|X���+�Zů�U�����@��S!��47>�D_�����Hko��T�f�̮4=���-�b��p�+�f���B�w�c�P�A>Oۢ_��޽O��}W�6*�#�qDO�{�*!�U�Sڤ�o�ўm�>`�E�����pQ�0O�
�k�b�QBi�9I�ҩ ��q�qTv��uk#0kuЩ{;�!Y,�f�������0Ċ�Nβ�f����ybjQG#`u��|��&�$�P�>+��/a�p����2�^����ݭ�:11w�w�bdsn"�KfG/k�U0����z�x�pَ;f��+(�#��f�d���Bl��-w>�,��Me��M�����_�qpm 7�)j�N
%Clx��%���Z+B� ���ǐ�m�}%[|{>�.U����s��r|���W�.6�*��(x�5A|�|���B�7W�h��8�@&�� �@��X��H7G cۏeiO�}�<;S˭�s�	�MFK��iL�>����.Ӧ�1n:2C��[�#�@ʆ=�Ep���Z��b*f7��g�q��Ro.	�[��řd�d��ങ>�j^^�䑛�=5�ac��P��t��*��cd�̃�ѝ�3�r�lTfd�y�q��	4�����&=z_K����ʎ^�l�>�R�'.Uub\�q�Trl��g���Lx�LW)��
^.C8p>h��2o���Xk���ŝ�C���fx��+�bKg�[C�� ��ǋD��7�5L�H��\?���J��o�����j9���`�gVǦ�y�R4�kR��vCX8]e'��x�Sr�,4k����!L�TU�l�U�{M�I`b�6���Cڴ��'[`���O?&�f&�� ���>�J���/p���Ը����1��J.�>1��r6��������:���0]h���)�J��j�x2�6��rV��䃕;���֎kq��3��`Ul���-�V���p5�U/u@��m}��&��+����]QRh�[使w�j�������5�����!�`�A��%`ʤ��)laa����HEf�{�&ck<�.�r9����f�-%tW���i���Uxpp�_8�Ub���l��m��F��@�����^��������3&�`pu��c�㪉���$�{��]���l�nvE����T���xkTʿ��oZ��B�+�c�݄g�1�؊AP�V<��Y]v>t�T�Bp�q����n`7%�S���bt��n�]e�#����P䆜��%�����ۻ�;���m�M��z��� ����������Z��嘆��+���N�4ʦ'���1K�z��o�y�[�6�����- �pUi;����FŨ���~˚�;����*R�<����W��!F���0����{-P����F�*Fqa�>'+;�WƓ�=Ô̾�[!�7����9�#~��x��IhmM�IuJ:?)�&�������(�Z��p#��qy��:��	H׹ ��H������Q��J�t8d�p�Ԯ2�d�{����l_w1M�Z6�p��4C�j� �eg�1UcG-�DB�1���U�ya�(�=��;���睭�F�w���#���G߂Gw�@2�_�ް�Q�%d�:��#p�� ��)���г�M�����U���Y�Lg�[_��v�9�B��Y�y�Y8�{�K��l�]�͛ж�����`�{4c)�K�rZ߂�י
+���A�'�_ �J��b�i���c�N�:�0Z X��>v5���Φ�\1��SV��p-�V�_����]w=M��-by�56ߩ�ԫ�����<8�f�ۧ��Y�S��6Z��Nt�h���%��i�7S�ń���_.'��g�B#0��ͬ���6|Ο\����w�I8���q��ڒ-U��r�Ҧ*�;����Y�CX6�߼,����3,Aj�m�p����5�r� ����P�3[�Y	.��4�J��5e*�G[�7�^�k��q?V\ 	�d�8�Wi���@���ǩ�Ѹ����P�&xU�#B�?��BX���7b
���B��aG(��eNYt6���_d�sM(k�,_t�e��f6������'R�T�ɤ[�������w�P�B��+O[�~�i^5�.�
${T|�e����߷Y9��d�4(���\�y�"y�X�02����m�S)*S��� �Fvu�YM������U��7�^\��������Ƭ�1ť:����1/��g��[� Z[�!��PWE��� �7UF�����a����*Okӑ���mv���$H_��6�~r��޿K��KG�(�Y�we#Á�Ml�em����;�����������.ٞ�.F� �~���ũ$�4yQ�UH7`��˨|)�Q����P�e��.|R?N�Y�!s�<��xg.<�r:	���-�u���[h�#-���>�0*�q��}o@�7�6�D����d	=ͺ�txJ[���Q<��B<�q��W�*Lg�#��-f� ����'s$�A�E ���gks���o $X�O7N���PBĘɽTy��2��:��1;�Wr��ώj kN���^]�6��g�'�_�[���wKT�Q�We:�� ����_/����R-ץ6�FX=�)Yt�;**�v���T�ڃ�C1���p[���E�R�,F�!�8&M��Zp��p�w�,:gY��8�X�쫌�f�@����2
d��E��	M1EӬ@�	ჭň�(6�����E$X�V�4��׭#�e�`ݓ��	A�� �V��A�B��k�Z.";��&�Q]��)��i�"u��(�_;�b������p9�L�$gl�s����¹GEj�F֧j$?�^z)"2���'"��kI���lI�IB�"�_sb���[�8��~�ȷ�2�V>���_�^J���_��fPWfW>ȊM�~����ez_?U�s��zg�Jn��ȎX?����3N��'d�h��ia��&�{��M���'�G��wKa0�87�UF%b��8+��p�o�zGN�AݎrS��d3ͨT�`X�nG����:1I`����J	�d9�sXp@s�,�i����KT��0�h���m�Ⱦ7u$�����	�B��	T#����������ro��hu���n��?�� �SK<$��#Δ��@0&�"�ۜUⰱ�6�9�\~��hT�u|5a� ����h���'�T�2>QW�H��WY~��H�wȦ1�[��<�pS���c?�%��B(ۼ���s����Tf�h���#vq�F�}�"�b��_Ɣ�_�rx�b�s�����]��c��}�뀏s��b�C8���[Q���@����:�4	����	)5M)�4���u�>k=I���k�Wo��ZÃw7���YE��~@b���]�I�;��{i_j	4�%�?Jc��Uޝ�$fB�`T<9��p���j>�ٯ�E8PW����^LL��)}�6�kV#tx���ݨ���{P�&��Y�ſ1���{߂���T��W}��|��"���sd���J�1��Y��(L�BD���P蹣�y��$%Ģ����d�xy����
�u��Q����29�@H
�9V���K,_qV�N�_$#v*`m`���*�����b��2�L!�� ��6�­��C��=�V�s��c�<����n����-�6,��$.��h+ހ��A	���<�}j�)����Z0�w?r��M��^��W�_�s;٦8��,����E$�[)��X�����,�����<�J����v��l2/|��{H���|���'��_�Q�iO_!�i�q֪N�����Vכ��L�N�~ּ5���-]|�ծL�b���W-rd��hp�,�J����m�y�f�&�HN�i8� ;��T�|��rP��B��܈����등�4j�?��P�DƗ�ԪD~8���P��3�êR/�(���)]񗒳�d��9M=SA���<L@y"�ݟO��M�ێ`�o93U\��=����G�p�n+�c�]���v+6No�d�Ui[��� �
�WX���~s���ܲ����K�O�6��͡����B�k�d`��K}�h j�����+<R�Vn[�����Ͽ�/����7�.Q�E��8D.Keuf@�-���Nߠ�[�^ß�!�z�7N�J�M1N�����'s�c�U3�ǅ��QW8���l+zJfBL숈8��}�L�Mn�fbHQxKRX^�xӚ��������XiD�d}�˫�+Fɼ�bZ��_��	�:����G\uS�zx+�:����Yvv�-
Mʦ?�q]d��q�c��nIC�!��H}��b�A����xY�r����СW�sR5^t[�ʣ��\��,�a�I����CW�䡸5F�x�L4���O�3�A��!�;���-�tr���z0Ci�F9� 5!�)����A�m�|����
�{��F����l.�6'�B�N���	#�d=)ʀ]�.������&!p�=:w��,ֺF�/�&NM��
yHz�0bn2��i��2΍�ik,P8�C��W af>-:	H!$�l�~���CF^V�SC������C����@���l
(=��"�{��I�:���;��f�>'ou �����<����nro���X9�4{Jyn*����-ļ�!�1y�W�`�R�V���H�/�~$kV��\LMf ��]q�R��?�@��~�������� ����n0
Ok�	�����u�9�b;��3�,o��������L��G�b�bC��&��������-���� zewb �G��S�	]@�I��'QV��^�5�Ҟ噭����\A'S0 ���'a�`���UkӜ���3�.��B�r��4۹�����e�����W����Wx��1IG�O�$p�:lή���[n�r��4�i�DU��t�7}�[ �j�Ĺζ�V�Z�����Y�k��eB�W��*��O��ZՔ$Uzq�ߪ�����M:�yٮ�}Ic����|NӢ�.A����L-d��NO��	�EWl<:�s-y�7꫙�#(��J���!���r\�����_�|l�^*�����w���o��|�&��>�d�NXw�SUG�Y�,`�.�A�x��A���,u<8\^H�FD�L��3�����ӷ���I&��𒉫{F�^��"�'�Y�� �#�����R��ɓ,_=�w�ڮE���
����T�ؐ���*�;�qe?�/g끝�^�6 3��l��n����Et:�٩�+�Y� r���b9B�ȗ#�_����7�1�%go�_
�\�f)m`�`)�˫�b#�fc�pl>�EQh��0�.>����p�����������%s�n֚�	�;��:P�.�� #%��mi�Kr�W�7_����w:o/tPU�ir�l�;M rU�+�&l'�]�ą㋺�W��pC� ��s�ė�)r<�s�o����4[�Wn�z��Y#�Z]T\���*��}G���lG�f��	1�H<����?{�<�;��L�G��X6I�!�9��P�@�3�i�E*b��ì�O&��S��p��9�����q���e&+�xM#zw�$��_/ַ��@ 9�@�,Y_*Zvq��	]�)$0=��G��PQ�`���8����-�bcgh�-�ܻٖlQo�}��N"�!���m�1{=?97�e�`�p�D寮(Eʫ�������	�ȱg(C�j�E4P:`V�_e��g���2"�}wY;�R5"zM�W`�e�p��X>���M���n���jq/z9���arI�������	V,�yx8d����r�`r,�w�0q�c�?�|ڦ��+��+��j��߻���SvyT�Ց� �i��ҷ~�!�<��ؚ+�|.�o������yH�m�I��jL��	|�h֌�SU3(.m����~ܞ�t�$�S`s��@)"�Â�K���Ú�kF���/�������>�J�3qè�n	�����:ɗ��Q	�퓐���=��\�� ���,�SwBɵ���SH{�؉�:&�#$��ƻ<��=�Y7E��)[aI������%�<���8ʊO��E��
@�Qtz��3|�;��c�BG�	�b�ӸLF���/��sDsۡ �edG��To��E�Gٙ�Ŧկ�b�`C�]m����a�����j��A���`7�Ê� �]� �6�����Ȭ=�e��0'Q,6eޓQ)q��P+��Ϩ���#�!�@ �EwR�Ye'p�T�h��]�yQܵ�߲�2��q�n2႓���.L�JA�܉6�U.E����{K�S�%I��耬f[he�`�6=�V�T��f����W�0���<?Cq񳰃WXi
�ȫGK�9�.ɬ�^�_�2bA��?�E��j�
�Bj(�x�ma�5�
��ģ�]�ǜ�|�$�A�����,�PW0�?�x�aor�j����g���xղܻ.c��;�=1ÚיŠź�m�!��9
�$b�y�pB$D��QKg�^��2 Y��*���gL�O�f���s^Abꢛ3���'����RHa��Y��)"�DlWwc��,��qt��؋�C�	N�;vx�����:T��]��"S(������t1|!��?��n��]����I��6II �,E��}�!���$�пq%��7�X#�`�+s����F���ଵ�b\N/9��nA��y*.D��+�S����q�<��o=7��� ����
��k�I�FL��&ԍY�׌$���S��m&�5٤�6Ȧ�c!ض�|r�	
i�0���ӃY>�z��xQ%c��
JҮ8�)u��^)��I��mQ&ݎ���
3C��)�Q`*����!;�#���E��D�a��B�ۧ��k׮��s��o�JzC�UƐ�'m�A�vOo�`��߰[Y��x�+�F<j+�Q�����&�q)°'��'��4l߭f�V�M��p� ^�ϨX�>5�F�(Ӷ�RY�(��թ�s��?អA�k��2=�	1,V�t�FY,�Cva��w�ۍ�;��ǀ�[�#�T�L"�&jπC��.� ��訌E��ҧ��}�����#S}o5�p�z,��M��x��� ��*�d�3g�eC1(T��N�x�����ݖ���*�׳���-k[�Q��0�]	����l���,ꯄ��K~�{z���c6�0sd�yݿEc�uW@�Pa%��ޞ~��9m:??n��V#���.X�D��A�?=�*g����:�,��~y4~~��ܴ�W����ۺ���S�~Vl�Y�:$�IC�����NsZ���M:��B�;Q/��Z��d������?�!7��\�Y�֧/�v�\`���b�z6@�t�>+U(�������_��K��*S�X��������S��e�CI"�m��{�����W�AP���r���e���I��X��{���5�!�9����3Z���ټ�ǟ��:�Ea�t�)�h����E�a��� ����q�׍~'O�H(,�fT�.v��R�W�N̈=�}��9�K������jeDv�_�Іa'l8Q�%�ơ�\���di�-gO�� ũ~$�-���ڗ8φ��{�E��M��Q]9<�W}T�1�>�r{��9����;�HY����q�	g��|�C���-�G"�T�]J��}Ѫ�k��b�껵nf�za�
Sq�Z�q_�&�����c��O-)bO0مP���qJ�n�ŝ�CB\^ʜ�����do���U���9_��M��36t�{�[G�MG��-j|?�d{�`}ǟ�ZD����+"zu!�Lb�j��а_�l4��B�8'�L&�����\��3bklYGe��m��Ҡ":��}-�Z�?ʱp1�5z�4��Mo��F��f�-�s9��c.�f�[	��9�P�7�H�,̑q�F�Dxx�W�"!6r\qB���$��F
��}�ⴌ`��B~�_̄�O��|:S³�Ni��Q ���PŹ������޹���.h!�i��q[�v��>��l����kE���ˎΌ�Ϙ=wiP�t l�w���3��b��w����pG�����d/�޺h>A4�p�*�Ga)?�8�P��񎞐t�:=Gg,���-���.�]��a]�8��<`�A�뀍���բ����-n`Bl�<��J]c;�[�~[�R�#Ȳ��Y͒!g�s�� ���~��h4Mշg�>6��F�d �:��3n�>��b��0�rE3 ���DX�c�в9c��]��*�2��X�8����/�	me�
+n ��p��W�X�-��	t[��ӭ=��Te��g�U�2H�1;e������B�[S��c���'��k�r����T4|zB|U�v�&���r!�6�ؕ�*�mm�B��G!�/$�>@�,mO�i�W�����h�~��� 02�*hËV�`���p#�I�
9/��di�81�9�&=j ���2��Ly�Q�e����΀f���c	y��I�!25eV@0�Fo�N�� �SЫ��u�4����ob���1��wt�,�N��td����u�ϝj��l�rx��f����֏����Tv{a]^�Y�f��{ Ź�[�q�e�ڥ��[�Jӈ��D���������[V�u����-'T��ᜢ�5����6��1�4([(���^���ٺ�)<����\WUg�*��-1���Mv�"�ۆ�E냺 	m�:/���Ge����})C 2�N�!B�C.�s/�E��o	��:���cF.:�N��q9�G+���e���j�k���!��RSn�-�����'�F�w7���k+g`"m�]xG?!�]6�Z,/��$�e�����׆ p`��XϭȦ��� �+��2v%���L�Zu�PM<�N�\�	cn_GO�������b���^��3��-v͐+��[еѪ��������
1�9e�ĥl�9�K����/_��=M�} �~x�.򈁙Z�7���HCm��G:��Y��hm�>�P�,���ԕ�����NX8�߽܁"wUv�w'A_^��$O�1@I%.�3���c9L�r����SM��C�mRk%�0atWW�T�p#�������1���	��J��9�����CN�����Ӎ�������\ٶ��Pq��K�_�)B>6�� �p�a�p�_�ۣ�S��$����$��_*�P�1� �ҽ[yJ]�ԕSW�a��D�	������@�ʷe���YIF�[:�����'>�-o-a��p����hT�;5�����$�v��8�}]���/�� E֘@���{T}�a�*��	Y,�+�ÓnϿ�`Iq� D�ir>ķv�:f��+b��mނ�$�4�K�ڨ�DU^5��_�BR���	�I$G�p��xk끡_i�y;0�#�@��h&����
��?	{�9��g��έ���,^�Gk"p��ě l7K�c�3�|D�.��@p��ױ�D���J�{�qܝ��Mi�0�d�
� ~F�	�|F}���6��ׂ�[O��v%�{|���X��v;sY�L�bi��$ڍ)�(c=@+��5���-�3؎JO��	B�Q����wZ�C� f��2��}R�a��K���g>O>��mv}(����SR�3Z�+@s�9��r�ʻO0�2[D{7�2��C,\͇m�,[��&>J9�}I��^�����8��ڂ1t)`�$˦��=�0^�_��(�ulCB�,dj}�G[�ו_�(]���
�&�!~�����Z�A�]JG�^��8M�h�rD�� �!�Ugx%�qC�TgAT�*��@ɮ@�`�d���R�LNC�i-��5!ټ�2ݭ\�0{2Л�2>�Kce�$�埄��p%r.�� �1;��c�&����\ر����	�&]P�qt��������2d@�=Zsւ�ʒS�����Y@�-���x�J�K����E�̺G}1��uO`à�,j���Pگ�XP�=\'Yz��n
$vP\��g�0KI��4�0z뀩,��5);�_gGX��\�q�f2�-V��:ե��κ)bp�Ѻ����S9[tǈ:����%�2^V����J��|�����l�2�W+NE�*�L'�8���0��\s��,���-89�˾9����8(�{Q�lm��n�ո����؝�����m��D��lr-���t4&h�U5SZ�i����ҟV_3T��Ow!#v` ��t\��W�K�
Q� Ba��qR"�ZK�1��P�Z�Œ^Y���ɯ}���r�dR�F�,[�-�b5Ex���)��ˇ�C '�g�Ƚ���<|���	�'<z}�*�/;�mj�`�VG�O{M(�5yC�����b�Y���d^Z� 7�� ��>{<Dx�˝��Qf�҅����^�q�c��Ҍ��B�{�X�0/zyn��%��JE�;��\��������'2�����95��c�G����hd�s�����t�e�f�4KU}�`O��ک�X;�خX&Ы?�K"OB�x��Kg�Xǌ��'*����J0*�;�J<)�īբ�jhK�F촂�sM���g ��[�b��w�޸}�b�	��8�A.qֶr��.�f���fBǫ�c��󋾰=���f*ܺ�Vh�=9(_���U)�P��q��"NJ b� %w��^tIn3|�}ȾD�͂�.޵�&�H��RA3I��H
H� ����=<���9tC�c:ؤK����9(J8���}�~h��0���+����J��C�u>"���`g�������B�[�<SAJ��*Up��Y�4?;��U��h�B�% ��B��Nl�Mf��C�qo���U"0�)yO3�(� �C�|w}v�\v��e���5R�t�i��M��#S84+��7�ShڪO�ȉ7�����r�Rj���� ��k�w0�ZB��hl�2٠ ~0���-c�%�$��[W�8:�H|k��y>q9�$����!�a,��L���ɍn�
��~ٖ�����0�d~��Ͳ}kPz^H`�Uv0v)�1�p��  �j�)���}�%��T�	s�MT�?��gA9�Q)fr:^�b	�B9�:�^8�\�hC茲��lF�O퀿N�;&G-g�W�Z��q�&Ut�W�r�Τ@�[�ɰ�U5�$�aBH���w�U�﬛��֖V���hBL�	+X/D�� �3s=�n����eg�Z��Qd �ә����wKVp���9��k�${E k�q�j�x�Mdʞ��Мkֻ�K�p���,��V�7.�<�u���R�K��%T�g�������D"����IM)C	<����~��tj �ݩ~;�8ZZǮ[�`o�����5Gr��ۖ��Q0��l'sa$��u�v��q~�����ĔΣ��5���j[�P(L�w��;�)0K��{bauv;�M\�p����jI���WtS�^dԽD��$�vB�&f���_/UzK�,n07O�����}�]uG�<f��H�\JJ�����0f��C�����< �:�.&�Q2�iNB�4��s�n�7��� ��8��M�����Ԩ���=�cOF%�c��K�����5�Y[V��^Ay4f�c6�����Q<�=@`�Z��U2��?�ȫ=Z���~�IT{�ui]�[�D�m{=g���d�10����Iˬ_}X���5�HP�b!ٚYlӵ?��6{|�ݸ�) ��	8Cg|��Q8�a=�^
p��¨.o���u��m� f�ה()K�j�ii�?#
����F%7�G0�~��,��2�B�j��+Mĳ�Ҍ�����߷��R3�j}(������+�Q���ٰ�h&��]Нz�zr� �(�"v1�������6ɪ4,��;�;�ꥶk�P����c���q���>�0����%�M�c�U���f�6���q�쪵[		?�Ծ�����NU��.��z�1�1@o��(��i8��Q9��}��V��#�g�fcKd7�_Ύ	��l0r�X���g��)�bI6���6'Pj��6<;�͍�8>/��;�����o�����j���M�wo��P%�Ƙp�~S�;��nh�&���ac&dP��0	E��f/˧��w��P,����Ǌ��c�3�Q�~�����+���(M�9�k�4�U5($�b�-�2� ��1�����ǋfF׮dz����a$x������ܲg����Ȁy+v���E�� k�}�������j�z<M�b�{h6R�C�(x�[��vF�\�ޜ �>�0�6����E>�������Zg��*���wW����=��#�m n�1���M1#֏� ������rը(�K��[����d�"у9�@�4��\�ϕ�sL�\&�aV\�ό*=���<g׊��S5_D�7�Cǡ�$�]5��@?�1=���2E��-�ƭ��"E�Z�|>#& ����|w��-JR��\��q�\�[
,�ܘP���S����=@��(Gg�O9���6��&7�ݿ�Ks��%�~�������0�u��2�����7#��m(?r��F�)k�� M��z��Xth�|m8*�z��� _a,8�+�f����7ut@:x�vy�ѡ��}U�=��V Rx'ni�c�"��G�>A�J���a���CS�0׬��(��[�#H�dQ�r����I��\�/�+?�Q*y[Yw'4�e��r���r��>�Z��P�:��sP�1lJ�c�a$8q�r�"�s�ϾO ���7��9��hN��IU׾�kL`2�7ʂ���Wa"e/���4��.����׾o6�F�1��8�XF?�\�2��֚���،�'��͉�-��7E����WjӮ���g�$��.{aʧ��.?s����.��MI���<dU�W�E�F:�9:S�6�TF傐z�-6@��%����Ʃi���ȶa�5�|��˳טj��꿠�*�������$��r���ꖄd�?�uQX���iq�����4Z�g8��[��72F��gȢ�^j�β�H��w���U6,�K�}���Y��n�Ш����J%�j�p�فz�\O�c��;+�21�[�ʪl7���]���0[�����}~H��MnBQ�<L4���=Q>�d�V�,����46�Q�1�{�(��މB{TrW�����&LҞ�q*y�9�M���Gn&+�ɦ;����,e��������v�j������0��'~p�
t�JQ�^P��Y�Wr�΁�Ϟ��~c��5H��AÅZ�'����pR��n�$�k,�瑢KK�9���8��;{�Z��%P��t-�ȴ$���ӓ�z�O���ަ�PC�Jc��W��G,��bes�P�ݙ�Z�
�V����:��w~��?�_it`r��w��)ݸ��$��e�&��ŋ���:���q��_4�V,v{� )�>}����q����gO��K��e���������	�4�t�چ�4��,H�.:�8�]H'�_h��6"���հ�m�+��}?�r0��4���´ �W���|�⮫F���$��k�q4�m��q���Ŗ��8�=�M��#��2��&��MD��>0����7\�}��Ҭ�{Ԫ�3�҃%,��a>uat�݅�}�x�r��E氕���,R���pܠ��K�/K<g2�u�J��IBj���΅�w~�^�?�>^L��zZj�=|�V�	mu}�&��~��#KiE�/HΡ�F��\6���v9�<�ĥJQj��_�� �7�IB�ZX9�➪l6ӝ���9�,~�����9ft櫀���\��`F8̒r��ރ�� ���ʙ���5)�?�A�h�8*�U����E�S��N9�o�z|)�d�£�w��y�r]����&�Q���,u�u�(��ai��!��1v�Ob�����B#t?��C=&gQT�]��*�&(���U�|Q'�
M8�ķ �X�;��1�g��������ˠ���i�=�����m_�z	�;u���[�퓧���`T���#�S�E��o�����亃�&p�>l�'��>�d��R˩�'��̞�J�4[�L\��7�HYj+���-QiN_z�f>�d(�����D��6���q0���4IT�ԙؽ�^�������¤��F��z�1o6�Rn��j\�x�	�u`e�ee���ZG��I��u�2���oBR�9��k�����۟4w�Ɔ��nH"gX��se�|ƕ'�z����c�m~�S9U�r[�D�	�B�d[E,�G�Ezp�V_��w���m���%��ld�+v��Љ�fx������ݐ��!��Dx�M��Ro�����
ؔY���sw��"߉V�R��2�^r傠�򍶰�Q+�T<�|*8@,,��O#N���jYR>��^�I�A�QY꿨�8&�lfxL�J����h��]�c|�3L����Lpy3{N��G
��j� �#$��X�>A	���'�2��o���~+�������-0�8�!s��s�M�z8]<�����uG0p2��BIS�lW2��?O�c�W�%S+9���X�\9E�NV�.�yBy�6}��Yg�[W����`2`5|�+�����7�oF��U�Oȸ��%8JI�M�g؄͚�vP(��{rkζ��|q`H�ܦ>���"7:Ŏ�U���Xb��`����I����=�����8o�e��9�05`q1@��W���9�AZ�Iя��+�a����WYP5�s5�`Ch�c�k�*%yF�5gѧ`��[�A�x����Nx����bd��b`B�)W��g���kE'ٟ�[�� ���_�E%�-��`�D�s+*{|��^h0jy3��&>���h�9Ǜ���/�����X8���ܠ�c�`u��md.[����?���#qQ��V�@m�q��!���(E�]�8�F�=�R�EC��� h<�����I�"�)7����O�����zjv=��jU_�cPt��oIWJ 8G!Q2T^�p$F��3Y�a�	�lJ��R�=@��й��9���Y�KM�GSM��}�1�q5��k�v������G4���a � -����A����tY\^"�V�0���9������w( @�]�t�X9�S 3cÅf�M��8>8 ���]��)�u%�s�S݊aǙ�5i�M��=��%�{�Y�M�eN�"��Հ�X D7�����f��@*ܯZ��Γtت5%���'�W�����n��v)�Li5���%���V��l�����n�i�l>�V�[��k,�{����XM&iI{��C��o�WM����=<ee������W��u�v�s�9b#SZ}��^(�pN�*��| ��#X�ۑ#x����'�����z����<��b�X�]�jׇZ<��� ��Q��׎<O�@x�=H�=I���Sd!�%'��]�2QÓ"�)�ob1����φ_ȟ���q�b���im��T��"OH��q����j��52���B�X��AF�ܩ2��$)y?�s�f�7Ӷ� ,o�U���ao�����G9���c[J���r��W�<���?�'�ȯZ�S���_�`AcL���L�h9�}�N�[��a�|:�`��iI�4�Wꖓ�:��:ǻ@W}�����n��a©'%�!竲�p~#쇻FA �A���}�~��L��J�Xr��t5�{���z�teCk㝎�4h�c��E�A���~?�;�d��_�.��]��;lys?�	T&L�N7��>0���{�tT��)g���\���C���.u�@��a���ڿ.��̤�0��KY[�`�l���S�L�Lo#`�8_�,�����g9{	�!��誆��W�*����u(d����{Lav"����N����2Q��F���p��̀�nQ��;�5W�]�<U� 'm�6Ğ��� :F;n���5�l��k�J�\��x't`�A�ɧ�>��f�B��sjr5�2R1�r�i�ME&�T�D)�>���$���jg���F��iv5��zC�_8��%���(e)NUs�,�����Xʎ�˞}{^G$��J.om�ܿ�A���մ)���T��*�߄�Lc;�-�H�v��3V�aN������?3���������m��Y=Uw�� � ��}����f4��MV����zh!9Q��@Yٗ��� X[�$�Y�+Pq���;���꘹.{�����P�k�OTB�pqM&��5r��I6
#�o#w�V��K�O�G�s�����$����Ѥ����}��	��a�Tp������N�	��wS\�9���蕇)R�:�h+"���+����B�bV��}�����ݖT�4\�1K�&����hԮ_���H��&��M�����G�]Q�$�`�ܪ�� :\��ԭ5��tќE��m"��lLF����:�#zp�r35ʶg��#�]�'��k�2��@�a�ʖ[ٙmh�v��h/"T��M��}~|��J֓6�8��;8��S�0r�{����o���có�8�G��V4p�M���O����X́e�<�x���j���l}�$����ȿ�������nn����4׽��?��_(!��&�ӜE�e�M)�J�yd������� �j"C	-j�g?�ؤ�70�Ň��b$�xy %������.N�-�߀i�k*���USipF�ع���23�����^յ�2�`K���<���C�r^)��A�r��V����>�J���f�u��gۀ��u�.�s��m ��r߳��hL 7;�ȟ��:Z��lƲIa���&�G/ݮ/Ӻ�ȥ? ��v��|�$(if�	辂m�|G<�w(9���y�Xƈ�U���v'����|�����q�	9����|��x*�AxНh<�ehsiB������}QA�u�_�~l����j\������Z$LM`��5,��l����G_}��L�G&��,����_?4�0�#/i�,�eUJ%s_/��ڪM�Cζ��3=��&�_�LaCy�Y\�a�xB����pq}d�|^�V�}d5��=vB�h�0��0+a7·i�Cm�fH-}M�w�z=jw�؞��U���O<��II�d7L9�;��&1a�-�����+�	�I�jj,��-u�jKO���{@���&�=�F�nE�X�N45 i+2Frn
�7����#dL�v�Fn��,v�g��v�CN�!7*/�Ewx�\��B%��I%�]Cn<��,_Bu�N�ad&���͖(Ek*G�+@�G�B����sҐ����=V��A��؇�^��� t.��I�����:�@u �l���c��;DB�
��q\��Q�O�+Y|o�F] �m1���K֔�{�d8�2e'�� ��E~+����G���R@M~���Ai�Z��{�b~�a9@[�Osa����%zL�I�6��+u:	G�I�1"�Vk{*;0(r-9��X<������������\qp���<�Y)������i򠙚H�>թ+F��;�⫺�3Qr�u$.\�������?�#�?��#�b+���K'�2T��y�fP*}���
����43�`��hR�W��n-/9�?5��ho��"�z��t��Ӵ^�_U@�d�\:j��עY�y:"�X���Y�Vu�AײR{"�JB��2�׹�C?�� ̂�%�� �{���梁��cAK��P�OU3���T�r�h�r�-�,M ��;$ɬQ��«�bJ�E�!��U ο5ʦ��م�$4�.=2�N�w�\M�:�x�8��7�?F����1(�C����l�ĥ� ����w�-��������)&��!�T�YG�����
��5�cƙQ� �4�r�7�qmjIk�m�����n/����T�b.yevٲX�S$�G�˧<M/�y����>�<���&�ȘK�M�Qٶ�U$M@�a@�=GDj�a�P�_8V��~�5B��{e,j�P�q���WH�h!s�i6?甘�
�p~]�R���)���Ox�������Y퀜��d��a*��I��)W@�~�[�G�Z�H67�63�`��� �upé�i'r��� v�f7�l���;;�a�7�u8/s�ʅ�c�n�Y�ñF��$P����a@�#���X�~���Mu�
J��Dn̄I�g=�Ŧ����é�a2Ȣ�G��K�`�~ӿ#�{W�|�����t��(��F�d��V�r�7T�w�.�iq�=E�(|!��J?CS>d`����`�Ğ��I���=��q���C�8�(*���~��o
�(����K�x��Ы���&��"`��4�0�MOEN����EO琇S��O�EH�s�uDM0id+m��E�7]|>��Q4�Ed/��fΚ��+��f��&	�1���֢�.�~n�gs����It�9Q�pp׎��sHLM�����`y9�3�ʈ�������'p)2���N ��zq�.�	�
6��yjP���$я����B��2���r�HV�Ȫ?�1C��w"+�1Q�4��� R��I��H�T���|P�6זϿ����P��K5gn�q�T/��p���PS|>�U:�5�X]V� �DHȃa���) �2݂U7�Ж�$�!�j���0̲;hs�@���˽�̛ԏ=����P�O>�����z'�{#N����h�����:-�K�mѷ��@W��]��Ik�6)d�F	�9g҅�)�`g���g����̯co�a�U k��c�4k���0�4?.U<�}�RfY!����4+�6{-�{�5xl�m, O �~h���T�.��7�F�l����j���pf˄h�`�:�`���Qe�+�,�X� lR3�yTEi�Ռ����Ccn&�� �q1*�%��=��6�f^p]�,&e��wiT�c��ڴ��%z
-��
!�27���D�k]��W>v?
+�'Je|�v������;e���E<�')��`�>/�
4�����}�����f�i),��$Ś��_���q~e�Z�m�-#����'���/A�
��pP�P�g�]hU
s+��"C�8�j�B��|I� �ǡ�wd�z�I>:���|jMQT2>c�
�K=�j��a��_1�p%�`�a;���]�ǳ�?�VGK \a��L-�غ���}�!�����'�Bx���X���T �ҕ4e:��}3��D�v^�O-�Hĝrày2�Б �}93f���cUФ�߃Ҷ�W�˞��M��st4ϊ�}��@�7�4� �J�x�8OL���2��6X��k�;�ѝ~��=��������@[�_T(P���_�����e�0_[�C"���J�?�gg݌þ[�<��Dk����y�GM��@u�p����4��,��Y�f�4`	��{X��'&�g���'�W\�_o�)��Q$ઐ�b|�y����h�-�h�O�܂ٕ"�p���Ghq2�E�jy-�;V̘~�{�s0�pJr�ߨSv-3]�CY��Kn��t�J�1�޻�>I�x;�	��L�-0�Vb����Lȃ !�[o�RA?��Ls4V�Gb�3�y�MBq�m�����A"�D!�+�P�Y/nL���vL��0���p]$��t�������4��Zj�&��&qa�6�%`���H�>�Nz#�Gא����Ub��iIC�ހ_ZLx�?���b��v��a�L��b�]��p��D(��J�j��w��D�+$e@�S���O�7./Kh�[�T�ƺ�I;l�Q�����4��*̑K@	26{s<��C7e>���I����Χ�����I\ �.K�^�Ȼ����xc��Q#:�`0��f.q䃆�H?�S&��(B��9�	r��2yҊ���uCɬ�c�HG������s�ۼ�O�^�^�P��)ϑ8K��R�Կ,�=���؅+�XV{s& -�"lG9S@��mP��j՜ؑ�5ye�/��vg�V8i��F6R����k��Z�'��i�e�&�Da����8=�E��+�����s��ގj��g�p�g\l�[i]�2�I��r��r�^߄�u����MU鮊p�U�����٘�&͑��pA� �S��DV�Kʥ��p�|���T;[��K�=jG�*-9�e��5��8o_�,|ݩ[��ز�|�A�{��1Cv��h�g�I[�0`@D��g���i��jO�ŝ��O���ޑ�%�IJ� q@d��_*m����0=�S)��CV&���8cȓ��b''�R�W����TBV�O��d:ʢ������s�@m��~���}f~nW�H��j8T��]��)���uY�g9:�O����]��O��i��3��5��Ӛe;�i����:��7�6d+�0K�c2� $���z-	��(�{=��۹jPz�1h��*��נ(�޴m�P���zX����}����%�2�f�
p�\�3�_�m���:�7'񊘱3!*�H��U��3�Os�h�+��7�:L�3J�\��f��N�Y�0�-�m�<�ZԜm����i5e�
+OP�(�¢޾���'�e��9�_�+��%��z�IW����Ɗs�{��jxC���ڶE�@�]&^�9�C7��'����W�D���v(@�F������̚��u�P�,�O�f����u42�}7,����Y�B�e�Ӝ�	}/40�4+�q#a�@Pw��gU���p�i�p��+!�aj����9���I�řިB���ZqD��y��bZC*�����T�G��u>��?����Z����lz�ݧ�"��<5�W����v�%X�'`+x?��R��ѓ� ^��^̛���!Dz��XZ�]��QF,��(��$}MOg�����h! �Y�-�e]|���Y͖jn�_��qC��7�o�/OJ�L�3NL����!�����V��
�򿸔1L�x���5�wj+4%WU�暑@�<-��ڏ��b�5���m�ICm��i��me�ܗ�QxT+<)�X��W� ��(�#�_�W�+B��f��Q�UT�Q?�D�?6x�|a{��jښ~�J�Į��N�Cq�mj����J��Mu�,Zq��-����n~�t���%:9O���o}�3���<�c��DjnL���E�I����B���8h��?�|w)����#r�f�����dW�*Gz�>�aq��~�y�|�&Uf��ԏI}�N�f�6d#���H/hC�V� E��*@�r����?*_'�i��AhWTZ��#����`��v����Y���!�h#S"~s{#�<ڼ���쎗�^W��q��;���ep;)���c|xԞ+�j�
)C?�6+ �*~$����-�h1�j�ZZ1�Aӯt!-Y�.'�gg��1�fȮtι�Iڒ�%�}�DӾ�~�]�q{��Һ��g=�ߌ��2]�v�_+�	 G:���bZ����A�����k�����;,ϭK��)�q_�`�Lo�'o�]�T�ɐ5ozԲL����M�i٪��o&M�m�GK��w ���ph��v��WH��|_��2z���F[�/@��l�qι�V�?�Ս�{�A���3b�Q<׾wch粢?\-�	JS6�G�&1ԃ=Hqo7-���n�ɲ��-�*�㲳/�K@�rpd�X� }���:���l�s-��	���h9���!����}(U`��_���t�/��Ю`�B��d�p��!t��6�k\npG�z)�D�Y]!=E,vJ]��%��F��$ux�m�ݻ�ۏ#>��V8��@/:�k؈�!.N���m�Abq�j��Γ�9�Bx$�\�3���}hV�2���H��� q��'53/�e�`#�,>�E@�o��\ �ᴾ����M��O�h��{m\�3��q����Pyd-9Ya�-�&xsP�+�l��1l:6�mLq~1%��KE�,�-=�"Ǌq�g�Y�,b�žc��aq1ȹd�*a��2� ��؊��̋�][�"�׍f��(��eI)`�I|a�} lU�*��3��j�޷�C�0(˺aY.�ΐRGi��;+G>���T�6|�#�o~lt��~�|��]H9Q��מbR:VH��S.uT�t�/�kI�a�'|c^ݨ�s��9���,	��_��8�C�ң�p$�����ٮ��a�5	)}�퉒Ц��2�	��e�@Oj�yӢ���ð��wU:�\	u�u������	J����a�M�F��Fr����+�,�L�/؟{���d�$U�
p|���ٙ��"w#�c��xB�nw�ѯ�l烗=��̳��������X� ���-
 e�e��Q�G~�zT�O��e��Z���Й�?��ϔ��s��6���o���I�2�eSB�WN6��z�|���3vx3�H��M��2��T9M ��5�O|�G�i	�.zD���ʃ����IW��T*����mo�Q���v��2٤jVv�2����cFC��bK���z�9����j��E�J��G�;�L��8��9�]Av�Hs ٭~�ޒ�_�	�
X��n]���sY+��JEW�=���/��{3��e���݈;+��dfi�����?Šdl⏏:��N̈g�@.�P�XC~,�ՔO��_�D>����h��s/�]k~��eD��շߙ&�&v���'�H�"�?�mZSI��V�����P��Z�[݇KY�]hMq�1�rQ%_ŬR��qE��0��P'�h���8�������z�c�&�+�Q����X�GǛT8�&��ۑ|Bo �����k��t�Tr�5�>W��8
�����5�P�u���(5a�	�i�Ö��9%�@%��,`Աh��%s,�JBT�����ȯH~d��hj+QK�q�DV���Np�J�C٬��4��|�v�٢�Y��X�gڧ�����g�N��6�����=�k�Z� �˓���DF����±&P��21R�q���V�Uɻ<���S+�3%Ǉ">��K�����I�f	���
è*�ws��C��<�h�?�W��~�}}�Zf��^:k�N1p�N�y'X�H�X$�N���C���ے^s�R������y ��P5�O-�DwVg~#�+"ԯF��K� !02��>~k���օo�d4
*�Щ��4L(�Ji.a7���Ƞ��j�r<?0���oq�fl�VlI�W��/�ڎ�����c^P{���#@�{�}�2�kib}�����嘼a"�����YG ���/)Y �s��"��<���:�!O;����v�e2��1B��[�N�H�z����)|�e��ٱ�~��g��ASf5����U��Lw^��B�C~u@wP&�`!���pY�iaRć	��	a_�śN�ի�"x�m�����8��FbE�0�n��8��d$�B�NT��ٍW�E���n�|�9�.I�Gw`�8�M0�V� > �0Ž�p�!�%��, �6�-/����I�U�w���He�o�F�/�o��c�ѳ>�YH�|Ԑ��E.�V2��cg}8�-��1%iC�����A�mdY��k�*h����p�g5��
*f1l. �U�cOO��-����s��y�U�\�z	�xʋ�> ˾��D���B�F�#AU%4���X��h\����0���JZ�!&���/�L��f萢R��,/f�W���t�����#Jv���_�F�~`3Q9�UuiL���Vv�����"mrݰs�c끱42��vwȱ, ̈h��8��Qzil(��ޒW��`���A�W|m�{��H��ᴙF*��:����I0.����jʇ���\q�-��<1z��yT5jv|mȈ�L������L�y��,<�3�{[�-�&2}88:�Z� �U�82(kC���N�P��u�{Ƿ-d�s�T?i�d�h�QfKUT�E�Q�:����r���7��9�hn����}귮�_�R��o���֯3s3�/����٦���Ɖ��ƻ��p7X��kq�UI��Z����0ɯ2���ΌL�Y�hi�PT�G�����%�9�rӗ	��%�ꇰ�L�0D�=J��+��橿���v�j������I�֒r��v��H+��&<V<���*̘7S#-G������ �O9M�f�H�|�������6`�2�Ţ��Q4�r5�ӭ�0��R��8f�1���	'�d��#�&�~:�3&
P�ӟ4dZ�Й�%�(:˙b��J{|n{	�W���"�N�1���G��NC����U�"|hL���; ���_��]Xy	��r�&��c�w�� E.�N��O���S;����Z��W|�@פc�j�K"��3;5�ߌ���Nx�C�s��N�[5ab�3�ح#=��T�@E�G�C�A���8��(yj�}?u4���s���Dfc�?��"���"'���T���-�6h������Z���Nj��@�Pጉ�5�gp1��F�5T��o���=е�J�ɭ�k@w�Ɍ=��M�^��tj*�$�\67t�8��o?��yT=<��Wm�ԍM�S����LIݷ�5�!�H�|jO�0`���N'qsv��0J�zb�9�Kt�(�U��M��(kD�`)�o1M`u�!�H�X<�>*:��ȝ@���6�Ds�(;e�,"Yu]�ɍ+�"aj�l��KY�
��0���TJ�e'��&����AM82q[^3ugNj�BYL���j�q�k�lu^��@���WH� �．�?�ކ67E�e\�i�
�� e��U��YH������DX������1�*.�J����N�̊&��Y�������
ה�`o�����Z�^Y;�j}�r�G�ʯ�#���1���>�(�g��;@�8z�([�[~�d�7�<�7,Q-��7�sk��4t�A� M5On@��Z�w���=}�-ں��-����G�t����_��+)�"�nl�\�m��&��ѡ�#��m�dUi��/��@�>���!�v^\��c/0��.1(�٘$����EX:G���%������ρ}ʗ񛖞��YB��AM�����#�vs���2Y���ZⷹD���^č%{��&�V����#r�?�]83>!�h��IK|�+m5=�GO�R����r3�V 0`��D�ӓ3�!ht��X�)��>;�����z�-wBƞH*�	��?O�����e�Mc�B�E.��S^èm0�����k)`��o�E�G����s=?;`�"˲my�4Rg�{БJ��u��7J!Kk ��'��������a��D�9<�믭���Ϳ���>�<&t�C��|��D?�D4:R^��[X�M"lf�{ZI�����_0l?d��g��x��^�O>L�m�Eo�+�}x�-���G�Naʀ�@�����y��[�KTE�C�_
�0�i}XMIƭ��4�����;�;W"����b�IH������=�FOM!�j`Q��+s�9$��	A�(��'
�b�N����@q���^�c�3�B�8��+!���;���_m��+R��ս����#r'Y�Bm�dX�P���\��H�Bw� 6� �ȼo-�d�������w��h�H����A����Q!���V�
�D"lfR��o�pK�~S�����؏EY�F���dxƄ%E�Ѷ����Sj��n���[�,{��?������ï7��R�eڏj��aB�iG�M�v�uPl�;Gv�$
�G���|*݀3�o �.����� �@;��?F��'��<�gV�R3��mu˺�s��/��`�[��1���!dҾ*��{촆��P�)~��)n�h�Sn#lk*{��r4���E#:��>��A&&��a�@P2��Uo����v�q������?���b��k�������j�5���{}�RF?����
�Z�T���ԝ�W��MOy��N��
��V�WM9�1�N:7�7���D�w9
B$��1no{���E�)70��������c��"�b:��M�͹I7��',;c�9�׻Jʣ��}��Z��l~������8���B�DR^���m2�3
\����
�3�["-3I8�h�x;w�����Q��hg�+xB$����\��C�����#�Jh�s������SvfU!~=�)�8n��f��Z���n�/�]�6E�p4��S �3�e�P1v����Cһ������W� Qê�B�`����2�M�� ���);}w���adW�;��+�s|wvC�*.Q���s�v�I7
ɡf�J�ɻ���;�OL���6�\���t�sӓ�����(�큑�j�NRJv��9���L�.���H�k���K�Ax�A����m�0C����Ǹ��o;�4��|��fN�s.��x�'�^[J�q�i���=_��,P�[�#X�a<��nY�����jD��N�?���:��>�x��T�����o���&Rݤ�C��38�P�b*�`ϼob�P>TDw*o�m����y �2<R
{��Q)W.@�\��]u]��$�LH�A�OX��̩c��Ö6*��P���Le$R�-k�4_3^#Ń��)!۷x�6:�<�h�*m=�P6ߚ@ו���Z�X?a0<f����9��7���)�y:r���c��9�A� ~�JnQw���-��_3>��me���~��S����ؼ�r*�=�B��n@��<×D�pF�ie|#�VS԰5��B�AO�$/�Ӎ+uT����h9�83�?�C��e��k.�ᐿ��f�&��s�o6ʉ�_�î)*\
+Z����Ɨf�3���G'0�%)锒���!>AB����+�k�;;$)�r��@��5�yr�>]�dE
h���#���Hb�+TG��{��c��)/y��P�"�t���n/�v��l]@)+I�D$P*$�sW4 f�/ЇO�ȦT/d.}�R�H�]@�
VPB�K5��A�|D�2l]u�W�E�P���B;��cd��t+&�_OnF�����~�/��x?ӗ՚�UQ�E(�k�4ϭ��f�f!Yb��ϽUo�~t%�Npx�f���2ܾ�����.�~/��p�f ��rS|5�lB����U/���oVj&�w�ʣ7.^�N��'��m���l/����Q�C¸����a��������n{�G��Oc�k�r7��V���9^�J�H	}Xq�XBJ��Sħ3�V ��n`WCaK�4�.P��*bxJ�ZG���u�q��vgR9��dݦ�_}"������q�|��́;V�qh�Vz�)���"Bm�+�bEud��\ 	���z���>��W� ��P��n��٣*N����|q�@��j�Лɝ�7#KA�F�D1��OĹ��cu$	��IrX%Q��.�B��<p���[��NMPٕ&44�(�XOb	�:�u�;2��;�D����0l͒����Ə�G������G\A�_��|�Sp�^)��
˱��-�_��t��Q�eU�^�1�ls<��������LT�L�v�]�=J�����V�;��]�C)n}��rPL(J�D���E�U�����ٕ'KP;�!�+��F��P�	Śu��`M:{�fd����G�[��z���a���?d�5�x�=+e۽ʤ��H��D�׽�؄/I�ŊY;��k v�'f��jE'�޵-`�Y$�ݦr��M��Q�ix�i�3������;�t��:u��o��xw��Y��H@�x�f"�7{'~��N`
Y����X���H��-��ֿ�6�H��j�d��JQu��1�,��������C,&֞�h^sB�k�]�|��Q�=F_�L/o����v3 �7�Hh~U�XƇ�	�ƻ@h���b�3k�+�
p�/2�䔦#�ٱy8q�Ŵ�i	��0���0--��-��C1�շ��֨�%�D��td~���:�ǌ�&І��w�כ����C��Ͳ�?kB|)�~��%��#{����y��</>H.��/]�Bͨ,e�m_EU��V%e��ɎA��e�{޶*I�~M��2���U�혖�Ī8��_�_(������cW+�������ٶ&
��A �[1����Eqg�T�1�3EB��b�mX���Gʻr��!��/v�Y}S���=	K�dR����MC3F�x�>l��K��x��dn��i�n�!�M6��T��A�UЊj2d��w,��d;j�%�TD盢�]3����+��C��Zg��NL��+L���*����(,a#�4���xX �%�~��m5A4����r���7�jS_̓��c�c����؜x.����N���������˒s]W`AIn\<�I�֊
W�-|uEC�X��b3����Yѫ�9�?�����2r��~����FT�U�N��!Y����S]�
���!$nj5�� �����v��f��1�����(� a�5�Ղ���U�|���̱
h�7ϱ�s�T�a�  M�����|�4�`��2��]�S9�5�5�~��d�/�zY���[�Xǵ(FB��+���AU�����6�*9u��8��S{�r[�J�U���NH�B^٨� �S�D�]q����WZ�s���Yf�����e��bX���%r�s�c�P�3��.�Vy�wL"�v����Қ~��`����9��q3�}_����7��4��x�2��P 
-�緇�K2�>;��?�9��<p�矌A?�̩�W����H��������;����C�dMgBv�.:�(Ү�-�x��>Lj]�O��ί�f���rBj�j�)G��{���Kx����� "��@��9�y��{e�Y9g��p�����
h�Y���g����  V��2�7Z��~H]:�e�E6<� 줯PB�쥙�AM�A���_��� D��I��uʺ�#�EqVx5�N���\)Ȫ+�f,�I��*PKR~�g	�$d�y�C��E������W��IW�Ω�?�����'���?-$�����R�oښ�G 0���M���5��׺3d=�Z6I𦔦�7���<b��q�����������'�/�0��ߕ���$�K=�	��������"���b����Q���38%����v�dD���ۼ���͏����ܛ��M�O�1��`����[�	 Y)1Cr���J8���p�=�8q�S��ۊ�C�⥇��D�0ty�wi���ٌPhd�p���m	�9� 2��H�%H�4�N����9��;�Y"[�Y�Pa�F�$�;ѻ]�]+��ב�X'WuHvWp��,z_�U�D((#Jn��D�q�C��rnr�x�`�Q�<������&�";4�`AN��h��43_�>�H��z��5X�/+{)|�C��r0,��fݥ13a�)�?�_'��[.�t����)~1:�2�E-Q��"˄ԋ�pj�
�~H�-u;���������C�/_���x��������c�d��K<��u]�S�d܃��\aI��E�̯�y����A���U��z_�<3�/@���qY�A�9��P��]c��t����k�T3匼�Ekq�[ǩ�ځ���)�O���,a��.�^����a]���cA�����^��ot����(��X1�OŰ��(�o��Ϭ��D�p�$�R&W�����ji�AZVJ���$B&�Ju-���K��jƠ��_r3�9%��Wܚ�1އ��/�����{�/�%�3�a��Y�^]��~�^��Z+��і��P���"���,���e,��Om%訷@�n���r@���S{W:S���zM��zfr��Ps�yGi.S��	q�h�$�{[�X�N��2���=r�$K����-�V���/s�|��͆�8��Q�`S�����N�AseȞ0y�����%��E��lv	7�J���~�2C5W&"u�S�g�[�&�p�0;��; F�<*�7�Y����H��- s7�|�;�Ǆ���]RCMH�jĨHSļ*ˍ���S�G ��x�]~�*���oj˫4��^���z�CI1�*���i�uӞi�a{I׮d�Cbj���O����H���[y�����dE�e���F��|,$�gPꑡ���/���KU��Jq�Uʆ��������>��NQ5��0�gUL����u�mHq�7�a�+��4����I��G�#:
2}@^Q�4a�ߖL�`J����&��%FWAk��4	>^��U�?-��v�4^�w�r��[�xq��4��!�S6�� �*������o��M}��-�-��{۶�]�lg͖�yٖ�A�	���շݺ��֖��+�e:K����߳ ��#��Yq������|!�F�����&�[�J�gAxC;@uI�Zm'%ֻ�0<V+���\K��ĽU��~���Om8�ܐ��b �ڙfs��g*�n`?�U�(���Z�rG����-yӭ �hk��Gc)댼AF�5؆k��X�M�!�<-��� ;Q�7	��<e�G+�	�N��M�F������ � ��#�&����]�#��t�ҩ���No׷�j�0A����1�vi�%'����φ���[>/,�b��t����X�m�ϋS��[P�����Y&�j| yOj�h��mk�OY�3k�1	�)�0�m�p�O��'5�95��k�(�B�����pm���:������!X�N�Ӽ��&�e��$��ҵ;8�&@�:-6�ͭ�v�쀖�bx���\�"��ț���5-�?`p��`����S�.R�Aꑵ:`�(������JrV!�D��������ڣ�pU��޲Z�jGԟ�B��V���I���桿�|y�!f�E�u�?�ѿ�\���H�gd���.��2EJY�!S=c�m�|!\!.IU���z�A�7K�X�F�vaY&�v.]��� ���im�Y���Ѭ�T���SX¬A2���VF�H��H��n�$&HpK�t�ˋ�B�Њ�-@̸��vpV\�{@tD�|�I��J_I��&o��e��U��l�k����� �m�ʜ���f�Y�v��@�xJi	���@�eY��l44�c�c_�����<���u��-�G'd�
��]ۛxF�`SB�?2��hcԺ� �>E�����ǐ3ؾ��h4��X���|L�L H(���@�`8�y�{�tEX.�L��"�YT�D�u�#f}(p����;J�y��[e�eN�u�]XW�e��Ey�K��K���
Jm+��\��n1�����G�
$�tѼ7AGk7[W��]��%���G"7���y#`ȷ��h/�r9=�<���k�@"r���e���,�=y?
!ا^���gV	0z�t6��&&I�Ը�68b֭��n�	�V�#��e��.�B�jE�9�[8�.,�ȹ�¸��r��}
~��[w���[g�΂`�&	,�!�(�zmF��7�Wu6,�Hҵ����Hu�9T�{�n$Ty�:���\�^��e�!
��>Oʴ���j�%-�$uj��>KI�D{���x�kwQ��]��j����!��u��<����͘o�����s���0�B�F|�:�:x8:�'�q�i�oT�A��,���V�ern�`����!�j�rJͦ�2�c �q^�[����/�2� E>�vn�����{�Oh�2��_l�	�{1�����9��X����`"�����^Y,qx1$���g�&�w꼼V�{rj`�m[O[����S��D��p�S_�)���o�4�Nsp|ӡ��}�P��)�#Pϊ��V�qո�qK��yi��r�WI����)�LqX���ܾmA�[�BȈzGUpeH�g����,$rM�8�R��5�~�O�����).�@�A�[o�z�f�ў5�v|8�`��b�#����nfbL�����#�h'
�*ȵ��>��\U(���Rׂsg���a�t�ְu��x(��N_�1��qQ[P$W�7�;37�����5N^�H;1Go��Z2;f"�퀈
��8�� �-�dquLU���`Vvc��&*j��ɷ�Q��X�;VL����5�r��uXRma�/'��p��	z�B��[v�
�3��P��
�S��z�)��Y��^"�����;g��lSg��}�`"�rg���!�����jug�Xd���>/�c���l��k��a�4ڒ�w��	d4䐅��݁�f/�}��y;nUAx�ԏ��2K���rnf�K�FaI�t�Z�8r	;�+��{���4V��Imz��C�I��/��%<Mϗ�hZ!��t_�b����(aݦ�_��.�����K%�O� ��U������GG3���5Zb�|_G�@qՒ0j������ib�U-)
(�|��j��dI;"{~��_��C$�(��J5+5���MN���nl.�-Sœ{����v}�����#��i�)�n�[�x΁��> u�������Ics���tT�a��6�F���oyY��`Ɠ�I���W5c ��p|7���'s�Y�Q��<mA�Z��OGx�5(Z�FߢkG�~�*�ݶ
�.�氪z��l�Kg��.� �͝��cD�V@���e&�9r�kP�l�˵ݠ�+���� N�ez�%�ī�����G+�XV�#'�D��٦�i����u���a�Y�-�	�Η����Er�L��|q�=�#�)��L��2�,������I����ޥ���|�\�_�#����E\�p}D$�ᑋ����IM��/aP!٥��XsZ����П����V_r�.��Y^\���s�a���bm�IT"4H�8��s�$��ـ�y\�Rk�hJ���[����j�C�_��������:&ә1�͌ʗUx�#�h:E�Pu;?x���l�a�:�_H�-�`Zy�jC3���WRO:���I��M7�'j��v�N?�5˸v��R����47�8��&Ҹ��^ H���m�կm���w����t������b!�g�
��&?\2ˡ�f�	L&m��'tԄY��FBc=�k�~y���v� �Ud���ek|�0��.x�p��hA*;�8ȥ�WZv]/8(?���=,�ܐ �NHi.ڡ o�{�{�!(�ah��h��T/�}��$LÊ��'�0N`?� �w�U"0��E�@B� -;nPo��iȦ�R�a�0m�I�P.�I�Ѿ"��6⤋�p��/��Ԉg-�>p��*��WH@��e;yk�J�B����m�D�*��p},�iZ$d�7��e���Sա^K�8�rӣ��H��B��	B��z�E�^���͈�Ju����ٕ��OE����|E!�JF�i4u�"�(������S��n�n;31���P�3uM f���9w�������Lh�,%���R�m�O"KI샫g�YH�L���6�bH�������$�0��W}t���}BR,D/�����l�t6���������0���>E{�ɻ䲈V[�Z}r��\�u���nY0}�5� �/�{6�[3>��`[���[��p��
�*`75�)�_�ꆛ�Wq����9!�f��-P����"OA�Pi��`�3�+�{�s�-�r?$�M/�K�[8@�e�i'��U�%�T��^�G;�� �����i�A������Ƴ���1���5p�Xw�}IͭQ�O�*5�>Vl?J��\�4p��=�z�U����Xpi	+|&��S~E�J�;�4��q�|1g�`�� ���	���	)�S^x��P\	�;�aÿ���RG�S�e��,��ŏ,w����C�6?����e�I,KO��2�l(�)K��d�x6ĥef;�rM��0h�,�ULՃ�*��z]��e���Y�� �r���e�8�۝7?TW�w�a#�K��ih;�v��	�R��~܁�2�n���1���E�:6��x�w>I�CG��@`��cە��&��Q"c
��V�y����Vw�pB�)�9��g�7�d�w��cY��Qu7�4N1 �i>�{�J,�+j5n���G}�9^p��VY����m-c�Mk:7����]r�����aB�E��ԛ�ġ|/V��:�4ۇ;��Fq�\��e�.$�6"�'^�?�.DZ����!��IwQ��K����7�g�
����7�((tn��ǲK�S����������P���k:�`��>�>ȟ���8n��n�랐o���_$�z��%��kKoy���&��9�Vޒ�x���9\i�>��$r�OH�Eb��,<�.(d�F,�rb
jKe14f�9���%��R�Z�8@���%<�~�̔�;ga�7�V�:�D�(�cI����~�F.���4w�I�R��U�~�w�!�R��4
��n��Ř�aғ潠�ĩ�)��6�\6I��oq4��҃�O������J��(��T�����zZ����wn�i��@u�cYJ�VT�(��u���Dq�3ڟDd����osT�?�Ĉ%QWv�Ɏ��$��o�Z� ������(k� �>���Z�^���!�c��Tw����8W����,H6³_�e���}�V����Od��
GUk��7���2�ZP�h��>F�S6�^Cv �8"���y@0��{��� ��&�{|61�<��ƪ��t3�g��ۛV5�bQV���k~�aW�r�n�o�0�Z(0�}ּ��E��]#��U�,���O��z����[X�.����j9搁���e#�F<�@����t���;r�2�H��&= K:�NO	���~�Bx��=�������߳�zr�@�8$�n*�eR��+r���B�&��OX����28��<�C*�A0+f�-{�u����	�=���|^{b�l�e���Gf� 
�jK�*z��]z�hU��H�j��g���1�ً��>���3�����|���&��eu���0_{�b
�}2���n�kI�Ѭ�/�s{A�!�����[�Q�p�4�~%���el7~(DP�?�ع��y)*����φ<���+=2��л�K�A�ڻ�K��F�N�w�%fv+�RT��p=F>�K�_����)��������4謺">)U�v��k�3��R��
�CtE���;�D��r�MO~2�LF��1{ot���u��q4��c�ðG��*��N�=6{�/�ɗLl/\��)a�aW��@�k(i�KϵN2ܰ��=��W�Dd&�iDE9�Z=�Q^p��n�JL�=^e�M��?�F�<�P
�'c�3�+w����-^t��k)O�H?���?��i�X�G��{<�*�;��� �eP�@�iN���+D=k�?�)�|�v��/fPspCk�g!yi>�1O�Ĕ���4��M:�c�RS��P�/��q)��!���fC�2���DG��7bK���@��6B���y�?V��57��C}e�q!�8��I8��x-�SS����z^����&�Xl6��_�`��Q��Z[.����vub�)c��i��cNg�@�_�	�%�=����G��U&�ug.��k��%�[vO(ښt j��Ar� }nN���>A��ke�}�aB/��XEg/#պ-������$���,u_��һ��򆧩̙��DA��O��Og��7�S-�5��'�F�1/_{�f��7���hq�cǛHq2���:~'�#��T-ϋQ	�'���#� nʂ(��x,9�k]p����.���+��ӓ�����K�b����0�� 6�bYC��BFޢ%Oe�)F>����Qq�4���P~爥~�����Ģ��j@*��G-���/�����:�بi3��9�Of�����M����ì��Rp�p���MC ���TC��#�>�L��(�B_��$FW�ŚkQ�8�ww }{��{�}�kT*�^�{�l�.�>�4AR�����B��#s��E
5)h16UKP濘��5�U���v_��t4,�����~�Nq��H2?Hʻ�٠kM����@m�,v
���vc��`.�˩W�؂�5�L=QS����9f��)��02��횴�����C˓jF���(��I,��$�SZ��N�Kђ�ڞb+��Zk�[0����E��g�&�A8���=�U��ҧ��,4ʕ'\|��@����eNG��G�כ�Nb��:#4�Ò�o�������[�l&��L�O��<'�0)�J���)����Rl�����E���
7e,߁kL��ID	j���1_8Y8��ӦY��Vs��{�A�
q����t͖i�@`�ʦū���R~_�=�X����i���#�-����&��Y���҅&�wc�!`]���&�P��Cͦ�p��D���B���wI���j��R�PJ�1���9<#������$H����D��㋶�C�L����ʽ�� �;	�=m+r��Xv	͈��p��9YMG�
��f�Qp>2�¯��"-δ�)8qhH�����!Q:�M۠A�o���T�Ǖ"�������Ji�~�*rbk�z��P��w�DQ'�C�yTJ��7��p�ȗ���n��V+Z6bؒ����w�ǩ�58���|
�΂�0:6\�ͧ6_�Ե3p߬�"���}S���!���Z�.��K���QGEI_(��69ذ���i�g�o�I-1��b�X��kDީM8;T��&�%��e؛c���Gth�~�%� �Zk����( ���V�<�q���CU���f�rM�ep�Vd~��Ņ�m��z���~����&gGh�Jx9?"�`����Pu�K��A?Yi;�C�^Q1�������TvR��3�.x���Q�OI����v����$5�D��Ȅ>p� F`��O��C~����-	��L�'0�ua>��QS׺�\/���A�;�pi��%�1�&Ī7��� ��x�9��=���Tu:Snd�RT��5�Mi"��y��~�ؕF�v[�cC�:Ӫ��I�A8� ��Xh?'YJ�@�B�*�����g��	Gh�X��%$�q��x~6`���ڶ�a��.+n/��)�0����mYiF�EB�1S=|��D�D7ʱ���pc<k���FL�k�n�p�BG>�G�\x���#V]yL��&ݩR��:���ʣ���G5K9N���	>��d����.�ӄ^�Z#k-�q�u���=H����$��>]��Nvq�R������\�}�2��/�QD9l*���@n��r�~�v>U��! ���+�e��d�=��0%��!�����e�	�EN|w���@�u@��B�"�ɷWD�7����N]���ì���)/�lD`%<��Iݞ��v丵2���<�l6A.�W��|�ȟ�r*���n�:�}d�E�O�n�0l��b�Tה���;���V��y��Ł�5�f���d�n�rgѐcs�NZ������:a�>�IY�����}�j�ТA�Z8�Ϗ�<�Z�w���Qb���R��*ތ��;�~{u�8�~(��Wy%�
;��A�fzF�r��ο���2�X�)��;���*3���(��-���
��#]�V�,8)�7���:QNT�!�uyd�{�Z���]�$�ó���S�)���<�,,��xrhb�\�`�������`eS=E;m .��Zd����&ߐ�*��췰�-�l�;dZ�u� I�xA|*ފLJ�!��~Ԥe[���4��-oze�05Ε�e�+o��1(O��JZͺ_��(5����u����q�2C7������̃�)ߒ����[Shφ,x�R�TCs,(2���u�fϯ�h�l���}|Oǃ�p��9ZO����K�;cĄs��� ���$ϥ�'�r]�i�s7�s��(�\���e�#D,d�f���Xt��k�Ha�o[O�z��*�l��&/�R=|��n�K(g��N�O�b(��3N�Ƿ>i����$��~�n`��?��G�\̝�L�	x����.ٹ�n&AI]�5=�f��߀|���]�LH�V�Ȗi�����K}��rc>�Ll��sZ��]pj՚��|�=�Pө�4��B�9�g?9��'���|�}��5ݏnύ�5|����E
�#����=t��l�]�ȦK@�<��;%`�@����x.�����"1��:u]m��N����w�_���Lc�v^�
b��_�Ԯ�1�9����8��q�RZ!�ǿ�k<rG�ضk�­D)pp�Y΂3n����;��w ]$���U�pg�ݓiQ@�H�����۲�P<���Ш�YK�De|0�\�B���q9w1�*n��Ou?	�֙�IM�ｋ�7bi�3y�!b�^�k|B��^c	�d
D=�]�H!��-@���j���-���~�	�k�(�-r�������� 
���1 ��ɺ�$T*$Xb]��*���}�_����Lь�z�P�$�.:���tCO���W�SP�2U����H&'q��zr3�V��� L&yh�i.��H8�onA��ͽ�՝�픍�w)��r}Ɛ�<��/��{���I$��x�* �L�3{N+v�uS[�|NYUہf�1��K����l�������G�H}P`:�/�Mݱ]�Db�?l��t
#��և�6�������MTz��ci��pqǶ��&e7�W�@z���P�Ǣi]�� ��KY|�:Y�����h*?�8�3u.�@Ϧ7�� ��<��JW�Llwm�+��3:��̀8��FM�Q�U��B�yu �.�p�W��-J$`<�O��[Ã�
���/����L��e�Ow�OF�X9�p��>^�=�ŤSӒ1��{q�KCm�Rw�� J��) &�D"�dѫ^�
�)!,r��ͥ�+P��{��Aˤ���T.��d��=W�(������QG4)|=(@�Ԑ��Ω���H���}R쭏�;�)��Ȳ�GR�)~@����"q�ZGs$`{Y�?�T�e�jV�N�X��H�-����<����, �U"|_��P�h�B��Os��������;��ؤ�v.s�>�
W�̄�;�^��eY��U� bʕ��D�(�V�ɣ����t65],��%%8~~�B�8V��z�r-6{�?���D�Ɍݽų���\?���������
��:��B8r/�A�\U�d�+�������b�'$�U��]cz�II��_� @h��)���W��	-Br�Lz�)J��mjt�IB~�ue1���r2�{��P�%~���1ɉk���p �t�hQ�9X�>Y�],�9[��&?ں����C�_�,�I2��X��T�E&�u�^�Zѫt$�R];"�ʀ��H������U��cϩ(�9��<�?+�
f�=M.���a�D]���;CX9і	^Vt=<�H3%���O������3{
u�`��1�FB��l(]�Y*"��� ��T:4Z.q�T��5�C��.�}���������b��Q���RIoWG~c�99�{p�u6�/�K����ߓ!���y}���Cb�I?b`Z_��K�-��Ɉ4��Ҝ
*�����6���ܶ��%�!�&b���y�8�|Ƙ3d�9��a���l��4TμW�%n�/���Hl�o��c38+v�n�,_��b��x-���k��Z`�"F~�6� r�v�4�+*�&������C���$��k����T�>�x��맇�&�ʓi���׊C��C!�T#��4T��H��p��j�+��zQ1�J�2�O�O$]�;�,T���Q}��H��,� �8w�-����{5=}P�R7�k����o���Gu�X�=�^�r�Q�r:���q[�� 8g�^��|� �.��*�g~a��]��9Wr�&/W:�\�A�Ed��F���엀��E;#�|�2�WRs�������_+�˅��ڶ�&���X�ep�����cx���x
~M��x�����������@��|8��xld�Jw�}�-��Yv`k�Z ۱x2�o/u�J��q��}�?8s���T�T�"��/�]h]#��$�G����GL(��<�9��o��h;c��������ԪͼP��GZ��6[D2�E�6�~ss߄��r��rJt���遼
� 2�4���@v�k�o�<IM�X��%7������S^�4%��&92�k����$�AM۞�WW�� �5�=�?��_^��K��\�TkG銑�͢��̀�}:P���b��)Fl#/yê��ݘv�vI���5�C��IS����ӈC?)4�� �_�.�˙��L���_��o�#�j���[ZES�W���;Dry�
�������j�ѥ,��c�8%qݑ�Z�8,��a{{z�����Ä�T�r��2�������������,9�,dk�����rɳ�&�!@��O�����1X�e��ڢ::�x�l��`�L�ȱAVe!w[�=Ӌ�i���Xo9`6dY!\�?�"��&>ᒜ�5�6B@=����9�ÿm����4���BB�+��WkP(�Y��E)�CO\J�o��XZ�״�4�^���siM�h"�����]Z֕��e���xV�8x�=)=�@����s��������{N*��-���&����	2�����'�R�����ǂ��wA���m�)7��3ʸ����0ܸ7#}h�Z�Ӟw��:�̦������.~���&]Kg����C|e����#A�Sځ�4"O
�tp^���H�2��9��!T��v������?z����:y�3��洺�i������0��r���
JR$K����ɪ��(LƷ���#OB���oJ�m��s�|:W7��:��Ѐ�Jko'*D�IC��ԫ8�S�)�(!&H<�ҷ�̂�~O��{��3�Ei6����ۗ��Sg�ӱD������'atBͦ>��u(ly�Tԯ�55j}�܀NY����팼�n�����1���, ��c��m��/J"�2�D��,;���>x��O�qi��'��;�!��P�r��FH��I�V���sK��qo�XI�ƣjoEe=�{:��.����ƒ��U^�bt�V���Pγ�O�3���}T8x:���-��g)^���$	���3���ꝗ��� �,�W���U4��(�s�B�z�'���"��pY(d�j�u/RQM�T��T���,&�	fƩjan���C�A��M�6���������`�^�c��=�5#Ov�F6a��޺�G}7��R
� �u���{NyX�u��%x� a����vM_ܗ�mY���СB�M�� sF�Z/���0���B��CH[:o���nYHmf%�<� �9��6�B	hT.��0�?�O0^�¥�R���/Dk;���k��s~E��G�+�K�TŞ��T���y����v�M��I�'!JIP��ސ����m4��&���;�|��� T�~�-s���6D�$��w��=Q"l��/Jࣟ��|hl��.,���L�j�Iw���P�'}�0��N�G�|-�z��6D�eA` 
���ׯZ�R���u�a�F�+*�9eKvOG� �5z�^�zxha�}��J�w-�"��F���`F�״"�$)S�_�?^^�M3��ϊ�ն���hѷ��� dVoL�#���dW��5Ϊ�������}��7sP1�=�B:��.p�i��[����<�W���fK���� h�f��Uzdc�>K8�3~����%�=;SO\�ԁ����>�[��4����L�#�o�*)��$��,��v���zd�=���#�������܍��"v�;��K��V~L�����?pG�6}Dy?P55Ex��/���Q߹ H:�
.���Y�>>�!3�G������T�|32؞�U��$�%���P�Y���;��܁*|C����������}T��P������D��e�P{l
|��x @c̩XG�ֵ���S{X�Y���x��%�u����@5I��|�>����bE䜅9��0�^�SY2�"��X�:���1hvŸ @ �b'��1)z>�K��Us�$���JL�H@"}'	K��U�x�$7ԾAd��)0��L8%�'s�^<�Km�(̘ă�!?M[�X/$z6Y�=Hk���<"0�>2��6sAWe9��K��Y���w�? ��2�Z�p��ο64{���dA3V�'ݘ���A�n���?�&�xMc�mT�wY�|[�&6��EEW�~��O� ��O�j�N�!1&V��6��"@�$�S��-e8&ԉ��E�3�{T1E������Y�$V-Z��h�e�����r���D�$�y���3�5�9�	^Y�!��x��7�4�������x����]��C��1S�����k���g�� �*q2��n����t�0fճ���ƹN���G]D�+�:����O怕�S[Pr�8x*-E֋��-p����ќsS/�}�;��n\u{@�B�ѴoqIi��C�e4d���^�j�f��-�bsvu=ȥC�Ug<��1�ҫ/��|��#]x֛yiz��uyr�2Q�4(�]��]2Y�Ӣ��r��O�N:��1yc�ʎ�X�i�%̲��Cׁ�Ra-�p%^�TX[8��=Ɉ�V�z)��4u�~����@�Ƈ�|{x>>�ј��]}Q��D���Qў̟�/�>�yh���~ �{�I3�Ap�3��f��>�]�S�Mb�p��m���y~��{s��B��ߋTɔ��	>!�6�Ep�/�n`�����#w#��@�H�|?����{@DVV�o/��|�����Lwd��(q�K����r`��U5�3H 8���s=�'T�=þ�tU�k�z2�"9(���S3�a,ed��6?Js�;+�����Ab#�J����9�P�x�U�I��-�ҡS�"tS^��ф�܇�p�V�ѐ��~��)��+��)<}��4M���Ňo'$$��V�F��_T�ٖY_��#�D��6 �7�2c���'�Xj�l���^��)����!vL�ם��:����A.>��b^�jL������� m�`���2�0�3���� ��U67{���MCtcU�ӈa f���Ąо<p�0%Db���a��Dv)��,���8���N#�
Ur�] �r�ǚF�ti����;"�Z��ȵ�8�UF�5E������~�*(0S})n��*���,�T�zD��fq�5��=���+W�����C�_|��>.��w�����ME�ĎL�B%`��xx1�% S�;�6��r�+��v|��(������w]�k�񶂨��\ٺp# "% #��k�+ezտ|ͬ��:�����4���9CH�Lc�vc���7�GbU��s�
<=��n��u�,٠!��^��gIA���:��b�{���<?Ɩ���B�J���#|�.ʝ�a8�^Z�C�,K={�7�t�� -�D�趺Aww�	��P��.��배X����U��OÝ��:�*�ڼs_A������e&�qq���<�[4���:�VWǋr�Y�4����h���tp"2��=[6�#L��4Q��cs��L��[��,�Ӊ4p�x���U@��{�wQ��q�.�kL�4�"����`�Q㥻�g>e��%|��d>��[���&�a�mړ��~@m�T;>`h��+=��S�1t�����G�O��cp?���Uɺ��������PPb�- @^d!���}�����[�~5���cf�I�e���7�î��$��X�BL�ᓏ+�h?��C�M��΢��B[Xژ����\)mtR���?w{�tI;@�eLk}O�N�Z��)����9̮|�&@�5��.1��ט�@. #��^�#�P��R��=����뺔Ɩ�mA��1qV�9a���h'=������Y��«#�T��dۘ��n?UAě��;�2��zkT ��_=7�%�\���#�z�����c)J̡�����&�1�G�:ދ䇲U�l������k*�Pk��8�8�]�����+W�=�[���x��x���5~w��{�~!%�e���3�UM��v��Lk
����A�q��E"� 3ͳ��p�	�Qm`=F���]VP���gbf�iE�V�g�D�zb[�]Y>�p3����\[0��� �&"��~��@PR��e�a|�h��0��hk��IӖ��OCa���P*�=���-痊[J���	P0
�L��䵝��<�b+(L��=l���$>~��i,F����k��j�jܠ\v��N7q���ױ;����6�6��A�f"3�v�ǋN�w�=$_���	�<%�����/Q��ʔU����Xxeӱo�������B���ʇǞ��ۊە�b?�d���X�1�Қ�~0�)>�ƾ։�#���5R�� 
a�Ժe���I}J��Z���Oq�L-��pn�w,ÍՃا0��_������CIׇ��F7U��SX�������<�!�cl��1[3����gqhQ��D���[�\�x���s࿿9C�,��o����X�p$0��V��Ʌ�k떘��cV�j����J#g��<�s�5s�E�G�mX9W���c�7���3��5N�(��rH�O��,�D��,shX��^^[���\%s=�O��<i��6�uqg��+�� 껯w���ab��1���7N�a���G��Զ��=�m?im�{ϸ�����<�s����Z*f0eėLן�v���%`��ۤ ꐅ�
k �:��td?�;���JM�P�������5�����!d�d�BZ�`f�B��8��u.E�)a�&p�D3x�-��`��l\�5
q�h���w�����_�gY$FGg��r�s�т�������������\1���܉70RU��iA�8�i��#�p��C�pu"���J�	�� ��S&�~,�z���~���e�:ua	:b����f�	`qq�A�,+�"��>_�8�u��Q��ձ��)�y�n����q������P"�`aF�U%�t�߮��:Tm�1���l���g�ş�4m]�3�V�tZ�ŗ%4--�h
�&H�,2��
tx�*r�2�UL6� �&AF��,"*�A�f��Bbp�&bd���w���6T͜+�&�ELv�5�I�:W�[���I����fT����FS�W�N�l�1���p�C2w�b'ܦ�U={��!z�.]��}��up��P�cw�_��̜��IO����i(U�����F�ţF]�����l���Oeۿ���3�fzz qG�����!�q����C���@�_�����E�����^��u��6dd���bT3Ώ���}*�i	��涩@Gd���S��A�7G������@�9��U�C�R]�0�V����I�)�L0S���!jU2tӥ�~��B6
+��!�����	H3r�~��:�j�Ѳ/{0�\Ց��3���_���k�-�`��E,�T�3�n򋫪s[`S07�
ŀ� ���P��}�^?BG�F͌�So�A�/�����&������P{������a��)#5�f�*ͼLA���J�R��-��)�3&WD�L�y�&������¼8��`3dZ�������M���+I�.���J4o���/F��Zz����8B;�Q�J9 ���8�&�ό`�L��K8m݂J�J���@Cij��|�g�R!�qYy���}���V��
b�n�)>%ȥ��MM���"	ڹ��#�}���$�S`���,4ᚣ��	/�E���;�}>B��u��0�F���*I)4�u�AvM�kϧ��ef��ִK6k��|�@.C����U��H�	��⛊5 2��J�9M��{���_4��#l�{{�	�:7
Wt�i�ָ���,:㯯���L�*��:'�o�w�g����\��$�	�(WCO�尣�jW��_�)9�0����Vy?1c��Z�V3r�K����#ܣ�o�q��qu���2l�me���q����lK\�j�,��2��co�͂�3���-���[5�S'��2��Fu���VX��n͇S�s���Z�;b"~��CP��`�,Ӏ�/?��c����Y+�ْ0�\�ak���pk�	����_��֊�E�)�=<g���#t�#�G�����ӻ��(I��n�f��B"P�y����bc�EyC� f�h�����mixH?��̳y\q|5�*S��z@���Sm&��[֝`�M�Vi_u���˷��-b��T�N9��T�a�D�����T,�΋�y�G���x�V`�e@:x��T��օ�j��N,V��`6O!���֝4Q��R06�&\ �����[]a�j�x��]��}>�;)�d��`���EMp�P2��-�l��,��X���]f;�o���ȩs��6K�D�.D�
{��c�����t�U�%��1^Cl�bփ�d�����F�O��������X�"�7��||���P�&䶁��\x0�0�l;,�)�w�8�a3Y%�o��X��C��D{>q���2����qr�#��:5��?a�4��{�qB&K��g�2Lo��:������!sj��TM��}�yh��9����߫�1j��7|��b�1��%��YP,� $�B(s����]��y���[m�eF�AWM]�;[�����i^����϶��9>��!�W����G�NT�y��D��5殳]��� �Q�i`4e��hg�ݮXE��&ve�@�ޠ]�j�A;sD,�`�v��33�{qi�7���[�i�8Ŀ�[����x�<Wbjb����7*�Rm��&��y$�`4�T�#��@
��ݲ4��Һ��
�\�ζ�3K�F�w�+�
�|^�m��+mS���0���Vxh5U���w�Xp���p��� "�����0��w8�K�?+�ǷZHݗa�&��ꇁ��͙B ��Ѧ����e\q��I� �.��"�(L��+��Q�w�I!��Y����a	����$΁@�lK��6��J��
�GybZ<����0��XO����ɿ�_}^�4��@����9�؋���dE�}m������Oj�(�O��2y<�*��lWQ���8q�S��%�ۄ!6�6��(n<$�E!��5��=�����+��YH$~H5P\�bR;�$O�ABI���5
�L�(��kG��W�cUݦ�����s۞������2�*��Q������w.l��lL^X^�6̋r�D���%�Q7�ľ٫�N%8f��K��uu8PX�L��='Oh�z7`�E<��N�p#3z��O��t����M�#�����m��m�r��r��@�ҀP#��h��Ć����;�Kr��Ȧ��K�h{?�c�'���)�[8k�Z�r[R���=5��E!M���xF�ӭ������W������.�**�����y����#��;0]���NC��>�p>�96P��Im���q��*�1���}�/!���y��`�ZE"=R������}*�4���էЈ�G?W�Y��b��Dǰ0���>�*�r�
$��&�k�c��[��j��6#~�ާ���z���	O:!JE�@�|����;5w���s7�v�,�o�ȑ׈u�+�� ':Q8�6���l{�M�E3���/2@�D�P��|D���<�-��!�Ce1�C�eOo������]�I�Pu�ȶ�5�h�;�I���1e�v������Lbk�̯�H��Fth�(;h�P�E�1�}[D-j��V�@#-7&���V�)��Vf=���3���$��+ǟ�0����'Ρ��i��sr�(�ti�����[�&>W+�a���4
��h�PEsõ���ՠ%�0�c��4���de����bf���H��֫�ܳ���"��H.r�8_�N�3�iR�����0��0`��[�+x�?�L�}����C��˘P�/��IsKڟ֕�D��� �����:��&Q��r\������!�[ B�X´WM89�<�h�	�4��Y+z\6������?D2����zq<����!v����e��bM�T^�2Ј�~�Z��&w�]�`P����"��}ji���x���+R�ף:�/�9�nё��n���������\�u ?��r�?3�>RL��E�bOs�����^V�+�u'8:�_� �(~ڄaqbc4|�6̵���-��g(�l+JJȟ���D{�L0v��<�O��~C�pP��{wҫyF��XJ��������o>��=�W�>����Gy�����X:&+/Ar�6ia�ˎ]o�H�x���	E���������ilC��6�!�¼�u(�'�w�CB�Lq�Q��j���eB0Y��ȢA��ȼ/1(��c>=�1�;j�DM�+�v��C��k`�X����B�`���רt�k���9Ŀ�J<?In@f.!`dھ
�u��A3׭�V1�d3�?�H��Yf75�4�m �G���r!��k���*��O^,�QNU^�|�;�/�-��<V���eL����_�sZ�G�[�����4SA"�{���3&�ʇ���V����Ib�t������4S���=I'�!��_Z��kU�KT�a��r&��*�g���g��SUģV�^'��h_��W|�Be��70�~�K��	a�/�x�;���� 2�/ϳ��U���.��	�n�������h�(�9� V���w��OZ�;��밝 ��{�/9I�m&J�Fl���G���U�81XN�^��5[�A��W9��s_����ק c�h�m�:�R(�,�	�S	�G��!����)VJ��xi�Iz�V:���T��+;��A7�%kjͱ.EK��K��EE��]�_}�$x�Å$���J�_4����.��1�^�CT��ݹT�ݖB������1| �8i�	���0ʉ51���T"R��	�O�(g$��Q���CUn�群/A5����\���Y��qmj�KY� Ǭ�͚IU��6ǝD���Ih���ZY�%4����i� �����Z�&�(w�X
���;JNX$����m��H�V�I緯��͆p��nU'��b �e�\�V'�`�X�8%U���T�g��H�o&��D!h$�(w�a>�]{��{]X�C�8���rQL�]��6p��<-��QA��hE����Sմ����ܵz������UkO8�u���Q8�!/ǀ���ʋ�k�ߥ���F�6���[m�Es�s�7�.1��ʥ�Pen�T��$����h�b�8J�N�lS�׉���%��֟���`&�Gg�R������n�:��#`�H���i��k�∾	�Ō �Az�4O�).'��h��6�Y�I"K{�~�]>��|��<sq
�=�ʖ�p?�������K����硫n�m׶(��V�����h\�ied��l7_��vڣ;�/�wa����@i�9�ԏ��*1}θ0g���;nȡ~D(XTTJ3�����-��@:Q�h��T��h���M�W��6%N=uN��ȡs-e!f����rR����´Hm�TG�uˇ��ɹS�����ey^�JY�w�d5�:�d��K���зt��dR���[��C3!�;3\��]/������qw����&�
����C�Y�#d75��T�e|%Z�5A���{�R��Iqa�?�!��Q��h[Q������:�0�Cz��|��_1<%2Ş�>. �0�<f������li�y`|ŋ�NXElIZ��v�5/v\R��y��EK�a��T�������|3Œu�UE�;�>�2:]�駃�f�ҽ2b� ]�=ͪ���Rsg�Ƀ���JyVwUE@���)���'�|�� S�8�H�t����a���� �SՓ�^fy�<����"�[�.7��u�(ĔՓ�N'�3�ښ\E�@�\�$J�]�U6 �^`u�qF��_�CN[&7�����2�i�[����cN�[Ŋ�6}�g����2P��Ri��df2�ڭ�_�c@ݧ�����9�H�yC���N4��O����6����&��:S��Z;��ĭB]
�����D��B�#C�.[�ON6ZU��7uN�;�}n���7��	6qe��[|��G�Z��e@��)�=Q{O�������&�50 �K�e�B�ڔ4�8��H3$#y��`�M�&��O@�wF���0蒚�m��}4�h>�%X���_<LF��r`i)b{)�Ғ�Ko(���/�L��7��aaf��DkɃP�܂MG6{gd�ִ��O3��S�t���u�3i�Bo��t��i�\���	�G�Ӷ�!�^�1��_�	�~�J�H��Q���1¶{5,�|{~^FT�mk-���/���݀�Ժ�ұ
���	X@a��%�0ۧ�g�$���R�{<S��z���a�f�92�S{�6R8$r���i�b�Z�a�\���y�� %U�{/�#��4��oG��R�����<B`�ѳ]D���X<u��<�0�S��>-[P���#���^��7�&��j��B3���zǃ�v�ҖS$֌-)�3üEǅ���3�ǩ����,E�S��]+n��BA �X4�`uGF��/��e,�@�D�c�ħ[��0�e����US���;g����A��?K�렶`��&��;b�EK��ڱ��t��t�tU�N3�W�I�֥��o/z]�W�HW�/��]�R㷷���XnT; �E��D�>m�f#��6αA��I�x��E�A��݉�O|/(uc��g�I��U�)A�aJ��g�dCK =�!.wdN��U���az�|�jG��E�y��v4���p�k�;>:���8�m�<�����l���G��rG͛s�0���)����m����
�w�SP0��b�9"Pn:�8��D�ٻ�JF���"i� ���P�A_��.������#E��>�rm�%$��l�Jۭ_���a��xq�6�IF�ǉ�]���ˇS���e���$E�KY_�q��]x��o͔W����S+,��`m����4�U��0�Q�U��.ZC�o�����%K{�F0\��萉=���T�i�X@� ؚ&����i�os�z�~�����v�X���������SP���sSJ���b��L/�T�"�����1��/2��R�*�%��j��d(�:Ґ�&=�%o��?`�k$�U�"�h�k~���u���4�2q�֒��L1/����B)2	}"�vl��Q��%�mH�n��P���	A��o�>�ɧ2�	�'�����O����+�>�?��04��=�ھ�z0͆�e]��Ps��OCK�Ґ�?����d�"���|&	><��3��_Z�����O�fER���LqcSO�J���Pi{�U�3җ\��~��b�nGx��`Ԛ���D��5*�	$���� 6��xG��	m����p!��{�q6�Q~6����iz/���|gO瘿����!9u���qL#0!%�5�C���u���vX�h����M��®��jt��⌚�����&a�E*II&�rGU��C��Fobp���?����wC�.�֮�P!RsIÛ�@.w�w�r��K�#��_�[������p�ab�RkiB��6Iϊ�J�@Æ]�pQ�s/Ɔ�������w���	G
�,����>��㴽/�Q�*c�h�rC���|��$P��D�$s���t!c�� }%F�X]y*s�nO�F�?��%@~s����;YC*�=˾���`��)ӿ�ݫe�@�����m4��&��Q� ��iX�����&��kE�+�����{����Ht�����%�G�ΰ��:�r��Ǘ�C��׳d�߫ÛK>�V\������ zVŋ��h꾁a��^u�MQ	���P~ۙ/!*�̅�Pr�c4����>��-d�1H̅�w��U$a�q>)�(if��%8��[K��R��5l���<��ZC��P+C}�.i��L����Bg�O� ��+ ��0����cȡ��T��Y(8Cۯ�g~��H� �A2lFڭP�,U̙�����p��{��u��Wd�T��`VǏɦ��4yay��T�R/g��(��/�T�p	͐R��rwb4��I�]s�)|f�w�ٓ7����<lG!N���	��(K5>Y�?W���:��0�ި�������_�7F���~�@nN#��) �U^�~��H�zUu��N.D'��#��Rvx'd�4*L��]�CƜ��F�4}ʹ+���X��"�D�G~�y8^(h������P�w�A�Bufh)���+K�$\J2l�[���������g8�LG(�"�j��@Y�~ۚ^㒠cB�^�oQ>�5wI���'h@�s�0�U�	�pC�p�d�~��fu��u�T�ёM�N�B��ޤF+�x������{Z*�����U���k��ӧ9�)�z��ŖetjS;m�s��4W�UЯ���Ѱ*<�T�\t�䰥a4,�H������M��Q��X�B�$�)b�zT�゘�@�\%��t{/����ǞJ�U�����F��7��'T#ʺ���\�1���Q	���yCJ����`�}8Ef*#��X�K��j�	�|Yle����`�(���t{�e�V����*]��	�֟�=	�@9j�F#f�v�{�~��/�|�����Om������Q2R��.���u�e�9'�=W,L�4�hV{����[9��0"��[?�ݙ��Ac�CY��yi!1e�������;m|=A(X')�U���p���\2���e��Zw�)[6]��'C���J0!���+��	_i3��ց��h`�H>�Ǉ{'��RN��/��'5�� ���y�a���@�u����' >�<k0�B�ֵhA�(���w�Os4筒=�/�e�gЈM��q���>������Ŏ������ ���U| �V�=Qܨ��+r�W���ì.[�K�3����8��y!d��!�^���V��`���=~�g�6�_�;����Ar��XA1�-���n-�fw��.����Z@x�������o�H8�o�*��Z��W��e˔��O�K?um��(2ߑ�=1�k�ks}���+�l'���RE���8��|�8S/��Q0|�� ���[!9�:J��c��Z1��<��KS���&�bO��વ��T�A��R�H��vte'@����9$#�I�	�ː�ސd�nl��%����统U2#yW^���o�:-Dy�Η�v�o�:h��aV���!i��}=b獀/��~���r"�(;�ïm"�m��������2sR�MD�dNr	�OzV�g��KRM���%>n������A�'�Յ8^�֖�Q�~�/B�O2�]���^��S��A9%�=��z�����2��V4��N��ćҏO_��z��r��i�w!d�T���qf\"�f&x�εs�b��O�X���<< �H�FΖ�>_ʢxLHaʝ�˳5�p`�98t4��7SD4�$�C��+�礙���" ���CM��с3x�"�T:��oG\��[!��g>�jJ��R��H�4�����bk ��ҝ�~:Թ��c΃g��zD.

� nR,r��͛� ��'����hU3��N��0Q��������:2�ǀ}�ێƆ���b@GB�����58���f\��)-c�`�*��@�E�V��|6���'����0I�W���3������}WƞǇ��p߂�|���HW\6Gxϔv� L
����M`@V���KRY�#l��Ao�7t�X�i�{G/I�ŏ��,Sf�e���<ۥ_���M�[+A%���}m����;��.L�Bb(S�l�X�M���:�Va�OĜ�B6�a�/��!�p��ox�U7�{X���6�:�D)���hn�ߥ���</�x�!�#��6��Ѿ���̻�P��s�)J �N� �/g�N�~�X)�2��EO�椾$y�C���(?�_zvw���oS\ݔ[�X�rn��y��q]�Kh��m�J� K���'�Y����͓H2���ϟ֚�:���p����]տ�I` ��������
3E�[�b�{Mn+e+2���A.�097�����i6�,��V����@�q�A��4缐ce�v���'�/�V���Nq�Tb�>s��֍��£>𻏈��I#F�	�wMTe�nH�똴91�o5��/��f�c�1_b�6��]}e��X���\c�����D�Na���r9�#kf��3���+�&�����p�����MI���Q�.�:rx�x�Q���~�L���h
��ڗ�I�y��o���U�^H엝�J�s�� M����I�\W�b)~M�_"o������ l�N�<�t�g-�jj��-���OQ�zO�֦�)�?1�(;%�_k�%�$Vx~����C�R�0���hp��^X����9�~&�^-�β;���~�P,h�����lo(��P�t��,��U��D5��QF�����Q���)59�%NU7!0f�m��;���6Q/��B���Շ��/ɵ��˥����rzz#FR>����/
L�l��3�k�Msuf�f�Q���/ՓK�B�3�)v�>����C

�+�t8~�5��g�]nr�	�*V�9P�/3��M�C�i���8I1:����5�A�Z|��DO���A�wZF�b\�P�:��h���2�m��t7̃�"����z�M���W�5wT�v�$*�����j��βH�t���^��|�*!�SL+ٶ�D"U	A]�8J�4��)���R9[�kgF��x�S��Q�&�١�`�����B�������0�v;�_��t��L͉0��P[����c��9鳆'�"�;�Ě�_�ӂ��f����8��Qİ�[v��d�wY 	t>GN��sto�v��<mO���w��r1���v\�&&�,��(�ך*�A�L�IwR���#c��?��n�#��C>��@4�@����k$���GE�ˎ"��P\Ľ�;���f�xhۆ�8�ѫ�r����$T�#�Yk8�am|ߌT����+Bן?Ab4q~7|����^��{iJ�*�5w}�Q�7��������?u��#f맮�YC$S)�A��V�mQ�ɗ���y�v!z�)�:��Ȳ?�nЃ���E¹[o�
���i�N�#[m?z�e�ٕz��Av�w(J^��y���>Sr*���k��q��E���������_(U�_\d��#��E^
�C��H.��kM�-F��cfPK!�h�M����G�}B�WX�Ja���Q�u8'�%Ԛ�z�������������%���0��F1��I8�=�w׳�1���Q͟��0:�~������F�	j�)Y�����ۿ�p`��J[�4�ߍޔ�f[0�%7�V�,��k����{�!�+�o'#����z�V�	G�i�3ğ����U���Ԃ��@���d�7tb�in���d��;9?��{��v��3�o|5h�7�ml�W��q��2�������v��%���?���UM&i�\��Vs��B��B3̮uݥg��$�����#g��Ao���T�U��s�����n�B��=d��29��T��g�s��o�ƪO���B������E�}�aq�~S |*�fn��7���P��/ ��<���O��Sd�.6=�t���T�_�=��hҴbd7T���A�M�����i9Me/���5��%��d�]*~I}�/�
4��oΥ��l	p�P�l's	��0�����N[a�)��w���U��� M���-H�'��n�m#�0 m�P�*:�	��I�5G偩R�l����V�h	2f�"���p2/���S��I����D-�}����&F|a��t�,���ӥ�3��+sʪ{*�}�z��}!�DG�.�y���g�%S��x���/��k:�X����)S�M#S5�Ѿ�T&	EMk���r�6��������n����+&
�ÂA܎2Un0��[x���m��?(���E�+A֬��z�o7�QJ0��9�prc��AZb|�3
3�6ր;\�L�b\7MKk{�e:p�i�B�f�Ȓ���"�����.��y|�I֏�7p�X��B���Z������>ͭ:a\����nw�;��̈�~�~{�G�=1@��Vt�&�:�mK>F��)_&%!�:�3�������,�\F(��M�/��[u#��|��Ң�<t��t/��!�X�=����3�g��m��=���߿��^t8��83�~�ӟ�F������L'�rl�RŬ�8Fg�e���T���fɴ��?�ȕ"z�8�X7�]o��~���AY�H>m�}I1�u����O�|��68�k�]6�ic+/�"�%�x�[�/�%�6��l�DM�^��qrε}�7x�b'֜��g�<���>��؏�'����̦�c;$��^��1	�x78����v���(T�g'����&�ػ�~kUQ�W���iM=���� ��C|�׍}�M\+��Y��$R�f���\i�C�8�@�o�'љR���"�q-y	�8G�w�lY�.�e�7r���\�c��e�~_�e?�b+a 0�!g,�������$���TO���H"^��pbS1��l����:"�.�B�]�D�l�:u�X�O�\	ZC�ػ=���I��6���	pj|���=��XǼ�i}H�U�qeB|�[�����^:ON�n�<���Ml���l�'�'���?*�y%lt����Ғ��mT�})��ҳl8�*�E1�0h8u�$��V5I�+f�A4����� ��!�o�� �����z����Ћ0C�rÆ9�ܕ���vh) �A��4+L1	@O9GGS�<�iD90MZ]����ã}+��ؓ��K@�vV0��^0���&x���cf��8� �r���#�uU�-��Yc^�ʵ�a���������1�͇����6��h���4��D���b7:����{/��h�z;�g'�ڋu���z6yh��$�X2̙P���f<����T.-����Q�O%{6��h�%|xc���d���LE�o�h/��Q��^xK�b�ꚌYj}.�Gml����3-�����t�0񥙠`z�N��y�x(v���)Y6������5B�^� ��'�j+�͕�	w��L��~V�)��pA����^�G�h8�;Y��Vnt�-C����x���C�����G<+ǳP�v�`3��� Z�t�ٓ��{K}�_��������X����_�*E�G�+��̲lb1�u��"�a<e�j��3芐��WQ�R7�`n�������踨%��E��V+A�&����h
px��%���U�<���[K�v�c�j)E�t%[����d��%�QN�O�݆O�sIk���6{�o�b
(��н3]�-v�'�R���
��=[�A�TkG�[�<z2������T֧�o%@�@�Qي`�~�q�L�O�arz�/���A�W��I
w�����k'K�}�܄<9�U��?��pbh���~ضGB����
8Wv^� 4��O�3�n����i�}��_���*[U���G��cK�e�� ���ap��3(A�LoZ��O�R��K���m�QN�aE����,�yab�gIQg�(;0�P�d$�ُ<���(���|nn*D,5I�V��{��Nہ����RTq��.�����3��-�=�Ӕ��klHʵ����|��4�{������2��疧��Q0��$�NO��b8F��9�&���C��Lq�ʝӓa�96��@F:;;�� b~P;|����Q`�"vT]p����@t�D}bhbpz��0(�EM���o����8m�q���yQ��Y���vhAX�	��/мw� #� I�i�lϳ���L�*@���0:�q��:UR8l��F��N|QV~<F���0�"���s�tb�юqS�3�f�R�P���H(#��.r��.��X�'����4F#��Gn�gmS%�n��
�n)��e� S<�w1��������KE7
����oT�������0C��Ѧءă��ݨP�%b��Խy<�ݙc��
3&Z^�zk��w�x��#�tSX1�̒��Ƹ[�k3�񩺜�=��ia��xu�zi�^�/�b��S�}�mxђ������H�p�Z�]�!�`Xv�őQ�dk����!It$�w�D���T+��܎�o��ٵ,8�V���Z繪ױ�z�Xap8�hY�!�z��%dy$,����&�>��7VXV~�lǜ�G���1o-!�3�F�3XT󋍞֍ !�VcC�ơ2���S��,��+�������S�ׁ
K���f�<F�Ϯy�0�&��
��=�x
U��|͚��eC}y:�����X���`�]�{Ƣk)�k��cАsf╒���B���7$�b�SHR	ƍ!��c�����+g�5��#�q�����k�O����ew�fYzm7C�;���*� ��P%�|�xx$2�Y)��<��X�oU�3'�|�0]΃<\����F�K�t���C�w@��ݒ�M�'������0��F���'9��)���w����p$�8���<ns�{�5i�R�='�6PRF@k(	`�� ��� �`�B��/p�+��D	����2�N�f�S���4*���	�n(�;^�籹b+��u�����ĻK�u"�4��a�2���0;��LA}���K���5hp�	�����$rL5������!�R��mp5|-��M:��R��å�.��R�I��ݒ�'A�o����\"��"������OZ?�?�I�Y��3�R�z6�_�jL#�u����~Q`�
�֍!1���ʹ�F)�MR����"7Q����'�1S����������N+x���'�T�ѓU,�aʔ��{���h���8�4�Tw���4�q
�z�oސ�I�é(�n�dkZf��LZa�^���������u��A��B+�������#Y	�m�w�g���Lq��9�/����H~I�(6�{O���H� `:�����ɟ�ɽ[|ÐǞ����Xڦ./1=�4���4y�qވI'�q��p��z�hu�R�A�!��=�wP?��맴@���Cs��m|���R���%p>M��LFW��٠-���Do��rpɿ��&{=MX`�8KǏ����wL*L�[^E�L��N�������Č9d]W�I\ȁ�7������(�f�c=?��P��&@�˪��-�mMV2f�
ڶ��e�[,e��G�C��1[g�s��G|.�i�����Å|��^Q�+�L�u��fb>�8�HH��m�4
ɯ�a��m�0%����v��l+0]�j�����c������1�"y�.��\�#�X�m�C�@���J�6"8Jq�^�л.�md����U=O��az�F;�g!��� �\4��XͽNP,o�uVa��m��*fLmK�9n(���Y��Lw�7a�V�&l��V2�>�8�7&~�b���#m���fɞ�d��Id��C��AM��* 86��n� y<���\hB���hM�Lݗ\����k)�l��IZX�w�r��\��� ��'m����*G�N6��p=.�+��(�o?+�s0���[39�\qa�F$���.Pw(N�^����c<`�k�-O>Qz�@iq3o�w#���:Qy�K�.ƾ� �"���A[Z*[�k8��X;���/ӽ����h�
�Rl�J��-�]�q�B�t�1	���E�;��,ml��Y�Z�	���y	A,�U�꜏���Ʒ���{�r�vݟ�?�]F��P��	�c�w�\�W�Vo�ᚶ~)���8n�4Iyar�7��h��cv~�ͻ��i����6`�̻�\�,व�[ؾeezv�V~�=�?�� x�j$�q�K�w努��$
�o�b��;($**U�|����0K�N��9>(�����cD��F�kzg��T�����w5�J"��vTp���5�3�]��\���l�<;<����aC��w:�3���"4ǿ��Y�4R�����c�����	G���� } �2�uI�~;���vXA�M�D��*6�����Eq�(�ɠ������b��u7�!{xQC2|s�6��r:����ǚ�M�	*���Q��#�Z|�>�9b�x� �x�YʒLe̬/'�`H�rL�*�`�p�>�w����6���k{��c-w��:D=�����F2�yʟR��$
IKa?Q-=צ�H|Q�"ܠ��#�ǈv#"_�*�s�i(3ٽZ���suG���Z�|�`��`!8D5�s�q���BU���q�6��	����7��/Q���ꅔ)��/��3z���`��;��̈�6w]�J�!�����������:~)�.;�U�ߓ����v9��V�n�QtW�!CDJ�q�ݮJ)����f�d�`gr�ao-����w�iBc�ȇ9�9lm��x~�m�A��+���սܥ M\�V�9gG����n�����L��0dVߙsQ�\!����?�Ҍ^�N��Z"s��N �������ְh{���]>�q%��͎��O4Q0W%��G�oٲğ"�
^����w*�ǬAMH�E0�]�	9��&)N� �ƎL#_1.����%Rw�)m��
z޿�~������?	��!��<j��0�a�B��ui���y��Ή�Q>����9D4#.{ۂ
L�6�
��`��I
{�f�����6�Ξa��E����	)�L*�3 2��u��`?�+{ejA�r
�
�O���1���P��w`�oo��L>���@�ޟ���+�ڢ;� yZ^��~�#�1&߭����v ���W��D��J�t���JU��x�g'O3�t��ht4�~���x�̸xOY���
p�k�7�:P�?�I����8�(
��٣+ˎ�P÷9_�E�9�,
����	��e2���(�~�5�ԧ��J.]%(lY8�[�cTl�E>]L�+U�Y鏶:���䎷έi����S��c�A$�>��n;�Ց�i3����vkv��QM81sT�P�f�KU�\=�Q�ȡ:�)������3����  ��]�x���`���;x����|�o�Nf��e�n�����|��{h�FOE{ �EIH�5^]��|@ ����x��^�`��y4�-gP8�1Cw�|b��0!��K�LN���E[(����X+�hU���Bz{[�i��pA8�{67^�fj��kW��=f.]����d���Z�*��9�0[g���ze����f/(�=�>!s��>�6!f��y�lj	�T^�c?M�ޔ{������$Q�V�/�<�A!Eqq~�6�����B��y	+[�EU��@=�����ɖ ��@Xj�G$!��(M��p�;���f�!��Bu�ȃ�8\m�����Nއ�"�%�t(XLy�%��)�כ�>Pv���~��N��NØ����z�V���j^�~i�dy�s	�S;P8yx�\�a�5��ܱ���j!�:�Lq�.S;�R]�fԂ��:�{~����&},�W�5����r%r��ߓ,��`
�G?���0L���Z��%P�C0Z�K�^��Q�Jf�-�ǁl�T�Ӆ�[w~~u��t0S��[�G �}l�5�]_H �m�Z�kk��ukM�:�|>�;��V��ֻ�|�Gt ��V����P������r��>nB��6���
n�{0�R"�x5
��;/���q͖Q���l��ae���|��N��sa���]I��/O�7�Z�B.��Z� �`��Z�m����Ud*@�+���C�)M���#��n>Ǥηh��k�X�5-�|�� 0,66N~|��DX��,�G5@Ѧ)A~U^�ٜ��F��c��0��s��x*1]Z��7z�+��;�;[m=�ش;�7�'���s�[��!�z�zGU���:��ޠ����pW/�b�>A�irH��>+7�<�t���:�_X��(K����#E����[�n��2(��ݵ�����'#ʼk�#kx��Зb6�-nU��:$'�ֽ�r`s�
�ΟpҼ�?��)�>��?~������[����=�*��èɒն"�HSGUg躑�y$\G_!y,a��� ��V����ds��y�T01!�b?�C��rA��tԈ�N���!r#iiC����3n"0r����Se��nve�b���o�g*�t��h5`�x���w�6��c��W�B�zN������6���֟����$�F�������t�+�Qa�:��D�T��b,rQ���N�kg�^:w&~��p���LM۱�����D�����kJ1��%�R���EnH
��hȫ7�ӓ��H�)�1��|(9'E��1�%�(yQ[��Y,Q���y���J��i��{�$Oe�hP2e
.�!|��D���N}kP@1���`s����"��ٺԃx�5�&7����d���ौ<��W؄de0�5���������6Ȁ좗]�d+���9ġV|%�����C�����9�2t>|��,��,m~-,y��:�H�1)���g�ԐJ_CҌ��s̅�<P`�1�Zx|�*+��_��7l>^��3M	��o�Y�E�M�̦A�{>��:ƤK�"@�$�w���C1� �R��͝od�V�?�-ľ#
i���J�d��������~�V͎呲���t��<>_-4�?��fm���&�E�X���p�}eMDj�Q�@�q���֘NȺ[��{2�	R�7X�α�nǗ0�>��c7��UD�ى	���Z̚���ԅh"r��I�e��Uiı&��?s��Q�����h���"z+;�����ʂs�7c�>���k�6��Y�_3n�5n���I�"n[��\��>F�~D��Ꙧ�y��f���;��F��v,�Yi�[�|`��Y�N	��s�Dw琶�=׃�%6	�?��2����F`y��Dh�7�:�d]�M��
4[8�_+I'�<��,|��5�Ck����4 �<�LRg�'Ů�Gp4۸�`A�	���Q��
�p|Յ���j���%����>
��al�E�y�,E�F	)��nu=A%@g1��C�m�P���%���D985\�Ax�~�j��F�>�k4�n��/�?<����5"✽f���[2/�'Q�SJ_���Z����\!3�J-c�����A#��h�֒8��+S���.!^��R���2Z�6N.��͑y/w�>��}>��oE�)�N$�S�;��="� ^��v��/3���Nޗi0�E �	n�~�"Gm���Ξ�s�������	FmGY�E����؟�F�-c�$��~�,@/W��^�q�N��ʑ�{9{�X LR�s��'P��i5�/7x� �6'm7P\$>v��\5�d�qQb���"=�o���gг/EneB�Q�@���_�<ji�N��-p'���/A�5�+Ҩ�?��+,�C�c6��c�t~���:���