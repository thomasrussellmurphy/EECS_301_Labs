��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|>�qT��>���r���s�#gcM"�.�a�w���H+��쥬����o��<�aR�����|��*�w>��6[�q�>9m�oOM:*����;�*�YI�O�뱦3E����N�,��S9G�I4!ς�j�s��J�=��l�������}���,���c#l�T�or�_� 5i����)����X�D|��L�7����׵�������T�y�KW�]��t$��Q}�$NU�Ժ�P���z�N�z<�G$�r
1�i�;�I�\~���1d8A��7�i����WxB~�O���0�!���Q�8�(AZ}��tB��2��#q�$
`�Y-}3Ĕ������PUA�ީ�"�lk��T8c�s8��++'�m012���LU����2j>Ԩ���mObY���z^ x��!����ˈ,�$��R����(��Y�I�@b�/44;Ú��5�%"�Tp���M4�>�c�l_`o)xCsT
�C˫q�V���\���&s���$����k�/��0ch���??�:Y��DG ��	�.X���n�-��MK�&L"GK�i0�$�,�π6��~�����܏��y0/W[�}�q�27��6)|�ew��?�T'�y����q֝�7-�>7�y��-�vC<R�9����C1�Ǫ+�TH}�Q
]ot>T���-4h�U�B��̟j�D1&ŉ)=>��KQ��(;���rA�P9�;qܵ�_�k[5�u����Y#�^D�GD�������)g��ڙ����>*�h��쇜	.ڞwO��1J��Rh57����%W��,!�1L�n�V�}PG4�5��7�]"<���WՒ�zI���p�4i��T�-���e�� �Q���G��;� ˸.���8�xT,�| �Q�4G�a�M#R�Q*F����@Nеֶr��Ӿ;���|��$��)��oPh���\��˒��+My� s�����]��}�5��A����"RdOA.�E4�[�XD� !ŀ�0�gH�F���Gk� �h��M�~��lH�L�Mi�� s�z]� ﳱٟ�"Q"J���SP�+�_�rI�ʎc?���h����):�>\_~h��;&�n9R+�����_�uJ�@�'I<�5
^f��`lu�?h^8[�u7waF�ݕ�c�W[v}J��~/ˑ��Tꃿ��裗´Q�଍�ff(�S&��sF!�~�>T���|���*��\��3b���{̆e9�<N`��L���^r�I��z�7Q��� 7��[�I;|l]�zɮU��.�/t�L��$ne�3*BKjfՁ%��c��T��B3��E�����W�+
-��Fb�6Y���@G�vJ4��1[�Y�y!Y�[�~�`��*Æ�Ng�X&�6Y�Y��&��L�=ػ�J3x'Q�I�_��<���5s"]ߡ.�d�e8U*���W��fQ,������HM��%k�u8���v.m*�����z��,ı�=!^]B+�%�Yq9�lq�����P�%!�?A�C�K��O�K���m �*��9j����I6Vn^_�u��L,�+ֱ�Yׅ�(�FQ]mn���{�дD�x��;!j�J��t$;�$�{��+���H]y!�(ږ�q���^�9�����q�Q|�� N��N2Q�1vqp!ğj�Vuuh^u��ѱ-��eۡ���.ס��Jj�c�|�f���C��d��&*(�X
�Χ(���*���V��qvŧ��\q,�{��"�(;��Ff,�ds3j�(|�����5�Q8H����������B�x�[ݸ��Y���|�� �� �g�)FS�M� �3J�a�#+>:��0D|���1&�H���;�Y���Kg#��ZT�{��r�݃z������ y�Ռ�<�ښ�5��jr�<AJ5n(���@_G�O��:.�H�$6f)�ZS��j�'{�?§}�!���O�I��&�/����9TP��� ��eEgs�D�o�����v�1�����5���4Pz~#�7��~Q|��bj�Sn����^��Lx�X���!s[�{�D[�{�@.����j�����Z2�P��[Ť!�T��F����ڶH�}/��E���p.ħ�j �^Ar��
�A|��.���|��%=�G�e/�lIr�����$:x�붖��z��l�=_P�Àl��JLu��̓l�c�\�ogژ��c÷������#R8�DO����ձ���P�o0�u~0D��J���U�G�)l��B����M�-$�W�[��ҋp<UV�g���ˮ!�����fe�:X�Vד>DJ��m8C�G�����{�*����T����9��Z�]b��݊.�CZ�`����ܢ��O��N
������x��q�Z)��o�b,L"h3�00ꭼiK��s���WԂ�����B�d�ɪ�&A�bI̵4�'�E���N���|U�@���"s7�6���	��V��H�ZZ�(?Ϭ�9�FW�z��rr�E���[���Z���J�h�gՏ����ǳ���JHa������������;�h�%;y�q�梻[0��N�[A���Wu�s,�*�B�*��t�P���	�ԏ)CR4�mgCqcإ1�o��HF$�Ӝ�N�G?�A��ɜ%&_�K��V��g��
`���{_$`�ň�����9�,��ٍ-�{I�YT���I��"'U	^<12��ٶ����w���'��;]�,c�g���~���C�4�Fe�wûH(�S�p�K��?�2�=�ku��'��Ө�Q�ݏ�3�Ch�5u��}����4�u�H��:��>!���ν���s�̐��qjYOQ��%�-�BP��MEQ�s���ҝ���^��g� ��ގ@I)4K�����W�����BW��{�L�82�HL�A�bZ̉S��z�?\�!k(?&	�8����GҀ(Hm(!��y�����F*"R�}WV�����߼J|����Bb<_����?�Q�\Tɰ�؛�5����.�	�1���@�w��h�Q'v�wi]�{CN���|#�N��fN��N����S�V�L�a�Lxl����t1�*U㶩`=�zSm4ٞ9�o���X�\�#~�T�}�,�3�t�D_�jc{�4J�3@m��M��0�V�v�R,`�{�Z�/OKRn'A�5����0w�n��
4����['�.��2f�u	60��4+;ך������C�H�rSȳ�n��*$�;��P)�m4<>��V�̘�[���F�<�"�^�_X^ӞW�A��N��_�N6[�\�|%=�����_�E$:�t[��4|vP0D&X�_�TL�<�ǉP6I�x�#zq�ـ�S�w� �,,��4gN�&���7ҹ����xȰu��+A0�ߑ{:��"-;�*����	��J�`^{����.z��t?P� ��`�������E�`i�|˂�b�Y�����Ec��Ey�����E�5��U.���0^��,��YrD�&��*��iY�t	��}Jbc�1�R>/g\֡���A�A�҃N��.f�sC��ު���r�!g��jB�ĉ}�|�;�D��F�yې��	�^=Dj�>($SD�Ű���2���45li�C���)߆7��C���S"��J�՝=iR��%B�,��Fl?�y(6$dO�*OV��cE�D@���uQ[O�5�����2�-$�a���ZĀq�i��+{w��L�V{�MrN�r�~�N{��U4�Ӆ���e�	��
��w�6����Z[
�����t�3S��VT�%`��~�`�� ��c8�P��Eڜ�I�����Ẁ`�k�f?��g>�/��[j�a�J;�ے����x���aOZ:��fU���#r��