��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�i��a
Α1S%� �uj?�L�3��TLei-3^5]E�$���zlUG�4�q�W3��I�i�bV�`���Yl Z~�sƵ$�a�m�X�/ p�f$����B�I��Փ���"l��v��~�A�mu�Ű⧘����V�8�g�iM^���7oT|g �����JLc���p���_��Ԝ���F����+2*z����n��;����p��J�Q���$�=ks�v�ݡ�_�ɓH�ɲg�a$�6�=�p�҂-I�/������U��c�p��`"Z>��V0���� ky(SJR�'�4g~;����@q���mY��`(������Z[C|�*A{+�˧G��42@������M�l�(;���V�@�"����g3�,�W�wP���
�1^Vhs�Z��z�h�e�s�����������[��{Z���q�����Vp\���-u\[��g�"���G�6�Yl�	�z5'�~)���=}3H��F��t��y���r�E:gU�H*Q�y�f���Jy�uG{���[ȳ�"{�AT�����C�WG��t������y�ԧm��=8��.O�ԁ[cj-�����`�-�����#\�����4�:�^O�C8�a$H�)��&F��D�`$���Ѽ�A*��@��J��	�wS�@��Һה��B����0Ci�tנ)q�>\�D
���w����~�Z�T1�� ��L�M |�@�l��?�?��^K�J6��4LjS<����!d��(@r����=7���Å8԰����+,V��%����gm�A�0��o��X�45���`.�~���i��C�H~�n���ҋ�^�N�&�ա�D��'�����	�Eӛ]�#c�����H�����
�/5�J0�$�����3]`��),~8})�8�y���G�D
F�����^GxQ�>���).&7hƕa�%�Ԗ��`1(���'5��>��>ӏ�=M��[�d88^��E\�isG�ՙ��]9�e���?����_���w��Kt�6���^��c��6�(jsqx��ۣ�#Y�����ّ�m�|�@Y" VL�
7�5S �)���"����ò�'��a�Vvʸ[���W�Y�e�{#��'��GۤD��BÀ��<�|~X�j����Z��o��GG����)^-|�0������Y�U���p�X��l/e��a�9��G����Cf�q��'C�y���c�^Tu�ӫ��E�Z���$Q92/r���9�@�a��i.����ߺ�{��;�/?���Z������>����fMw�s>A�HF�G
N�=�K�:��qy�K��d�Ph8`F���YG>�5꘳�����)VmX��椌��Û3Kz��ubK�oNꡗ����z���1����9�w��a�P��7���K>yd�W�[q_Q��ڟ�(��D�mny��J��[���9�"��զ�U����Z|���Ge�"�������pG� ʈ�q<[�cI�@�н�v:����R��`�K��|཭u�%�ra,Z!{�sU�v`]�?�y|��|�P�a�D+U�f���Yr����5,��I(_i^��fZ����Ɖ�f�g��vH��[��Sɱ�6�Q
:߃�h5r)/����i��Ac�E��^�R���\u@��ZE�/f��!G��;��V���R�M٩���m&R=:E/�fu�O���8��ulE�@	Ãu�Q���G�W��T����Lπ���-�� �3�[�&X5\�1Fص�`����I�bZ�5�3_��%������N���u�Ǩ3#EÝ^k�Z�:�L)�����W֡��H�ኣ-x�eQ(,���:y�����moa����E̸$kKD']�;��S�W��/b�N3I~���ӄ���T�`E5��P�AW�����՚������G���<1l�N�8�l�G�E�h�V��C���	����E�}[c�C=�۔ w2LΪ�KG��`�zT?�2�	���`�Zcz���D�%�o�}8�d���j�O��V���ha��_��@���%�T�2}i���g�vd���|��(ٚ���|���F���=���p%T?�"A��� ���uw�*Ē������	�̽mK����#�Z�)L]���}�Ҥn=6�A��g�&,�*���v�/m|���%�����uЛ@7ΠJ�E��}qG��x#H��I颖+�%��A���r�(k�=*�C|�y��Ԁ��b!H���t��7f��K�?�H�M'����V�G���-���n�c��O�6�g+=�i�~�聍�'�J�O��!\��L�Tb�h8���#�L	B�s�ڊ�G�x6�X�Z��@��`��h���s��ݻ�>�"��r��LqeLU���ˡߌ_s���;��Ix5�ѫ�⥜�yK�+9:j��2���&z�q���4R���=��c���c�7��	Zh1S�������W�8����M�+r>+�&r��e���O�J����M����-��9JI�2�p�w��>v�!۲�o��p%S�&h�5Ք5pf�Bmh<f�2�NiBV��_M8#�:��K"���`�M��GA��c�d�)�����I���z׳;Y]A�jُ��{�K���K>�Ϗ^��LrWAO@�_���0�C�y����t[�]k��j�w"�Q�ҧ�8�DQ=����a�Ҷ�$߾�F����	߮H_C���g���$u�x��B�k����\�Q�!�E+�=�6�yY^��풖g	MA"��r�{��S� \��(�� ��`�spW�P�Dm���(	}b��5�K~��_u���b�J���a-���W�KcCt�)�i.A�'%�ޓ�%�F1󷬲i��3E�+��R|�s��v�|��S3�����8Ce5ho2��j��~!sޠ&�v�u�T���y�u����[J
 ���s���Zt���`z�f�#s�
�R_.�gw�f��+�����OL��S��y� �j��݀UW2�0ƹ2��J��:�!׬��DG@q�]�)�1~���O��aب��+0w9� �73�@2�����p��G�x�}̕TK[5OW-@'> �Q4��p�h���a�pV�2p��y1f����[�]��1j3D��:풅���m��Aa�d9L��΄��×�%�
�+"f������FY�M�3��S���)������it����O����~t���_o�0��֖����{�[�G ��NP�ps1**�����_��6��"�"a���ʈ'��X�_��Տ���Y(���"���]�+ذS�3<6~X��|�'�Lp=HI��h����&y[�tK�>�dq��� wn�e�m(:��?����1<%�w)ha%kv;�fS�C�b* ��+��n;��&�ŀTv�N>�T	ppo�$�Ic���/��[އ�K�x�@�56�9F����Q��?�a���l�l��y�2�P�g)-�P��nΦA �)F|��w��[Js��4;�lvj551;<��U�$������-D�0�|A�ZL�s1��0�aVJ�p+��<��Gl��a��a�X�S%G?De��d�MO#"��'�
Eƨr��+�E���;�/��&�l~���(�~q �o�h���R�ٻ�UA%^���7�]���p7s�ޑ])ja��q@��u�qV�S�oV6'TѪD��� w&Q;�c�`�zv&�!�An�� w����7��АѪ���~(;��0j��� �*
��#����>�D�$cK���y|Z����X�������(�b��uI�9��g��>��Ţ�B��F,Bq�Qv�o&�h���W�b�h���n��M\�����@���Ы�Jp�(�U����`�ي���e���C��H�����WLU	����}B�М���$U�I$
����Z5��h�Oi�R������q�� X�܁��v5���_vV�8����.�IЇaL�V^aH�.�=8%��)�S���� ��"D�aa�M���;�����r�,&���R	��zy�ҘKI
�=��*Nʷy1fY�;�J�l��%�s��P�$h����x/O��捻6����kW���[�Y���B?!Cj(��O��m�f�&@S�|W��2��5$d���������p�#��/-�2�S���À�{�)��Qq��Yz�k}�w�P��a�k|=��َ;#$Q��4�"�����@Tx�ijm�������#�V�L����9��1�2��	-�\����%���RǪ4t��Ύ�a0��4��a/���YM���@ �bt�GV�O�!�A���8nUO 
�6S���{hװ��pں"�u>�_1Sc >�5)u�%Y5�8Z�3�:�F�*��:kN�iy��=]N��	��_�1�e`��w�!�[t@���lO�m���Ei��W�����~���"�鷥̒�T�����~GP������j���yN�M��3k�Ą�+�l���+4˩��J=@�m��D2���������z�ǫE��gcӣs~�N��fb����S�t�q��]9,V�pB�2�1�Γ��8�R��|������\@�hR^�� �mk�7�$��C�=A&2y�o)�����O�9�ȇ��NK
�ò���>che����Vr�6��ʪY�!���
W]�7�{#�#����Ff ��
�Z��d�f1@�Ֆ+�u�0���U�8,��щ%�2"��vV���� ���j綌:�H/X�2[Y���*����{L��g�QEV�P��2��g�;�k���]�}"�Ym�M�2y�`��/Cń���vӓ�s�q��a�!,t�}.�*{(�m�\�9��hL�H���%���g�����S�Ϋ<RuCF�����eJ'5������qby���@9���x���sPV�>#�Q'G���#��@�g�é��.u����juI�`��C�d�m�"w>��1=�U^����v'��[�-gd~G@��$k-�h/����/v�8b�ﲖ��[��NX��ddO"劸1|��,Y�Ѭ��-�6�l��s[��ػV���n��WBF�T�� [�yz���S%�<���CO�w1�.܌�|�`D	1?�"�x>VT��µ�@�����=:q@c���d1�$�h�+��B>u��4�|��k�����sb:kK/�v�L���h����F�J&!���>��'o%�ى�rM�4��}�U�#�1~W�U�_7_|b�:��BיV�������x��]p4i8ޔ6e�N���Th����պ��L�i���"��YB���M�Ĭ�\��3�؇�#��/Lq~0r���EQ�P�h�4S�x�7�\�1:q��A������Z�%1)la���D{QYu����-��L��0Z�^}���K�Aa�H�������u����i�D*<;��(�^ �/�h�(ҙ��P��}ԋ0�o�MI�, yZ虞��[a��P�CF���@&��\3�d_;M���M��l�S�/oD�!\d��������;զ`;Q��R������E&�"����ެ98���T�/��Ű���
 �����	�!��Ԅ�L�����B�=���#�C�ޕ�{Gm�,����w9(;Ha�| ����T��<��rB�4���5ִm3�� �Gk�sdwD?����1�cofy���3#?�wE�x~����G��o��z�-�;H����p)U���q]ʕQ�M2��xQ�8I|��}�~��Ԃ�,fl`�J�VQ�c��>�%�1���Dnc?F���}N�?����@�q�t	w|y��ʝ�#Wc�N �` ��U�|�G��	����s�FV1*�	A$���=�seo���w���3��'����,�rF��*�zޑˁ��(`�mw ��_�C��0{!����.0�[K�r��I�L8�9*�:����:�
��=y�J��
�R�8������O1�4��z -�\Zd��Z[�����[C�D�½}R�Ko��bDг ͐��-CoH�&�H�{��I��h�D,���` �R_L�T�zz.�R�Gi`@������X����{W�k��/�=v�ȽX���&��,"��Pӕ������ݝú�!�Y�C?gN�ʾ� '��z�#�e��ƕ�0��ҟ�9��r#y7����N��/��J?��n9���������u�驍���v����Q����0��� �-W,���$KG����@G(o��H2|j{�L*��,h	냊s�P�
��=h0u��� 2.`IU	W�U3�G�)��|w�*=)��/ffS�0"s��xw^��e�=6&a���.��W��s�D�V2{�w ��|Ѩ�lk�G�*�
�tt�h����M�7v2�+�����_E�KlG瞨�b�"�������Zyd!��U���8�C��8��X³�g\��K(D枰�pp��Gtr5>���!r�P0Q$�&��Vj;{�ݺ���
d҆�j"z��f?)6�1����7����� 7��yԐ�R	$=� ���i:5��ڎ^��E}e6x��a�Q���5B߷�i��c�6��������[u鎒y'Q��t���I=�.�v�&|���pb�u�jՊ$��:<��֔uR���}�P��&����}?�w	k[���$�f������h�{m�%���q�%9�M��yS=�r�z�R����
ܙ�c�鷨^7�֫ҳ���c웲�M��Ij��cw��T݇Jv�T�J�2+$���$��╪q�X���%DK}��o{�y�}գ�E���)b��*L#�%x�Z�K�����H�i���0u\:w3	�e$V�vQ�'�OCVp�Ư��y�_Ϊ��g�ɒ�9�eLi�)Y�TDn�EO�at�fSC��௩`l��d)�O���G��nY](��3�}���K�o!g)9�A������W;���)F�yD����+�k�W�Y�bL �d��~�wKn��n�._е��#��~����i+�"!�$�������1
�RPêr���%������	<򪖀:x�i�;Ja��|��o��"�:�x��������h3;E�VEE�Β�|F�)��Oq���7�R{3����z�N���8�7(��2�2F�Gl=�!���c���[�e�
�����G���ic�vM7�3@�	b#r ����D爳�+��PP�c��Tj�.���cNE�E�%�ܖl֖㧅~���Y��8-�A�2��`�t�|�ϐE�@^\ĩ�s�$����}�#hֵM�A��$����|>�c��0Ln=T��� �Im<nA���Tz���x��Վѿ�͛���4:�eZ�@8(����2̷����=�3�ɺk�zV�* lE�rvA����H����fe������͐�N��ˍ�a]�)B&Y� ʼ������"o(���baZW�����9��4�׋jA��sN�o���V�/��&���X@�꧑����m��=�"kW�X����1*�CY�ug��#�!	
V���is2)�p0��3My�n���G�ťZcO'UH�28,���W�]�g8ȭ�3���_��'{��u��( N�� �D���pՠ!&~s@r)��{��Qغ)�P7?�{��<t��$Kc�����7˓���N�i]�KҊ�-F˱�>LWM�6*-����p�y���<AȠj?Z0�%�8�}"_�9b���{c FF��=.���x#��3�:�=�:�3�E���5V�NB�).s�!@w�������9B�~�+��I�JP���3��!�;��\"*��og9GG�$WY�O�xK�P��;�p��[g���&���z�wb��xx#���6�%	��K�0��t�l������h#$�#g�Ph�ke��R�����Iv(g�{��;�Bu����B�I.�$�4�+��Źr��@���@JŗO�@ؒYU�(����i���[Eigid�v��:��e8h��3z�9]XN�+^��!r^��@s�!��9(����X;p������;�"��n���y��� gZm8�q5x�Q�5C.�D��G���"����l���F?�S4�?�
q̨����pk��l���r����8�����m�Ę(T�%�������	'0  ��'Lhkt ��.�/�W�O�8��O�։h���m�Q�\���*!��X��h�:ĳ�sNK�T��5b���@�y�Uf!�2��VW����/�Ch�p�g r2C���PH���[A���B�/��'���ze"�F54ɞ�p%$~;�/���
 ��o��W]������<��c�1������_�2�ɖeA���F���*?���t���ɠ�JCi�Tn:��ry90H�1^��H#�����ԧ|�ƃA�32(Ç�u4���^_T�v8��۰��;a�mh���x��T18���S��x�͍���P�2��*0YrP3�Zp,�r�G3[�>C�3�ף�e]Rb����fhw'u� �O��7M��Ὧ2��ZQ�U6ţ�|��c_���ok�0�ip��*��5�?���X���@蚝B��d>��G�8�L��Xy�������Y��<:���9�Ȫb�0�/���W��x�I����ɓ"إӜ֓)�/�����C( p�.$��SE�f��5X<��ZL0���y!�����'���vObfg~�԰pt��7G���ne>��a�י�UӼhcm�P��瞮�4��I)X��v�8�_�RM�&����ʴ�4�jD��#7^K��%FlL����ۯ&�a��%) �`7SJ<�����<ڨ�o�y��D��P~oa^O����G�����&��&�4좮���������K��'
�����Q�jR!,TE��d0jYb��=��>)�,�/�"���*��]�f�ůڵy#jKCV�nn�͈<�]�p4�de�8H�"�n�,*�ⴝ<'�������j�蹼�_�9}'��4��4�f���(�'�=��'�5-�+�O}hx�ܡ�^B1���E
];ky���A�ƿ���=�B3�Oy��$���Q;�Vuْw�m��mDh�\�<a�!6 <�z��(�]�W���~7��7�GYe�ٛd@�	��E����;j�-��(��eQ������L�|Y.�%��@����6;YXUH���[K��&���}�l�,�6trgI�`�H��*:�P1���ծ4�h��!�^��8V��������:WjY)�/,\}�@��#5ؕ�M�p�VY)i�k!�䝯?L~�6��)a��]@#A1⸎C&Gޠ �`�V���4��?�`����~��$�mU��J m�t�,G�n�-�|9R��w/.M�=�3�'��Mi�7O�a��tV���^���-H7�G�e��Z�v�Xi�GV"�x~��q<�$爮޼E�|��)G�{�r�����C�-�-��aY*Wd
���bb߽m�Aط�Q�r�[[/�m0���f!���Z����尼V�oJ��
si�����3P(~(�l?���S���!���0X����k�К=�B��c�fU��nR��d�0u	<����	<��Ҏ���\֦�_i3j��Ėf�:y@���QV��J"�'�>����i0ǥ��#��]�U�L�l�V�C/�3��qC��������]؈�.@��k1�[<]�iê^�P�0M[��)CP���:-k�E�;
�^
O�����{��lj��N@�F)qy�)\���_���������*�Ӿ���wm����7&�OJq�t-�����WP�\�#l�
�y:ML}���7n5F�Ɯz��Lf�Mv^�w�e�v5�Ow��3^���5��E��N/�?L��#�������[�V �,w<iJ��@>a�S}��$�&�&cI�� �C�>�muQ�]ׅ�j���*+G�O���G���$tOW�L�|�eڟ�/�eI�����)�ב����qZЧ� ��s.ԛM>�Sip�Kݿ���aװw��q�5�~?F��g�;r�B
L��0��]��3�5�o���	�P�u.|1�����Xщj)7�6��l���K�B����NFh�)�㊍ͣ1��+`L�`��{@0=U 2j�B۸G�02�z���R�/�;�8�]o��A���`�MJ�i�
>ӏ���b�7i���h��|"$�z���K����mt�0s	��5U�T���vr�W=�%/�)�n���ñ[<'��h,%��ms$�m��4>@^�G��Rv�;2����HY�J4YY�`sܫBk��Հ|��.֤�{����~,3��I,;w��K,�/��c��Ej����m�*AV�ln7vr��m���)�gԻ���)3��p�9�S,�qD|�L�ӵ]i�U1�Y�����b��x�磕���3��)��K��;�F��1����Hy�lDXr�T�ݪ5��e0����r���\_�4�]���+��u|B��$?��6�n�I:Y�@��9�A�&b�À$��ɫꩺ�F�*?��3ݠ�'|Ε�}��*����Β��#Z���0��!a�H�!=����s����Ζuk	�&�PG�7�L�0$j�wNJk�$��1�Kc�E�y�^.K�\��L?c���4͓k��������q��̉7���������v
�KT=5W���F��:���\����ˏ�p�/\�����W���]\%v"ěM�%��t����HC�>,@i��)Jb�U=r��R6�+�٠����2�pu�&���?~:|������|~W\{�y (�t7�����S/�S�=,�s|ua_��X�I⥩���$�1��ug�����v�ܖ�?�Um���K1�#��A���=�G�*�߷�Y�Ȫ�A�`]����/̲�`���� �Hz5�hH)�rd����ʉ��:�i�d$��-��`=+��F"t�¯���u����|G�QP2�"L4Dy���2��*�ʵ�<���ܖ>6~~aeI�t�WI���i��9��U|W�ŝv-��\��S8 *p�m�W�����k�$lc9d�'�`k����w.5zU����c�?���E6���/+�&~˳j&�$aIe����m�����4 m�R\����t?���	n��+7��`��؜�N���:� �� �F54�-9`� iHMX����ZSF�~ 1�+x��5K�o6��b(��4�A\�0����V���[��\��"4#)*��\������>�d��!���n֌����ۮ
R�WM���1$��Х�ē5]ч<�K^����{�2.�͂�j��n������J�>�8��EO��#�
7AF�W����'��杋��xt��ϯw�)�i��㼊�,��;;��,Gx�m� NB�x�9����$"�
��9��8��������<(�� �h�Sv�3� ̏�h�ƿ����>6p��ܔ��q\���	�C��G�F�	�A����&컉��W�r�J@N��2��N�|7��m��B;.�E�c��Z���p�3Y��;���1�G3�9%��k���ltq���󬓷!`A�uV{1�U�~ֳzk�����^�yնC�K|���ϓQi&��2����3-�����k��ҢK��J�����Ñ�9�<6����J�m5+����aC�d|�븦-Qm_`���*3�h��L9|TK��'w~~��ަ�P�|���sx�?��˴�d�[���靆��9R�t���|�F7������t���1����A���k�t���Y!J���k����A��㡛�@���*������pyI�
�S��(ǹ���1��/��ǲ�%����,-CzKTi��33�2�_���,�����*_z�#U�n�w:U(7vO�'�k�~t��ܡ�ĮZ^b�zH��-��r�hG�"h���CAef����c��Ma �to�*���Xd(�{��~�\n�v�3�f�c�3[�=8V�O����	Ѹhe����)(l4Թ�X���f�F��{?�^�Tx��?a�02�yBd��!�#��x��X2�
�e,� [74T��sw�g��Ԅ���kގ-h$�2N���8�O�w'k`�FD]�&7")O�B�9A�!�PX�`2�\��h?�u�ӌ�]���4��fV�=Wl2��P͕��rn���7�f����A���t24��+�L
���U��2��e|L'Âd�/�N�
O�����2��+45���VեrG���S��YX�W�%1.�9}bC���� ��6x@QM'�3����h�`m���)e��,lq���=9�F[;
��Ϣ���U=��W�ءf�򎺻�ԑ=��#]z��婅B�^x�n񸨸[Tԥ���?	�q+�;=��u�"Ÿr�ק�߄�]C\��fZ�!'xrrȎA���c��:�<�u�Z�/p����_[~ ��2=L`AYq���5�Z��`��6��U���W]��!O���& �1)����X��N�6(Lu��������{�vĔaN?�Ȋ)�p�6�B���0����7�{pEXR�M��2£����G���~��e:�?Rf>�Q�}B�Qy9턈Ο-���=tQ)z:�������ϺƦ���Pq)S|�\��f�zm���'t ��"��zw�ۼ"I�gf��w�C�0L�w��a���'�E���|�t�KQpDh�t�l<�$:��F�%X� W�,d��ӄ������N9s��n�#��=��pT�f9�fA�'c�m	@'}v����S����!q���r5�4��G�W5BvPv�F+��e���7(H����TŖ{��db �Uq�L3���-9-KТ�!�W_��!I�0B�kҷa��wT�v9M 5]* |t�F'y�jqS<����Lc�lF�|�;�ݴ�d�/Ä�;3�����ä�c��)-l{)\k�y��,ZPƤ�}�ğ�����%�! ����(�o�^%���y\�"�8�Wd-��� {�V K�>���>�V'�J�N�1K)� ��m*1%)ޕp��lͰ:����������gXi�[��X������̚.{�T���2���?&"
ad4�4}
���p��=��|C���$X�3PG?1^�!�h�t+.���S�1�c�q���R�t>WRm;��؍z�'�O���¬�6����;H��yl�p%�ek���ej������԰�B��_G.A��}�ύ:�	�}� ,r� d����%%b�
C�S��kd����%��8�޽.<n��;2o�r)�.8S�{�V��Z�D�;98(��E��)�wp�r����e(��t�i�5��b�uq )� ��4�l�K������3�����j�7a��l��L�S!��R��$ >�
{�4��!V\]�80��a �53����?$-{[�|���3}b���*�e��X!��c�po�R�(��������݄ٕ�%,H�:t�=�L�tw���ɜ�P�s�*!�u��lI�5L��܅_st�e|j���v����2�^�d�+()��4���CF�7��S�U���UG��h��r�<�i��@t�������.����
�E����Ql\�s�
ϩu>�܍��GՄ/*`"�&�.3��	-
4S�IL�>(^]_�jAn�6��и�18�����[7}R�PF:����#H���ja_���x{fP���'��/5�S��	���&�\���O�C�ܱ՝�,��a*xI�kMt,�X,��4����������:V��&1��K�6��(��[N�� o"��|		}���a�:���?7h��� n�.K��s� �u�δ�b �����lB��������u��j+ȍ/4ݐ�R��%h�o*��E@e\:���D3��`���`�O$5��>�� D���*f���;����Y�`}AJA,���;�n�8�UN,tĥ0^}��8%6�;�@M��/N�V���e�X�1\s��#�`sx�������4؃])��P$^�v�b�<%M�����C��f��7za�z�bc�Q�,�"�ٳ=�ni���+#D0���s2��(#��t&� ���\���hY
a6���(�{0Q��� �,J��0�Vrf(��fS�� c�4�I��D���t�4��3^�5Z���)���+�u����H�ܑ蘒� ��H:1݈�G$#2V˿�-y��eU��+��^A �ɺ�����N�F;_M�'�H�������<sg&P;�9F����7P�
Q��f�]��2����= :��$j�鍃�R�W2M&�ae_�l��7�+�Q��4e[-H�6ڜZ춾�ί�<���<3���&���=0�N*8��������I�ǯ�:nukOZ��@sW;���d���i*`��u�{u����������U�^����k�.�AY�$rjl����O}JT��{n
>�7�{��8b7�a��9�؛���en$?x�]����:g\�Ga�ތ��`rpvm�M;��[ (��k0~p��Naǎ�v��� {ۙr�L������_���������=#L�5r�����s��f�-��0��nȚ4���
S�ʉN�����L^�����W�q��k�Ѩ����j�UI/�:��<I�	��<3���~ Q.ߖBM�"��?ۼ8� �Z~+�k�ǒ�������_��:������rЭ��a��y��>�+�.MJtGඪ��U@�L:�3�m5����6D�^���z݉��oZ⏊�ĲR [����l�h_j��0IQ^a.��ղ<�Q\�k|�^�=���Z���6�URp���t��sA��q���<�%"^���$�~ 8����F96���4g�vy���O��a�������f�A(��b�3_hz�1��J��`����� ��br���VW��e��F����%�[�F��א=q���ɖ�������z���&(�9���)
�Y��l]�,n���:���gsb�c��Ϭ$!���y#�K�"!��)�y�1z�����[,0݀���֌�% LmA<�/����lI�H)�yщ&ۤ�j�z���yX�e��%�A�O��\��Nꓯ�� 揍���߄óVJ�L�v�N�!�َ�l`�Rb7�f\�4UW,-���pG5�?���( ���i;��g����|��P���`��z�`1���,jeaF�sHkՈ&�i654�=^v��g	�$�� �g�<�&�id]���T�8�v;��.\_x%,���7��A���`h���N:	�@D��4We0:��D�dJ/L��HKx�Z��р�����H���"v�ڇt/h��Q7	��.{C�"�
�Ԡ�Q�_3�,�F��3�k��g����Fg��a��\�Q@� ��Inoԛ��Y�A�%ҺVK�lq�ؗ�����AW��DC}�������嵀ZSݨ��N��֖����èK�xF�(p�C]��-G_1B����/f#I�>�WG���>=T>k�+z}�����;>�{��v�<�����kL��s{b��4���ub|����[��~����T�$�1LI[��m�Vo��$Zr%�yY1�[�S�̈��Da���pE��'���4��m�S6�-U�8���}��)�P[6�-��h��S���K/�dy�ke6W���]���W>��fPݴ���< ����GOK�"�;�ɂ��_�Xu��G�J�O�߹���'��-0�A��}�C�d��j���:_�%{��mJ��:�h�`��	��«Wh�T[� �]����g/���N%lZ���q�ĳ{�Y�=��*Zs�A����q֭��S�}�]�T���ns��I�!�����;J�9�q=��wG�f����N=$�}# [t}~lr�qS�&����Vno3C�˝ܳ��� �� ���e�P��.�VW<�!; Pn����)�O��f��M� �%q�k̜�?c�7����V-Gu��œx���K�m��@9!!꒑�8Rw�0azMd��H�X�'�k�[���qJ���6a�&�	:��_r��+�V���:R�v�X�ᙒK������;����oB��rO�]��5�Y��h�+�lwGv�d�sAB7aX��r�o�`G'�I�w1�M��޴��C�0L�F�6K��,֏j�9�����|��>�(����nF)xvo��n<��w�c�
2�V�R^����؎�o7�*M���Б%%�
�~��֕ΐޠ�p� ]u�ظ'�D�ӂ; �{Y�X��_�w�T��5J�yh�4��Gځ&�q��MY^^��@XYڵ��>����^n��h]qs��y��J^k�I>8�%U�x*͘M�yHI'�zbj�\?�h޵.��W�mbg��`,\���0�u>1BK��O?r|(eԑ��r��MB����o��"�wXāg���l��Ψ#e'OC���0�;�����X��dU	@?�(�@�9{|�P��y�	�]��v��~��o���ZT�zn����� ���٨t�vmd�-��P(�+�<�Kl�O�4B-��ˈ֦��.�����)�z!G�8�q���N�>�`�\pC3DV�b��jߜ/��I-�Ʊ���֩=��Z�E����5J���yAw��Ԑ���!+���ji�ί�J� k>�a`Z�5?�i�ǩc�����(d�"oנ^}Hh'3(�5_��]�{�}x�����T�$�M�m?��ߒ�'b��1��D�3�'�x�N�l�a�[i�;Ѕ,F��+� ۉ�U
��!n�R�H��j�L�����SAU��/G���d���F(C[1�){{dP�	�5����CpY9t����=�^��� � U�{��< ����ں�n���1˶�c�N]5��)��ގgK�w�3SI�M�T¨�4F�,,߳r��*�o#mgh��$�
����c����{��q!��I`F�r��I�Y3�R��I��<T Ġ���w!��fW9�5c�Ex #9Aq:��?���7��/]IB��c黁?�d>��;no�a�;&D���Ü9
=�<�X@��Q�&�#�sLm��[���UuC�.��;��A����//�7�N%�����@�;G��m��T����FZ�jRpw���Da�����㽔��Tv�`@�#5A��7��8���ք���ngZ7枪flw0� ��6O�rY1|//^�o=�Lyպ�O,W	���u?qy�q�:^��k*	��-㣎�2x0�e�Ko{�f���&��M��(<�8*������F��i5��Z�>�&"4H^IY-��9%���*���2ZP��dp/��N�P���S%a����SIdĥm
�O��y�����E�����t}�c6�*	"��j��R����[P�pS�l�g��]�>������b�h�e��A�M��m�Ch]% |�:iߪo�1�?�@��/���1F#0Kc���P4�p+_�9L�w~5��	�n'.�Ee�8�=w���ꌞi��T#����D�C' �H��M��Y��l�s��ص5�q"'5�T}\�
K��[.�8��(O���Hj���0{���il�?ߺ⋻��[ 컼�]��<;֗�iP����G���z�&�vf���+Dowi����s��A5�D��V�E,�����dT����	�d�HL��lLi.}�����nE����8����ڋN��{���W,U0K�ǩ�t�{�*Y�1���-D����^)�#j��N��S��㗶l �����XaCJ�y; ��	տ�ݎ�\Ȥ��@`w!�_��v$�������>�]��R\$+bkT�WFRT��2�Q���t�w�$_����w���x�����JGC��iǮ�צ��`e������p=������N5"̫��T�+�� ��c�5o2v�7I��rK�}��~�f��g���\�J@�C�ȷ'��6W����p���#��A��hU�F��`��|�Ϲ6۷�4�Of�� o|��C���}�I���b����9^���;�B���
"R�#lv^��#t�]8	�o�NK�LjLΪrzBr�܀�����P&R�]�0L�9C.��x�S��d��Pی�Vi�_aR�aC-:O�!�U��: �T�k�+�G
���J"#p�?��C�V6�'�dy9��Q���;��.{��+H�ou}����.��
�\���Pl]~�ȩ�煟uMH�j*>�V�f���o�S�P�dUҋ�������Y\$�Fd��"��{LT�M�6��i�i�7�n�����@���n��뗛�k���@>k�w7*�I���	�&���_�y�X�Y�TzDYSgX��?�����q�7�L|4t[S,7H)>��ڏ�)�?��ITI����*�w(h��SR�z�ru0'�*Df��FŃR��Y��(`�!�=�+�nYn ����B4���o*���:#v���@�� �3�^�	a��]KeM_dV��Qh$*�6Z��/�,�pM�v��z��Q%9�Vf����hN�-��ly�6舀�[�n���#m|`��ܲ����=w�m�<��s�n��)��TEX��Ew\Ѭ�XjqHrp)��u�UgՈ��ť�&
Ak"M=���%�_�r�8���z��ۖ|?��b>,^����J.1� �2�~�����Oz�����vXe�L�fD%���S,�B��<L���CxQ).�c�e�`
#+��ַ���|dLB����T��`�:�)�t�T�9������ar�$NF��3[o�+_W�IAy�PΡ��@����L�g������i��GP�6�vqw4wJ�^�j�x�Tk�zL�=���᳦��;������9͆�]�����p���D��	A#o�1�-�����(9ל�I�ʷ[��-�/����ONN6�'�����E�Fmc�k�M��f�]����h��7�SАZ��Bؔ�]�:�
(��+�[\=@>�经���Ķ&��� WXȀ��n^a�R���P���e���X��S���00����qu���#����L<���P:���`�H�.��IQ�7H�U�K�'.)���Q��`E�Q
�g�g��l7�%Y��H�����a��;�i�ͅS;nC���0̌����J�>�D ;����f�*������a�� w��h!��n��¶�^��h�d̀�|i���w��T���K��N�30{�z�N�"���\�qc�I�����!"�����q�d�����9΂kG\�j���2�Ҩ��T�31=�W�(.~���O�n�!��{���8"�,�(\��	F�3&�R�r=�i�g��z_����Y\�ch�]K�NQ+#^`����"����� ������'v]I\��e���|��4
�Ϡ%�@�<��^��_vǱa?m��3�C�+�$�w�)�i���E���� Xkݽ����Y���1�@��	��C�4UX4n�������Y�^p�J�7AR����d��������E±��\y�t��±08�c�c{��s'�R5B�}�R�h�-fG�q�&�tm�
�� 2�-�h^ĩ�C�w'
q:��?3)]O�8RO�^�����#�X���-���N1�g����^����Z��h8nyj�K��ӆ�*����x�{ ��1���T��1�����I|J a�EMort�[,�ɵbe�>+�ng��OS���`�Ì���f����mU>���$������/P:/+����-N��c�]K����*O��	�Q���N����7��X��<E�L�m�� W�J{k�~X�����I�^F�=I�����yOW���c�����_��?؞yr5n��&���ܑ��L�7��P5R'܃��]�"�>�,�RI[�>Ι^�B���	ݼ�"����0���FǇ�[�.���h�a�jd�U�
3�
IؽFUjUn�Q#ͽ�ofi��=,=NP,�o�����z�,Gk�]�X{���NTy�O��"b�&����?��C��ù�]:]Y;T��~��9gZ/6l����o�y�8�}�Z���z(�k ;j��s�T�������!�p�G����V����V�E~��G(���W��)Ҁ�aF��E�<�{R��21\��m�@k\���|��l�����o��0)�P��8�MA�'mH�f�h��t[�#ǵ��Z�a~��<_��Kiu�ެ�t׋�h_l�"[^U��"\�%��7�[��b���kjV���+��W)������W?���ӠP�WàQV�֪TPb����C-���u�nu���_�#�9�o�����n�읾,�ɳe�5ʞ��&½iљl����EJX�+�������<����~Ig��~Ԉ躰8lBz��P{65Щ�%��U����i*˘}��n�==
i����z �e��'�B�� �qX'p�+o��ºW&;�C2U<��χs�-��ֱ=��I'��Ty
zɖI5�&C���0���/zʗ|'�1і�tmEF�W�pn�J~Bd��@y�Q�>�a�qם�G7�<U��)V7)�hu��G g*�G��ߘ������}��'�<�dmrD<׉�tM?)�a�rp�^	?i�y8>�1(�R��%�o���n���T���Τ���|��vƖ��X�],ay�O�$l���N� �y�E�z'���gqaf�޳�~���Svp�)�s��{�8�c���h��2��7�x\Vv�Yޚd&��x�j���C�Y	{�o���)�����xNwQ�׿g�c���T�+�$�S�}�xMsA�':�uS�����@|RG[�.+0Ӆ�(>�3�7 �����/ź'T��'� �Ao�m��Q�A��:3��jWQ��ρ��[~��am��Ώ���z��]kĶ�P�?�-������m�;9�&�/�U��i��-{�%�g���ŷ��ٸ�@�ۘ��M
��@���J�F��* }q.�Q׊���+�����RV���V�%9�n��zA��%	���G���K�Qoa�_,e�X�Ŕ�-��;��YM �[d���"���C���a�FԽ!��&y�o1b@�njw�Y{Zs�z)��]o0D�}��rn�[ASv=��r.	��*���3V��jg��`��1��k���--D9	.פ��cS�vR�wʬ�K�hU�*|}��j�Gw��L�Q�1�5l��Q,7jdB�i �-{t�ⶱ�\��P8���7�+�Dw�p���y7�:���<U�<Z Cʺ���R�ﲂ~6��E�W:�<�IM�; ��Mx�λ��a��R�,�yfY���FS��1��8W��eC�M4T^4�2�G��:��}!"��Wmx��W�Pgw�OqC�0����&�#�:6���R���@��L>�HaJ����e���uC��%����	T���f�^৪oA��J̹<~L�U�u�U߬r�WUoTY��l�����<}e=��;��:�XU ��j~��dҁ��_��	,m}S�XJ�
qo���[	각t	���Tӱ6VS��e}�[�p��D���F�����&a.T�$,\ћ{J�a����W5F�7��pȀ��S
��ʬ���+��Ҧ6^��F���w�ˮ��
�$���Ta�â"]�j���s�A܁���03�U����t`l�ƐⷞL��J��Z�a�G/�1���j�p
��ܠ�Z:'�`�#H1���V�����Qw�����&۪���\��)��4<ǉ�hU}}�v��p�c�F;��<Nr�\�](�2�x��w�����ϻE���cva�K�G`�UűX�����b������#��-�O��nK7<�?�F���m^lmb=j���עV�Cg+��[N���7�����@�?W<}����х܉�X2l�횎-)��� �s?*�����(9�:��Q��9�����֨��0'rb�:��^O�$�`G�U��ĩ �����бtV��$(�ꡫZ�#Y/%�� ���*�ܸ��㙏}6�ݩ�a���qRKrfA-@���ƭj�(��'MI+$4�&s[m\�nuݭ]�n��=9�u��0|��p�b>(綄��9����վ����{)�zN�.ӿ^�|u�
r�9�m��s�sǕM+e��!��}�3���i�ag4~�6�B�����2Vw<�9 %\׵�_�񐴡t�=g�^���%��{�D�+�1���� �������@�izؓN�T$�8C!�B�4����x�ڼ�@)N����qB�ҚD����Q`��䙩�G�?	i�E��?������������µ�C�a�m�����d!����}[#�� ���8�_P�JؐGP�%-݄;e���#� �ɻgp�bj�a*.O��AĐ��C�0������Z����*x}�L��-���֮����Cd��%}���g����!�=1�۸���`/"韾	�TV���:�sT�p�S��Seu�[.¡�@�R�u����![�E��^<Ј.��d���y�����QO"u![(|PMw<.n� y��?I0.O��n��!�ZBi���E��9`���C�qt$@l�3U��{@�M�Db����.����	���wU�\{���OZ�0���p�K�V��Ю �l���ߦ_(p��[W��(4s4P�|�rdG�~`v��o��]������X碨ݝ�o2qK�d�{>�I�(��X��6�(���K����?��mǭ�8�M`�@V��O18�h�P�{��Y�?�MX�%t��K�eN�0ʥM����O�\=�5\����̵4�+�h,"��&A�RB d��ί�|��wv���]���p|�8�@r9ELW�8�z�c���]�]h��N�W
e���B�z���o�ɀ�9t$���FL�׶�v�����A��V���e�\ ^�麀 ��FS�\��BYn;�n#�F�y��Y��?h��l:Rߠ�'�&y���%O���Z�'������-���b�7��]��!�ZͰ=�����|�/�_S������B��)j�B�Q���jYx�^�ʬ��+f��7�wQʆ���I��$���ۚd��+�����Nu0\��kα��� Q���G1T�7�o�}<}߅;�O�j�5/�S�ܻYh,J��$L�	���JR<:�s����ߡ$ �U���B!����D� =&�;V�x�ϱ�'�ʧ7��T��یh�X�����ˌ��������	��D־QI5���|i;��7�'�.�}�ԎKJ�O��`��;��{���B����o�@�,��~`Q"e�<�DbR�U%���x^�����몹(4�Zz7������q���J��f˃MI�v����Pe�9��o$kFq��>�p�:{�S�i݌��ݣH����~WK�������6UVj�����_���L�\,S�|�A���	Z)���Y#KzUx,�)s���B����8��U-fS�M����ļH�IN��?j.ء'�_����dl�dP��\ԻEy)�A"`%�"�`��`y�I��(��ǈ�^ͺc�!
V�5Fj�e�#z�V����*����³��e%ʶ I-י,� �Ș���a��5�K9O�S߽%����{鯕#��$K�נ�\Kޗ9��ȍj���:�F8~��??�6@�6���.:]e�L���(a!.��>-1���=��M����q�F�W�ޜ�ڷ��n�,٣�O�C%�ء��>L��'�utY���0�@���|����Fο��ge�ҹ�#
Sw� މ���ntk�����.�a�GL��h��]՚J���uR'�C�0��+ea:��Rp: �sq%u��p�Ѕ�#/f�$""�;��Ofe�67!i�1
jg�>vǶi�o�w}碜u���Xr�`��6&����]�}DR�]�H'I���Z���oH��:���)1��oZ)���si�U��I)
g5�����vX�q]�h�ˏukބ�6v�	\�r�~&gt�X��|]i{k^ө��n�__JTu���qf�;i˻���g:�J�08:��7ܬڑ�*�K^"�ҢyX�Y���"hX���)͹n���P��m+�k��t���B�I����5�V���x����	�d�����V���x��S���硍[���BRo��b>��r��m��H��O9T)���&���֨zۜ�H��'�����ڼ8J��{!%����/ ��#�M�F����Kg\-�,���@~p�{��t�� �J�^I��2�d�,�-��|Sy�%��e͚�$�g�[�G��:�]|H�Zy�k�BS�H������wj��Eb�j��ӄ"�}�HU �![�;���W)?�4G"B��w}x{���ɵ��~�}�?��⋳o���7�{��^��������oB�	?�C%��U��r[29ہ�8��4�{d^�������v6�C�t�?5�Μ*�$fD'0%
( =�UQ�6��,e2�*��C�Jy3<[ "� `��n��:������x8�d�{��L��x]	��+Az@�2q�P��͡t�����ן%�#�MW9�������H�����K�I��uk��o�^�P��'������U�����O�-�|{�rdI,�W���$�~��jXa�ÜA �ݢ|?�^+�� ^uO@zQ�r(�4�j��)�h��&� A��#�:�n4���-3Hť2-��� Y����j�;:��T�鰸� _?D^k��_R����B���c�*��I��g'�5\*%��*!�
�E�� ]u�����R��%c6�Ji�'?YiȎ٨D0^�(G+mN	���z�:׮���� N׷`�����,�SW�C����n��� ��}	,:j���;;��o������E��o�HP��Z~��h��^�s�F�Ρ4����A N�^{��ժF~�ݹ�>{@9��7v�]o��Rb����9��I3=��m彧#l�0�τ�-�Ǎ,��M�fޔԱ�};ۏ��{�A+��;�z�m�j-Մ��ЛS(u��5�EG��Q��f�?�z�(Q�iM�b�z�Kn��A�ԟ-�����N�	n;}a�c�hR5�lÏi��ɔ?�@"n�5(���L���%���C9���e����W��S~�Nt:�k D]8dÏ��U�G"�_%����b�"M����۾
�{�6�r����Ζ�?ϧ�;fĞ���	�����NLv��!�y�M�l�A\I�Pr���c-M9�Rd'6�$\cl=ż>���c�A�:g��3��	���@�/�-o�3v�l��7�*w}��|�%��֢�RA�X��m�5
']S�/�`��q]�ӑ�\�I��}9IҲ���Z}n�����m��z{\'dT�k�>k�����:��q1�d���CŮ�w���Ce;����������qU�#���a�H���ic�!.����?,|� ��irB�����(�'NƉ�S�RڝBJ h��q�z�W{Á$�m��] �>�\����T2f�/@8���O�'dkB�o�f�`$��hݸ^���*(-��+�M3�m�ͣ%	w�U�O&*[/M�]����T���פ;<T��e_	��u��~Fd���Oz�ϟ�W���������֣zV�O��?4B�wK�h�Ν���4(sӈB�~�9�]�	h�1�"��+(���vA�We䉇|��)�a�3w���� 6�z�����_�Ji�9|�yn7�kt݃+��-���̍rV�ULf0�r��婛������F���ث�]x��h/7��f�g��a���v��E��`l���3�3EN<���Cm'�byі �a� Q��J��WfA����c���q��%�����)��K1txk�J��Ge�z���彷@>�Ԯ,}�&r���R�]�/`|%}�d~�UK�L7��Bu����}��XB.)H���o�>�5��}��/}��F�`xR~V��,|��Y�����e<� ��&�d�l���d���Y}��`7e����3�##.���ES7�}*I�	��vqȝ����k�����@5�'LTAe���ڗ�ϼ��M>�5��C�+sp�vD+hK�L(
UJ-Ȱ�K^�Uuھ �%2ٲ`�n[����<�G~kr$���\�s���)�~1��I�4$C�A)X:n9��º �X�]m/JF��1��g���Όg�"L���;=R���'t4�?��@�h�t1x���O��_�-p����)����R�;^�

���}�H����$�R_�F�fa,���	~w�P�[��]4gE��EF0�M�Yn���R�pi4�>�d���m�0����k��������%��D�_y\*����\{[@Њ\o���F2��-��
�-ZC�?��%&�g�ԑ��M�C��q�!�p���U�>�e`��0�/ʞk�L\ ?���v+��?���$�9��ِ�^2�g�����?`/u� *����8\�5�%��������<��c(�����n���m��:�w�OrCi80��eq���-�ăX�Ý?�����e�#�g�P��E��������EO?��8_&���90+cǧq�}��)���Q/�Ƌ�C��?�A��J����1��8ҳ%�������uƛ���Ud���f��*Ft�����.<�A����E�j�g�1:��z���hMѦ[�o���8)U�x0h�Ucy���e�zfr�<����k:n0�T�X]�E�sqy:j�
��Z������&�(�����'�&�XT��������`\h,sd+��!�(qZY鹿��\��s�Ĉح�1���1Ù�Ě~�n.�gt�a:-���E��L��â�jn���`]\u����0~������V"��M5*�J�8̐��s�DN��hb�U���r�@ט��O��Zڀ�8a�� i���	ܮ`/'�j�]��Ƙզ�6P,!���hfۊ��[H)�Mʢ�yή�>K���R vF\�����4(gQG�9}�x�9����SD1qT�Apu�gd��@���K�%a�I�ƕd��b{�;\��yr��knWXq ��։�Č�
n��Z��.B���,p����� �S�)���"t��Ɵ(�����[�c� �}�!%�}�;�\�ީ�軰7��#��VdU���*�6m�x�}�3=��)�rn-G��q���]�"��$pNA梩�'ۗʜ?,�,��<�a�#dl虿�H��I[�wLk�R*�������n���BW����>��{����X��x�H=%EJ���G��օ!���w��Gf[b�h����ݦ\��D,͡����	2}k?	��9����L��rGɤO�&f���H��"Z۷�_��n3���U��@�����P�>0dB�蕎E�����4�x[O<�|�f�62�Oٖ`�f�31ǝ�兠;����Z�{�RR�% �f��K�e�ud?��#�$[������H��z�}m	�jAeq��~�"�pF�sa	X�UDО/�W��H���
y�D)X�u`<�����*l���kj!7\�R[.��6wK�����7%��}��o5�5����WU8����^�����e�4+���I�k73�?-���IA�P%��Z65���eZ^����48E0��O�$aZ�	,)/ �@���	3���C�,�.l�z�F�Bk'})�`7/��Ŭ�-�o�m[���������Wjc�9]}��E/�"U����鍲������C$�(/jU��?tZS%.�"�9O'8�߲F�0�e6q��YP���)�B�7�� ���_�_{�<����7��?~�ѨX��V����6�Y��c8_�����b\K��u�
��S\e�,��d�ɥ���;����݆J,��
��@n&��h��j0�t��;�>�����e�a�ns
�DV�Tm�(�m9`�H�m��k���`3gm�-6�F�����EK��|���l�!�1�����eo�`oS�#��I��1'-��5a9��i��u5�9�=N$�Ê��sϮ��bә(�JF;�B��M�^l�/#��''���U(湳	�GS"����߲,�gOݩ�H��
��bWgU/R3T��i(#�M���?a���=U�L*�H��h���uX�]�$�C����J�O��_��*��j	`'h�l�1�Lx�>��iIGu�Ȼ�{��l�R�>��!L̈́�|�1g�x�V�B��F��iHm���v�kdT����ʹ��0��u�+Y<�Y��X��qjK3��+^�V�S0U�z)Z�����7��s?��^�"�Z6&�z��w:�\�+���YJ��^ҀM�,6%�:p����ʿ�Ά_퐏<�	���� 0?���,05��B�ğH��7OJ���Y��T��T���I���ς�C�*J�o�ye0�i~���s�6��~�����b7R1"�&VɶKt5|�EH� �b�����)�t*O��]���+�0~J`�i��`j�{��Ё?��xxЦ['�P;>�?�M�pS���|��"�CI�����S}�clᬃYr1,6A=�i��e�x�f	���_~0�qe�lm?E���c-`#gnbﺦ'H���Ī��0�Pm%Ѿ�����Hա�4�/Lk��1�1�u��Z�V�[�e���V���S�H��-����%X�Ċ�W�cMc���%�-���V��B}���@��ʤ�^Q�n�
�CH/$��N��ؒ�z���(�
<�x��1ع�t�`��@sb�{���3�JN�5���X^_Du�}bdu�����E�B�O}.ǲ!�&N��vS�����ׂD�=iF��;��s؋8�3�90�4cRq@��v��i*2�Z_��4A	E��?�k��p"W`8ϓ��z�b�n�dHa��?���_��y�sf*H�]M��T�J��Z�G��Tkn�𦛩�5q�O}W��&X�'����*%cc��! �p=�n��7��H�7m�1�-g�ږ��pַ{i�J��M��Vti"����eh�D"���_�:l��������<�.��e�Yq�D�?Gu���W�G!�z_�קK����7pMX2ތ8�(��̨�2^�9@�4��Cȡ�5�I~���(���L�uŲ콴���h�ŶN/s�e���h'�W��g�wpF���$4EĚ�$q���2���FZrf?��b�<��&����$�Je�Z3���D><��Y�4r��D!�/4wK�Vt�ֆ2��"��d��|;�{��K��*�Ck�El%	���Y%!��>���u�:����R�azɡ�d��~ܸR8�����le
@�ץT�>��K;ms:�uf�{\��h`h �N��7���>K|����P�
�nriwW��SyB�A�i�fU�ŭ<��6"A\��5�d'��oE&�{=B�;�|=l)b泮�A������E����Њ(kNl�y&�}'b/��%6,��l���(�=�����_�����Շ�9�������+&���/h��cӒ�(A�I�����W�r��׳��O@��8}�)�Ť�������i�n7Ez��3p�͘4�ݻ��%����=}�n��~F�hW��%A�����2::G��(�_�{X_�����,������+� ��>��7?9���F�4�R�䨝�$.��P�ϣ�+<��qYr���~
!���<���<��[o2N�۹������P� ��N�y�ph@�T��pÀ��n9+��L��<62��f�-'4:s���i�����$��'n�+㣸0�R<�x�@5��Ҫ:Zf�V)�Of	ί�����V ; .��*�&�Se�y!6�;~�`��ی��O�h���.p
�͡WrM�"�j�V{�����&d�+��A���W�_���zd�g5�x�z �.���Qu��z;V9<��+ ���3�{;9�	֧�2r�ic2������$�\2!�1���G Kx���`�����D骶a&p��Ԟ4�0����d������b�O���