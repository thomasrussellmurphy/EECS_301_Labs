��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\���V�fnvx��ÍG_;�ȅe�~�>���9�>��Y;�0G���O��������Z���G��A7��e׺o�o�ծ� tR�I�3\M�XŊf����mq!R��i+�e�ڶ�H��t?%y�&}�(X�D4�bc�7*)��M�2�SNM%f��N?���؀�?O�H�o�5�|P�!]{a��@!?jM�x�稍=	�x�&:�_F�r�l$2��c�bXLšR�0�h �K
K�4�pͦUN 1JĐ�d�0�R�������=�b�`���Cx��`�E��/�gӛ�5l��Tr�r�܊n-yƥN�'f���q
\#�pm�0I"�<��Q���g����Gؤ3ׂ�aK�d�T�7��J��9F��;;�(�,l�O�-]��FsIw��~���R�|���uj����y��峵,��-�&��ca�->���r5QJ:���+ ��F��|��Y�V����s�6b�k	����6)�̶�����[��X�^t�z�%Z�f��&@Si4���4�n��YB"mq-���Q�W��sw��?"M��q����իf�`�8m=w�	yi�:7���^�&��u��,*  �.���!��$���L�l�m���'� �f�$������(g��7��9⤮��~/ 1��c�P6u��� �$��{�-~�Ee�aV�C���gT��������L�9�ֽُc/mƊ]+ї��~) ���yU�PC�U�����&�¹��^��8Z�݂���V�w�.���:�ۭ5PG�y�'���uXH&�O�Mе*y��uG+)7V�o��^(��o[y2qs�Cb���?#CX8��
��W�a�/c�cF�y�GZ�JwC�mb���!9q���m�J�?rj�mE1J�ce���]u�\�4�<�+c)5�p�%q��[ ���Oªf�bDg�.˯�6�F瓱q�Q^��R�W��A"�r�0���_��SFrHTe3UeL�L6���ƘSD����lVt�s�^���7���|���"�]g��z�n�8e:�.����k��M݁##0?L�*(/���\s6��&*�)ED��}�����iך�+R�$N�k5v�!]Pt�(`���Y6-����ح�<C(�
�)���8�R�Z� �ލ{�`S)�巾��sz����M��$J��N'���T����N� �~`�g��W��@����D{���gp냬3�����& �7�G9"hr��Φ���Qf���6�L�]5�Kh����w�L^�t�ۻ���M_@l%m^���}}����&��S9�-�p��;��-GKla����c��MB*����O4w�1��	9ߣĒ��z]T�<*d\��ҴkOB'֍����j��b3��L�JQcKh�̈́��9���Qfh�)!����I�%OS�kz����C��Q��t~6����?�0gY� ���
�/R�4���M�T�MNߡŬ�q���Xr�z���k�X��Wd�����7�dN;{��|�U�s0?�Wm�'��hq�rD	p�}Ҿ�_�ݞ���?�C�B��'"�Ͽh���ˉOf���~ ���á�S�y�xy�<h�e�%�/ёng�r�w��H��M#�֣�$��~6kix۽��N�|ȁL���������]�n�Dn�+�g�ɪ���s�lH�2�K	����eUmKr�բD�^���mH jp��nF+Ñ�T�Xwi���>�+g�?�w��Hp9�j{R#l�ge�Ix]&��>j7��h�E�{�1E�DI'?�|n6ޠghv�#�#�Yb�,$p|����F���0�\�l��U�ʔ&<&���ϯ�Pd�]"�j3��G����Ԡ��9)�P�R���Өk��]�����Ƈ�ҟ80����mf ��m��$!��dY*?؇L&1m�O�t숬,Cr���6Z��0N,e��^���D�K��*����,����	-���/[��W���{��o9SOF�P-��C���f�w�8�,,�����_�fU�[�nM^}��#u����|����de��X�o0�&�h��L�	Iˑ�{�qx���'mX��u�,�r`�;�W5�Q�^jԥ;;�� q��w�+�"�.2���4�ʁ��򡈼3�M��g~��u�^�U��}@��ↄ��V�]�<���^e�;ᾎ��i��vx�};�Bk��0	�Q���p���dKm̜ w$TDe�2�~�*̀'�u��?����>u���c� ��!��R�Z���x�ʚ��4>�X��XX�5HS�"�S��Qt�1�����L��μ�#޵��V3�քۆt�w�Y��#���[��A�R�G3���Ht��)����:9�����$'��U;E�O�H�A�s�w�����p;|���"Ə_��� <�_h#=��dQ�����ya��c;=�PԌ�1��=�QqWS'j�?�G���@��]�wx_#��;���%+�kK�t:�R,�h���7����|�����z8yh*�q�����O�Qꅆ�(���!z���h��G�UF�p*(GL�KpJ�@JT	�����:�L��F*g���^`���r�\�+�IPRe>L+t��ǎ���b;�	G�^����,�&��?�ζ?/Ba�~CUڠ��xo�������0��"o�ޒF�f��tw���]�r��T���/�[
@oIk�"~����X҄�]z�<���~B�>q�gH��w$�Fw	�R��fh?~�ނ��w���?�)P��>�'a�jD}P�B�m�+ȇ�f�}?��{(����a�J&�u7听d�V4�s������N��b�2",�:��@�_j�xڠ��j��dԖ�(�*ř
���WcH���y��v̓��G���v8#L�'�/����P� k�զ֯n��9п@GO����*�|q�p�����x�����K�Jn�VT��9�jl�xl�A���a �I�_���|�z��63 ��vC DDK�� �h"q����Hb@�����vI�@0�8w3�r�"�f��5���E+��,�@����k�����]�J��CF����q��C7�����G_�	��[�|��;��p1��)xs�*$��fZ�-p4�~��3���<����A:��1��{�1Nw��Ӣ�Q��<v9��2; 5����.׃f"�K,�XV��a��c�đԕ�b��O���L"���K��\�S��W��'_}�k���d�+��y%�P�2�@��E�p��� 62��ʮV�9��ӳ�{#���MGQbq܌S~UU|6���\�@����3?�y�w	�eh���57.6K��V��Ψ��%�q�BQǄ���*���{I��.��t����(�m��1k��B���c'�f?�4��k�],A�:k�X �L��l[*�B ~��x��qyQ8�[��qX�iH9X�����/7Z���G:+���K�����/��EK1rBY��,�8/%r�q�|��u.��{�CD�:�m_�*SA���}|g��M#m�3D�]5����6��=��Y��S;��/�<$�LՅv�����y�!h�G|G�3s���о��D���0���OV�Lj/�糆=��|V��8!Q��v��w��
��-B=U{*X��ο�0CЫ�m�,E�H��F4�� �{#��K����ԙ�E<Bݯ��+x0d(t�e���%��� ���B^M�uF�Yl�#�"	v�o[ٗ*�
��־]��d�t{2�����\#�)uD5}�*�_Z��¨ʆ���Xv��u��#��9�6�pR�,�g����Ï#�7�v�c�1E��)���T��ﾉe��)F��&�����0R��<����\BZ���Ĺ���!,}��m�]4��zk��W��O�uF0�\���*��A��-������.1�6�$����qPz�E)��Xe��.�FƮ"���[|�j'D��sL&3D&�i�I�����#�0wP,��߉�2����x��b��0)���zU��=��]E�f`ebG	��r�-��o���P�i���&P��;�zT�i�Ep!#��ZM���y\�*A�l.`�����#K]���1�q��5��&2��"�StN?�> O��֍b���I��etssW4Ocs�6��\~�/�)y�ɨ��zl
#g6Fq�\��Ui��0oi���jPGۀ��6DE�J�8r_�E<U	(m6xΕ���f�@˼�\�d�T�Z�OW����٦�)���i�?P���o1�1��[*�R]A���2����3]���3�0�j�
3���oKօ�7 �7���|�޼]��=Nt���Ȇ_ /`NN��.���MF�N�h��|��*0`SRA����m|�w�߼P?�P3��r�('��Bqp��`F4<BFw��*N��L��v~�:ADh��ݝ���i�;��9�O"�������ZV�p�-S#t���p�M-�X<p/y�JEY���s�P��h�>1��O�w�cf���$���s,)�>q�C�J���� �G��������ڝ�)��	7��R��	4Vf��sbt�VE���6..]J?��	~Z���	6�7��5��Y������(J�u�{��!1�k!��.};�V�)C���J��&�����ޙ���v�w�;� �jIR����n�L��9ֵ`�3��~W�f�Œ��J,�U���L���aHJ�e�R�?'�� ����� n�6X ���Qw�����!�NW�_q��T��b0�1��i���n�qŇ7I�W�v��V5���/eq~1��\�\��2�����> �4�(!���?��*Zf�ٚ��,P������08���p��L��˯���3����we$�����z�LR{�`֐O�u@�=S�N������{2�S�y.dz�C�����3�l��������^��Lp�U,.��Ϗ���W]�^�ȿ8�Z�J֊E��-r"S��K�A�� $�FHz��Ԋv���U?�W ����.y�*��8��$�qɘ$:���3��0a���E�Qh�D�g�a�}<�IY��&�m0��露���F�h����s8>���CJ5+@|{����=(EV����_�Yc�`b�R
a���\��~K�6ъKC5&`��LU�
�}NL�����NwV�ձKb�gT��1:h@�8ʓ����u��y���G?}R��}��ӣ�i"�4� G0��=�e�+Qq����"5
u�}f%l#��J�:�y4��UJ�ony����G����ϋ����:�6�.���a(:��Z�� �@6@���X
EނJ�5&w�5
���sAq����M	R�p�*$�ĩN�CwuV��p��F����@�F�$#��B;$T�3=��B�1�50���u�M��9�
�N��TAAڊ�AX��HBiIᛌ�1�F�	�l�f�>�&;2��2fߤ?��T�:qȕ �l�H�rw8n��#�lS<�#(k�H-ڡ\��ڞ��&� �i������f���~��@�
n_z��z9Oa�|� �e.)��K���(N5�mA�˜i�/���s���7Q2�>%�Z��cۼ����vUE�d ��?�H>��~�L6/ޕ�/̌8����͝��2t*"�F�*��G*κ�Qf_��~�ʂpJ̐�h[��k�\�U�6�{8˷����/>DwB�C��>�>��1��:p7B�JA�ߖ�i�Y�'�M��N�ޕ�l���A���F�|:ξ�bJ�x4]0[��2&�
U����K�a�1�$��*Hvu,���ٰe�BZ�.@]�HvO�m&?8���"����#O���&�,V��p+'��Ug݅��k���O����'Xn�葧��??&�jpc�h�,^��P*\�"_
e�Y�џt��rԛ����/Ը���;�5��"IO��>�0����U?��������*Ȥ�8v��E�q7�Ka[�*=��E�3�7y�}���h��pqދ�^�%c��L�]�9[V�&Q��2�d����okhԈ%�"��6o.��-y�ҩ���~��Y���o%���3�i!@0�����nY�G���0�����1a(~��H6�[�._y�إ�8szY,F'k^j�(X!��L��M�<��j����D~{��6e��<����է��F��*I会T�!.�5�84QlE���E��B<y��;��y�4���:�,�J���#�F`2p�3޻s���DS>m�k{R˛"�üJ�/�������կ>H�K�����4�;�g�X��ݬx�{����8_P�_
񻦲��v����)���Y���I���'�R�=���Ȉ�ͥ�vm�%��b·�S�G�h�����b�$N8��[O�T+���DB䊖~+�ɲ_v���_z%�a8�	/�j�-���ք�`�N�B7���;wP��~mѸ���s̄̍�w�j��C�W�٢7�^�]5�'q��t[�O��1Sa���x-�#��/i�֬��>S���3��an��ߧB���X�q d	n�~��|W�N��M�&��_���ÖLRD��JZ�4��`N@�%�ȹl�{��$g;��y�M�R�<�f�j�nݓ�� ��e����#)�@�*+�x�Xs��q��_�"���3D�_k^T=�ǉ�>�YB�g����X�'_�/��c�i#.Q� ˏ�ůb��4/a��һ�e�a�/��4�8����;��n"x�`�)�GQƅ���3s�g�