��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\���V�fnvx��ÍG_;�ȅe�~�>���9�>��Y;�0G+��{��d�=e� +�.�~��)!~&r�J�d���K\�{[=�I�֙��;آ�[��HZQ�-�i^���	��7n3F�:�Wu�Μ�/W[��}A��LO���v3*B�G�
�ھr��U�y�_�X3�<�ĳbu�O&�"�F��������ﳳ�N>��pD��Tr�So\c��o��P���sJ��٥A��eȶ��G��K`B�Z���-8r���e��Y�x3��O��c��k��C�����0�����E��'LJ��`��N�c{"kl���ly�*h2E!���Q�a=�,�o;k����XG�0
{0��< "4�O~܀nvI�7($c�
��,tb��]
�]��0*��v����kT�:F�O�]w�z�fZӒT��s�-�Ӝ�)�1�P�������i5�2�z�`jzݵ���2�z��tLD�2Q���?��ګ��&0��;�\X��b��V�H�*w!���qs1.ӑ_�d��Y�#<�Q>���w��F�}�ـ����ё��ZW��+�M �����,D�ע��%��7�tw}�RMG.އ�4� �{w%���
GI/��,��(I8�k��v&O�~�];���'J�,1EC�����9��*j�#�K���Î�N�d^��C�����i��z�g?e���R�i��߻�C���qU!�"޹ي��<�����V�� ����Sp��e\lfmϴ�e/\^�.�B�`$�-�0ʶt���S^�-�o�.�r�'Nhwc��(�6A\��]�s� ������T#ŠPߔ�`�8��4Ch�_��j	[:�a4�R���%*��h�T;D*f�g�\���cR�a-�8E\~.�kY��_��f���߽�K���|����I,WV�|�s��@D%�� 
��y���
=������6��?f��I|[�5��C�D�b��}�)�~������c����k�z��f��t�� %］�s�N���;>���E>D:|㩫A]�j�;�۲�άt7Q� �v{vN���f���L�ӅGAUK�A����y�\K�RN��L�.�!��/�{rM��;si�S�X2��,�T� ����̌�X/���j��) 	���h����nR%S ���nD�H�7F�=�{�	�k
@�.椠�+����u�{AN5&����
��1κh��y���FO\�g��<t��U��s>�E�D�0]�67�-)�h�c5_�n�n�h؊�A�3�>����	$��U��6@��»�6��[;@>(���I�e�G�j�O~N��T�