��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\���V�fnvx��ÍG_;�ȅe�~�>���9�>��Y;�0GZ�Z��H���>��< ��V�ũ��W[g�3K�E흳Z�6o{z�Y(*�� ӏX>�4�UM�j0&�]O��ϦfPt1�\��_���Ҋ�]���p��m�	H�f%�Χ�5t�T��u���m�9F��=.�D��D�K3���^�P)u4]�u�5��?�l�FTj�x�Y�����+K��i�����Q��KQ��_�)���|�qN;�SXg�J��kst�7R\%�tH�g=j�i��%G	��K�J���+�[������@[$S��	HF�����:�=z�}�Ceͣ�?�}�'�LPXG��pV��k�$�
�5N�B���n���'Zf�	m:|��L�(�

h����p��rGI�R�����c�Ů��_�sL�sQ#�抡hiUn�"�	�A�6vfW�| e�d�f�Zg��<}��!�6W�}qIB`Die �q�'����rʮ�O��J��-�J��#Re�ra�40v�/���F�=YM�q]��Lp"��=[)#9{��4B��zf�^��}�~�F
�	��{|^�/��(�����4Qy���=�繛��Y�?Xh��hD���,A ե��ժ��H_d:�/�4H������/�4Sj�����]}9�~<B8�b����(͙k��|�t�{�� J��fZ������P��Z�H�f����?��k�������uX��>TzG�MI�9�8���F�J�Z!�,¹�0��k&��;YU�<���|l�d����ɄL�$��ۂ~�2�Ի�_��f�8�����H���5O�i6):��LS
Ʀ��!�Ih�M��9�ɳ+�!R�l`��G��P����R"C���{64��W��jX���5G8:����,
���s]�!9"P؊��������X� 4�\��|��=)�i�kx��E!��6N��G,��Gh���E�F�y��CȢ컇����;M�N^u�yW�(�!v��8��-��ej�3O�W���e������d�n���V�+�e�|�����byE��]���)�6!0��<�ri��~ka�u�C��xɱ(/pc����H��
o֠�\I�Rn�?<�����1�[RwL���� �w,��ରl;� }:�l��!��|�
��tI��́ߺ)���9���=� 71�� J�4Y�����L󎒁h!.ru��!/3����$��&5�����´����7j�܋Ӭ�
w��N
�)�ɰ4��Q����e�J)V����uN��ݺgԈ^0:�aF��	�a��>�5��bIV�P��=�Ҙ��cص!EM;q���w��4s�}0���ܾ��䩻bi,i�7oZ������:6��I�,/BR������A��%�̛vj�_��a�[�=Cl��r��+P�+X�
(�>|d)z1V]�u��agC[ф#��Ǩ�H�[T��$��u��x6l��ŵ�[M;o`K{��Gq�_L��|mk(��_^���^j; �=��;�k`�QZ����־�f ��&
jV�P$%)�#��(U7? ���2���,�\�&1]�M�)C�U\g��N���m4�Kž�&Đ�' ��YA�c�yP��9Q�,�=i����T�n��7޵O;�ә[���rX�w�`����D�x|<�ݪ���s�/�r_o:�dC���'����Y��KR{�L� ���Xry$��\�:?9M���WPʨb�2�Zt��j�h1��Ø�U�4;KTk{'+���.F�
��{�H��z�ڼ��﷓�Ӣ0j(�%׶�F3��(�3D�-t�Q9W�(��[]�&����i��,�<!�u=��vs�}���$F�X⹣t����?��+1�f���H�,}o�ς�+!,�z��<f&X$w[ޚ�>A�̙E�~��ߟ�[���19�L�S>������=�
}ـ)�>�ma"|0��Pv4Z��z��!=��[��)�`r8��Xy����ga ����}���AIt}X?�����ǯ���[�I��\߀����z|������V+�\t�0�M�U�j5�q	 �:���"-ϑ��n���V�s`���h6�tb�r-�N*M��w�/��X_
2�Q��k#��L������C&@�W'������οa3�[[��9��&R��tE�
L(����M43�gC����b���~p��*)3ܾu��۞�ʬ�XJJP���|!�;
�IY� ?:��v�����S�g�Y��j��� ANi��������b`������4��ߝ�'$����9��{�s�L�̩Bcu�m�,�i���#]،�&Me�Fey�^jL�{2�B�:!˔- V�7A�����i�j�tc�0�>-��2l�%�����G�}<���'�x�0�()Q���Ѽ������h1@��=�|r�"�O�e3��k�8=8��TêI8#���K�b̈́� �:�*H��
�^�qO���P����ov��'ø٩d�y�mۆ�%�9�B���Ji�~�&�X;��`j ��i2�B��X�QJ�l*��fg�<�hJ� ��-�G��3�	7���s=*p�~g�\�f6��ϟ�����\
�2�0��v#�Zd�A�H.��A�T���՛iKy
���	Ez 2���~��#Xn[7���?tTt�7���₮cƙ����=�.��-spzH(t9�wPHi��S�pn��u}�b���q��؜���8d}�.#�v�Bcvךb��۹�C���4P��?��7
������7B#i��d�_�/��f�cgiD+���0�=��]Х�ߖtvm��D��Jp���UR�1�ܷ�p����-YiDc����C�ɕ�&����R�_��C���zAK�O�d��]���ZͿ*��7M^B~�І��p��4�� �y7�(O��?Õ�iM7ں4ݾ����,��LS/=r���<��x�o8GD�g|ho�4 ��ȑ��)�����Ό��Y>���OKy	O{T���O*5��`���V�?��rp���6����Ǧ'�+7�ֈ�g4���;�b��*Ô;l���*��ㄼs�C[�U��ǔd
�H�����oG�����'r�\�6ؚ�[�'��#@����w>����y��L���w��0�������A��ӛ����ign��x}���w�b���Z¥� Oo����)��þB�a\��m�Z;oq@���'�����ejI_���Tzokp9N��w�<���D������\��rt0�f*�p��Q.(���+��?�pߏ0��}���wB}u;-���<�{��"ثr/..}_�+zǥ�
��ӥ�D{����L�hj��rո�xyM�!(��8�����t�޵��
�eGL6O���II�K�me HK���OewZ �&9�be?�[����"���#,�:�����Qlɥ6�P��K�0�9H����q��b�%;�8#w��.<,����t̽�RJ�������B<��{A�i��
�� 3�<����ͻ���pU��!*�c|w������B�$���lz-��=��	δ���;���gQ����(�,RPyS-�(�O_�L������O����8�_�^9����i,"�4�m3eW���MX�jjUP�89jƒ��� R������#�8�� �o��'۟/��q�?C#:���fȚT�+1FL_�S@&-}{Q�H�QO���:��cSv0��[�q���gY;�;��6x3!Eb��f�y'sr伥�4=o9��a[7Z^/ۂܶS=sx1Ʋ��p@�搤��M޸������ ���D�cW�g
�����ml��w3�{$4�J'$�ù�i5/���i	a��\��o�7�3�V��tP��,�`	����
��\��S"���=���D�ĦmW5X�x#�	����Z��	��#Vl��Y+W�&"bx���i��%�	1���I�ߕ�ӡ�.���]�O{f��w��I�_����*
`���9�ΐ�cwR��c5P�~49^ �<���wS�贏����U�s�ث�2�}i-Zq�­�j���7m���yd=qo�o(́�H�gT,a���AEW!4�j=��ĕ���>
���h	,*@�_j�t!a�ޜ0�4�ݢ*�bи�C��7����iN.����=�T�|�G�xvOPn/ڌ�wW�;�j��Q�Z�冷�� "��ϭ�5@bp�$�&�]c��1�ώ��T�,I��1�[ �*�X�<�?�?�����5��a�*��\T)_��(<��H�b
�%��Ϗ뫧��ȇ� �`�Ptkt6��.��FOo�ZJ>�pu5]xe
��(���,~����a&<�+c-G*������rjr�uk?�G�*4�}w��<e^�ѩ#Ly��K�� �2۝�*��GX��1W��f�)�1�,�ɑ��C�%{����IO���(o�Z'�ꐏ��]�
Ў���v_�U�g.�V�!v��|!����w���R��P�뵤�+ba���ޡd2�Z����6�n�G��A��| �.DpY���(�MG���F�T�Φ�l=�0�;��ǼT4���q"���F�/�u�:&�(a^��T)HY��A�G�}{�42�Y.f�غ�w�uŲ�/�����R��]��`ÿ�uȖW�q�<O����ݪOf�PT�9�o�JHk�����c���H�V,ΦIİ�y�Ǉ'��.+����()"o�t��[���`.�˝���T\>��kƜ@�(�+K�eNB���ؗ�f'��OэX@���QRH,����v���=k�PYY�#G�������}i��1�da�-LT��Ԗ;g�2u���髸�(q�>=$��1
�n��M,��q��άL�!�<�� �ϿHq �q��xe�"n�en������}�2�Ӏi��iOw]\�b�3�QX��Mj�;vD�c������6^�HL�Y��W�H�xOӇ���-f��,l%>0��@D7�`�~4+-�)&p����eDO�k��AX{�ѫw��x�_����j���E##y�U����fM1�x�5���@�1)	��6R1���|��#��}��J-xG��ﺈ�s�M{,\ڰS����I�L�
*�|r)�ƞ���Y���+X�X�B��xb��]��ϥ���WK� M���x�pWk��=֝�޶y퉝���M���ś��P�<;�EI��	74���v����|�����u�IM�E؂��1�O��6#�^�p�S���F`�����%v�~��e���������-#�i�"�|P[��%3]��_PI� ��!�`r��/F�w7�"ZD	�[/a>t�0������GpX_/�_�3����,���������ǡ>#s��6��@�~0��e>��7u`�e[�}�)�u���� �>t݋���I��!�z�&4�M�4,����}��~#�خgbx�֜��#0��t㩱��j*+�I<](�p��<��g��`�xE�Ч�I꩗9��ce����b!������;ˡ<bxp��
T	wae���=^@��tJ���=(�EA[ڠ�Պ�[z��M�K7+���r�����N�MZ�I��-��<X��ҁ�V�����Q5�R�t�q���B	Կ�� 1I�}��B�`%o7O�}�ef�ū��x��#�G�2��U	��l�ɼ)Y�gf@Q�xY�nr��$\�T��}O�	�ৄv�/�2��\pdgC����i4q��Y��A�}�������:_`����as�BsK�V����˶t���׷���Ы NºM{yK���7\�-M�Fx�P�(Zj��V���y�(�P�j̅%��0�^F��>�<9�J��2�&�T���(��0��C���A���,~�����Iҭ�lk��