��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|ۧ[�����Jˬ�\Ũ�k�c�5�xLt�Z9���c�U�G� �-�9kÉ��!`f!��P��,�S��8�
�zw~%Or�w�:(��FK<]Ğ|Q���zp)�bH��y~��h��;���5�-*D+��[�݉w�]�P:.��i�j�!���έ:��i���	��P�P�}zR���}����ju�u��eK�C�4(�A[�aov�Av¨ۉb���?���+�����O�CrVQJc�1��c�Im.Ze��ƀV��w�Gg���)`�'���z�NțF���Է���8,ָ�f����B��f����]RȅF����fX��k���Ÿ!��u�/���ڬ1]@���vN�m�N��h��>a��vy��]5�����K�l �ƒ݀�,�u��U���6�r����x�����������e���kEj�,��u��B�>�'iQ�������\����}��+#_Ae�hR�$|?�}��ٓ��cd'�v�ߖ����c܏��JLkIĆ����$	h��gI�]�4���F[MJJ��=�Du���D�'��C�Sx��Mn<�N��,���
�.��l&�Y:Or��ٜ}�?�ieY(��Y��b�r������	�}]��0��/b���ב��+�>=�L��!�I��8�>����jμ�����+gmO� L+����{W��f���R��M�K˔g�&G���}��]F��@{l �1�M���W����j1 ���Z����AI`�[Q2�8S^�c�k�Q�H$*���J�$�f�j�Z�n�͠ԙM�
�����*&M��ۨYE�z�����4� �?C���+��O#���ƪi�s
��M�S��幀��\f�3)��������i�B��n���[�tP���6����q�]��V�M���� B
��ܕ�Jp~�%.�aʄ�%�uF�'f��s�ĩ�#1�ǳ���6��Ɔ�"�%���h�
��a��I:n- ]�C'A�����ʆHy&�v�Ӿ��3&ݡZ�J8�3,uo�T놌:��g:5���o܃h_���7a͊:5�1�SL����OB�r�C̽�p�����e���H�j�)@��hI5���7XX������)�3��U�_v6�*3�żvZ�s�40)i.m��cF3�e���8�X�/,m���o"D�#�T%L%RA~��h0t
^�do�S����z�u��p��^���Y��b���:\�`��<�ч�ӵ�d�`�V��R>DPz�R	�o1���+L���/[��=�t�aQ�c)��,J3� �H�d7�y�(�i�ֽ���w���N^�o۷еkr�<�=�R的��Zr�͊8��X��eBׂ�wf���ԂR��?�X����f�u��B<�%�R���DZ��?���~2�Ej�5�'���C�M�YJH�����l�� ��GG��B��3
UL�y�����ҥ��>Ges9�[��sK��`�����"}땷��c�&U�)��$m��o�� �f��.$@.�Oo��,&� ,���%̏eb� �8~������M��ovʦ��-��Ӛ���h���"k_�N��<��$X����"����Z�d�W8�>;%l(r�:/kѮ��
���c�0���K$=���?��!�L����?T֋~��(V
�b	�~MD���E��h��	!�Ah�g�ľ��QK�槽I�����|��j �=¸!�?�=6$��8�h��aA/�=p\z��0�^� �%?rtI���!j��ÎxU`�%L��[��$GeAJ;+��/1������p�%��rv/P���4�+X6�Xh�̵4j��QWr�{��m�X�S�#^�!�V��M�7,�57Ȑ�'aD��Vio�9?Cɲ�v�cp���1�j��B�h���:O�q+6�W�a�4���jᨗ<pF�Y)cuNeF���P��ڏB�ME�L���,GɈo�e^�+�T�?�y}8��7��h�`w�ץ��MS�c`��[ƈ'��1ъW:�c���/�ߥ��/�=2�b[��g��j�r7V1M�م�݌��|��$R�1���9�uc�P{.T0�=ȑM�tj#dBD\�3ul=�2_�ó<��MW�r-c���-�����wllD���.��:*d�g!}R0�qC|U�������3�C���C�7����u8,1�F?ύ@B��RJBg�9�iD�Y�i��W�}�u�?�s����s����`؅�Fr� �z�.�pL�kn� (�iD���3�N";�§�mu;�QV������tU�A�vn��K�I�S���Λ�J�-�ۏ�&��R��JJϚ2X��ʾ��Â��b:�]�_����6A��}��_��_F����@��D�4j:uH��T�@
m����^EX�j�&�w�0s��=.zc�<M�ȵ��� Q޷�Ss{e������������Ķ���r���#{��9��u1a#�����LKص��E3O�*47zvq�]q}X!3���}���l)@v��A'G�m�ct��%�f�=u`?�է�߮^S(qP�qt��5I^i�N_8�$ Hjy<��=��\�k��϶uT�w9=�l�������?��`)�)e�-�{Uw�.�l�lgw���0D~ת�'O�G=RVmF�;�8��7z�<\Y��&�>���A�ۯ��_�VU@����\�4���؝у�dF��}���?"@��0	���ʳΕ.<F5Y�X5S	�ZVl{{˜�ъq_�Zjۮ��m�"�������0�B�k  �R̐VMy೽u�u]A4z,[�51�7��CgD������4Oܶ!���,J_�[����A�� ~�<@Ȭ	��y��9����x�t��pR���`���.R�Hݓ��A����4�Lu�9�?�ss��.t=�pԡ�%�0�ѯ���`����(:U��m�_�!Z�Y1����r{��zT�����[.lSB�y�jb�9��Zc��t�w��"�_��!�'C{�,��sлK�g�{��W(��ro��$�/3Q��ĉ#��SnH��؀Vh�1ӥ�iu[��ڥj�T0�U=��/��Pm�F�ԡƄa!T���V5�<Ewn���VB6l^���'{BF��[+A+�R������J�!���^	�fE�S@5�9e*,�.�PK>0��&5��AE�U�!�˵i���3m���u4��nd�=D�^��hG�;.Tz}'e"����,KG3�@P`6H7���^��* ��HL�/Y�,��;�[y�]�翘.)��hc�ȏ�&L�N�t�`H�[�Y�#�B
Q��=~jX)�V�S@��a3�u-B�cEk��lHF+�!B�b�nA)K{6ω�
iV�FW]rz��ŵG_�y��LHp\gRq�k�UVc�
����ô�j��y���G�E�[�Hs��u5�n�8$}���a $�����\�&_�E������^Hf�	��f�~:9�yF��*w;� ����8�"���p�E_�5�ͧDd�}D#�L�/p��_O���~.^��ƛ��p$A����3�?��M��캶i�͵,���3�|h���`�y>-v�a�j����f�C)�v���<!�ќ�R�m$H� �4�3'���o��&N&�j]�2���j��~���S����\Jb	Z��E�jȜ�H�j��F����#1'�\�|��]��o[�ω�=�(��3B�A�hm~�]<Z~���G�����x	ۗS U��0r�:�}���\ =�^�%}+B�l��s_+x�vn��{~LFc HR�%(�\?��ڳH �0��kY�����ߣ�~D�zdc�!A'ٯ��eF�8�~�sKx���ӭ6\!�"p)}�g����3�5��\Y���ƶ�~��èY��0��8c�iC�F��8��,aH��m˺+�wtq��~�b�ͷ�KfM(	�f���O��3���vVײEX�������t�a�HC���Y��ê��X���W�Z8ÊA���|��t���򁸧s2���v}�Tu���DJ��qr�ݤ�] jqO�R�΀���E�)��N�v���&J�����(>�/+�*Tb������H�v��^R.֧��n�����c��@��l"�7�0"����œբ���X_�~�U�����!�9ۖY\Nf�bl߲H��¢Z�#�����O,�U����j��H0i&o ���*�,Ls��0�JI�$���?):ϭC�����ԞJ95ӬR��K����%�O�Cy��
�9�VBPj�;�OЭ�22)����G��ᦇ$,������X����X��x�s*Ql�C��.U�W��'!pw�n��m7o*�b�o��Z1 ��-Ǡ�gI�ֿQ�<�G��?��˱�A,n�x��$��a�<���4P��t�i��� ���'0l��W#��L���ND��R9�3!�H�G��Y��嫣o"��K��n�c�u_FŲg���k���ƽn���ٟ(���#�~���V�﫪�GkT�A^N��
o��@�vFc��`�/-�]�y
cۆ�֐�m��5���<ȿ����n���A��{Z'�bh����)�əEx�)�~��5($�M� ����7G�(�B���a-���5;i\�iV	�wE�3�̨`�����xg�RZK"�`͗6$~6�&W��r%��(�s��L.6�)V���/�9h��R�{���A��\���d���1c�mN�E�Ж|������f2�;���cc)�3>Oƙ���n�J/9��_.���F'��R �쟯�TpO	DKC���7f�R�L���i��-��\�R�{3� �+j���D�I�2)��aGG�`�/�º�������B׺���B��sS�(�:=���B0b��l����Z^��յLcT�W�+��B�Y�����F`�����%Q�����J�#�8s,c}�'|1g�NnOL����2��tQ�	T�!Y��7
��c���e��
��T��Ĉ��)�s/",��@�o�%[�PsC��d_l���$�b�E�rd|����\�ܼ�K����$�J�uҙf�E�����?�^*����ߴ���F���;���+*�%FXv��)�o�Ua����U0����l�󍩱?�yZ�G;╆�ib���.��#��D^^�gw�r>��Sx�$�YxL>��%�eSP�<`��m�P���.8���IG 8c��Uq����w��,�I�'yH�N
S������⮹����8�2Q� 
���%F�4L?dh��x�%9��<���Ė5�H�)�l4�g�|��G�Z:sJ�B��l����8����ź\�F���U�gŖǷ}OV9��ᐐQ|�_5�:��� =T�x�X���F��6���s��t=�v"ó���?��ҔwW����cˈ>`�LkN/� p��M�+����.����^v�LB�R�M�$+O�Z�O�fAE0���0�"�)����?�5j���!|�q��)y�a;T#�v`w�Ǡ�oRޓ�ƒ�����GO������ho�W�H�M��\jg���{�4��������^4a�M�S��6���I�իs���Ǩ"a��<���4y�����d�ˋ�W���b���Oi��h�*�T�TEj�_ �����!���x��8�<7S��$�{\�-5�t(n�1��,I6��198���_#&S���`?)|�s�;2�
�k���Ɔ#G�f�������ξ��Љ�����.sg^��u��G����$Pj��ߟ�Ŏ�\<����βz:�F�������<����W�
��A�[ `R�R� f'|�D��
Y��Xw�]�����y�4&��ll2�p�c�wx�$�̑����ŀ�F>��n���f
����pP�0 �#i�̤4�_i�6�`��V�W.�JY�7Q��<�`%�s�QhX�#��C��|�mϘ(��A�#y�{��$Cv���LR!_�Iq(��E%	�o��C���?p21�ȗ�wކXB�-kl75���}��6���9��n!z��V/�Nr�hd��o�p�li��aa!/t��T�p*Y����w���gg�1u�#��Y|T�7���hL��	^�{Z�"�lZ�'����F/ױB����M���h�C�?�D�"���e7S��ց�@�,#.Z=)�ݝTP�>�"�cȈj���mc�)<U�תZ>�{:e�oV󘐎��oL���F�i�L�!,�sgCs@൯ ���_�u�vR\���Q�;y	V��˨?���|����4���Qц�]�7.�/���(O��mb��.�E�qS�'6��Ҋ�!+� ���aV�@S��s5�K�1T�@cږA4��|��)q+ϒQ�N� �l;AZ�}���ò� �Le�Q.]=~���A"�9���!��Ii$���y��[���g��(���Bb�)��3B���(�t,�7���2֐"/�H�pވ�3����e�$|~j$�D��9J ��Vi��$vW��@��3�;���]A�`������j��ڀf�}���k�y��	>F�t˒�&T�s O3
)�vykٻ#�._Q�Ģ�(rԚ��]Z���x�\� �r�b����p,OO�q�4K��:}�u`����ȹE1�,.�ja�|ɺ���\�
��Be��F�3�m�ag��t<J.��|.��R���$4�ؑ��wg�eM���R�ĔqP��N��'yG���YJ��lM|o?��6���W>8%�q���m��w�7����$�,�'{�yӗV̞Bt�^fx`��|���8�m��	�EK~햔o�R��ߵ�9Bљ��g�vm�ʕ��3~�~!��������V��X  Xk"{�{YhY(-���?~�:�}e@������a?��3Z�x���kV�ۚ�� ����/R k8�Jj�fN{��ވȶ��S9��i�-�9�kBd�e����6�`,8M��aWlL̠��V�[_�ul��E<��J��9��x;�^��bs�$��V	�S������������h���������I��^��Ӽ�1N���F�sԟBi�_x�Vޅ��վ�S��*
�R-�$���f���,��?V^��g�j_�z�y�"��_��OV�	���Gk�����w�v&���G�f3:�٪l�b��w�2����쾋��@n�@v�=�yb������0ʋL ���{͗�Bn'�*�%��zCp[5�Pi°'{'������u����T1P���^^�x�JJ�{�)���A�6��@e�=�� �\ر�9�j��e�JƧ�����Da�ޏ3A^�O�PpW�Ө��ӹ8�ORl�%�l<���t�0K��*ט�t�^H;is+W�u��ol41#gf�ђ�-�����$�U�TWT�&���x���<i����	�"������vXt���&(l(p��c�ʄV���R�Ͱ�\A�\zuLQ9I촀�~
(v{�g�h@Ԃq�ĉ$�#�^Ƿ}.�a�A�O���2�D]j�y(Mȡ�mq$r+��eN����Ks^���S�qi��(q�?2ʆ�����-�x@ި�9�W7ŘrzW��� �=E�j��_���.����]|���Hn:cE8��^� �T�b@bl�/E�!"���i7��g�7]=6��T�
�'�8��l A��4g�n���)�7�?��C�; � G2N.��@�z�bя�Ȟ�C���{WK����#��M<4@C�M.�M�*y$\��1�����pY4톐�4��q���Χi��V���u���7U�|�n�B�E�ts~t<�yin�&V��8�Y���I�?���nZz�[����זNYD{��ԯ`�`��%bs ����B�@�F���������1������d\M&b:e�ߨ;��ͳ�`C��TT}�ug�X����.�E���?=H:;J��4�\���g.��!���\��	�D�9��w����g�����m�$�U�\���>s\]�P���eR�j�؆�K����/٪��� "?L�
�kwQ�~�8�)Dfq������w*����݉����0'fD��|u��"�[Ŝ���Q9��c˂t��o�n*I��M��j)Rn�D/w8�O�����9e��>��|�����l���y���-l��x2�.*�$���6�Q��Y�(�7�5��b��\�+;.�;f���T�����z 8��E���$/�G,`�߈�`���=W�B�A����r��G���V�	w�x������ }�5u}�5�?�����z�1�},������M/�))[/�MM�A����_E�����0��u���0�_���(YTy�(���M��"^YA��of�Hk��������p[�mig�����nB���1^O+�}_&��v�QXO�nt;�k(vB�o���H� �_����h`��j��UC��68����US�P���u(.`�sA�
t�A7�%׹��C~���I� ����p�NZ�߭�0D-:ĭ,�����нR�]��ZC001t$��T$0���%�|���JNN�Hr���B2߸�A�z�p Fs(X��#��P���p�1��Z;��28v�Aϔj> 9Mt�L��"�^
��/H�Z�A�@��Z���k����o������?���Dh��k�<�;�h��k�G�$4삉�%���E��o����f[�W`� �^a�)�������uӐ�:��k��e ��g���U e�:��M�۬b�::�.q�������T��r�����XaQ;�	]5��q��G��U��N�&`�G�0yח�a����y��%ί�J&�~��pJ�u�
#,n|K�M�o����\J�Cp�\�^X���������y�O��}h��?��_ܠf�����W3�8�teT�=�6ϯ`���!3�S�r��m�+��}Di�i�A��@���V��+�Hw��#S1O|p��^@#:�4�+YK�����ۑMj��v�C��+�5�~:�+̻�q}}�[G=WH[7wU� l'@���MiA:כ8ySf v��-R�X�_�-����*b��@xm�����X>��8���p_ �Uw��G3���A���\ɌE�hn�q�8��(ux.�V���/��)�'�@�釱��ny��!&b�Eo6L�fr����u˄��گq��炼Z�]�կ���m̠�w�am���1D�`��_6�}Ϟ��1� æ����7m՚\�<�I����q#�&����� ��lU�R~F%��m\У���t��{y^�:N(?�OKz��NO��F��$�ί�ws������?V�A��l��(�g��!	�������?H�nKDǻ"@,l���e���xp�9�"�w�kM)FK��^�e��ؽ��7%!�EB��+a����A�P��>�!-������#��C�]�_�S�Ȃ,�������>�~>�YfÛ�
���h.J���t�pwTr�u��C��i&��q��c��A<�,p�i��n���D�p(IOw�*D��tN��֣X%+�?��o�:r, rDh�&o�@���t�#C^̽n�-���j���}�*�}���:.@R��k�I�_���S]��Ж<�R���5�D�([�,u��x}�W�������������L/���m9���E�9���h�n`]B����Jњ��"���y�~ДM�v�y	R�ʤ�o�lb��x������r�R���������ih�f����r}^\8_�ER�(П�B���&�\3WA�p�l8X�`�'|z'�u�Zs��h�gx���;��B�����|O#'7T[��
UR:��t���d|ax5��~��&�O���!^�:q��!�P1�r�(�n[H|i��}���5n瘘3�)(z��0�����#d�8a.�H���ZvK�2h��
�R E�P��]�t[;b9#7��.z¦��H��l�@���A%�؈�$��"�!��XC��A��%4� Oj Aa�i��'�~r�Mћ�f���^��a3`nu�T�vzu��5]qYk
�>"���Z�t89�}�-�C�cy`
7_֍,T��t�1"���a�^:�/�N�6�)%��N&��7��',�ZmG�x��.<�L�񵟐	��G�*�:Q�ƶ*j�T)������fb������� �<찿^S`�r��3l�
N<��{�3�g���sIΘV�ъq�J/	[e��\�]���5���W�[��ƻ3#d���:x�
���� �tV9h��⥶��t~�35��O8b�f�rIQ<��o��S������1�X�ѽ�^����4�)ǻ��M<[t��I`�{���N�����JJl� #'�7�+�����l��ؚ�W�6���@9���(�%�.��c=�/�'*��F%��7f�mԎh�P��$�¾�S9�
o�������wH�X:D}��L�*�%%ED���Q��?mGו��@�Y8�O�R{�t�*�?)��{?ۘ�A��Zw@���1�i���ckj�:Ŭ�|0�U����F��vא����e&�|>Ei�y+�?��35�F&K��?ڄ�!�"�@�\Ò��K�]7�$��1o�D��I������]L�u3w+k2��r�P )���|I�aaRMC�<'��F��K�\�x�N��!LXzsj��<�f�	��������5Q �?�L��qw������]��s	n�����2��*ԝݗ�0N��l��zM�@h�u<���C{�y�\u2uM�.�T��{�&�>Rg��B��ɕ�@�z tá~l��"� ��^��j�?A������?��r�LTB�9��q�(w���/k,�0X���L�O�[�I��������*$OM�q� 2��θ'��ό�zZf<��P�C����\Bϴ|�~uQM�D>���
����q�ee���חA���f���l��,Ҹ��A���Z�r���|$�{f�J*u��Z��SZ���*/�IɈ�J�VQ
��I�z�� 1*���⻱�8)6+a��E*c�D�|t�1��T_iyCJ���#�N�_$�#5�e>�� eȔ��,�׬U���\=��;�]�Ӈ
�5
ӣ�)���|��Fbr��U?�x�0��c�d#?���x���m��V�6G/���fq�5�]7�Q׌)��{_ް�ԥV���%`���	�*$U��/�AKzm^^���SgWs���{��z�p��p�J6+M��߇� �S��e�Z/��~�c�<R���_�5�q��9��u�	�#4*+�D�!���fς�`HFuОq3݊��$)�AH܃Z,��g��#�G�OP	T��b�KB+]�� m���9���y�ևC���\,��(���/�ge��F�az5�#s�Q Qs���A�<��[M��X/JqQ�8tk��o�W$�SWvm���a���+�������b��W���W����фq���cu^�g�?�һ���]��FѝΟD�Q�@3�#&T��xs��2��W��Aή�2�����_����Z���lZփ��h/^�QonV2��*�%����Ǵ.fS��u�ãsj{� �#y�q�F˟)����o��RǟIi���P �<$����F<�<w���&�;P� ��Np�܀�L�������Ef�� o��qHK����s�>!d:R\ؖS�G>�Z��D��{�Q���r����\�~�u�رx� ���.�j��? �`_�y�jl�'|�∙���A�О����:z(�ؙy�#s�z �T{�Dw�ᐮ�P5���v���+c�'Ů<vs�;�D�X ɓ��E*O���#����@��	j�%,��{NbG9�t{��?7�Bb}����c+C�z� ��=���j4��$����}��-����N���������zi$s���Z��P=����>�2��,�+K=GܷZ��>��)PA�,/�ւ��#����' S�Q�4ޘ�1��CwbO}�gņ��泘�,)�˲���5X`Ç�сs`�7j���o�����,Ԫ�\�厲՝��L�L@Ԭ�D �C�,J�r>E`��@Q��j"2� ��m6L-te���ْ�.['l��b�"����|��x(nq1fN��4��x�p�Zn]?��0İE��ΩYPً\�u��$�e�M��m51.S��0X:����ٸG!��
v��ׂś�ڲB){|H���h+B�uΟ�����t��I��g�}*C<���y�>2s[�T-��ۆ�_x��yv�#� ě���d�t}����TPdh��<t9����T%�#@36���6tuʷ�G,d���j��PFg�fm��Y�����Y;���qKa9F(�O�xYYZD��lI�L��3X�&ԇJR��DK�J;�c�h����g�O3XзE�2J�<��_��� 6��31$�X'���G~nT���>=|�?6�ˉ/�iu�>�4���t��yU^��Ms0K˸��z(�8H]"L��l��O�j������6�����J},��D���<@�B�@�4:*��IO�di�z[8��$Uf��d�o�<�4�9A��Դ����8n��c�	 6AF#��������w�� ν׉�I"��İ�@N��IJ/S�(��$����.�v��Ӆ5PC!�>��3n��MuI)��p%dm���vmz�v�8�ꋽU����������4�⏉�W��^͚	�xY��ӑ��<ʕ{��b����
��\���5�z	iB�`��`�Zj �eB����fK�v�57L6�t�F=�2o���H=�㸪J5�h��(a.���#��9ƊQN�����:�V�����Pd���<��_����k�i�KqP}i~�	�5IQFq�R�(Z'����-.�>��ص��}eH�H��+la�`��AړG�f��n.$C&�n77�C�YK����{�+$9r�0���P��~�t�BQ� �$�S��)^���@�I��I��oC�Bc�7Lz��q�!$�%*D+f���bZOu�klv6B�&�� ��K鑶g��9�ȌR��t?�1�({t�Đ2�`�B�����2n�Nyٚg���S���TN�����z���h"�J���N{��f��]��|%����k�;j٪�p��V��T@j����{�p�r������8>x���� ���	!��.������73۳o�> �8���H��x���Iyd{-���i([�<�k�塻�`��~���"y&�wY��K���M=��b�Ӝ�q�c��)������͊?�KZؠ�R�6�pn���1�1q� �c�:o��dnM��Ƴ�����jƁ�.�����E~w�ꚕ�M	���&B�E��Fޅ|����_f�j
"�7-w"�\I{�<�,PN��8`ױ�~e��d�V��8����{�9�������UM��ڳ�]�yD9jPjA��߃��>�1`���-~ltj��	s�,kE��I�9��lw#��=@P�)VY!��fi�P��O"�u��ׂ�gXǭ���=Y�r�4�N��PtC��-M�l#�k�!��Qc�0�Pw*=���9°��������R).���f��*B�X��$���&�	�R	�$�����Ip2��m�3�S}L�w-B�"<��a.v�XK�m�bޞ����a962�7�[�2-��{c�T�Ye}�S�� f^�r܈�s�<���k<�(��/R�#�#<��=�sa����|XLs�@�{��`�!��=ya"g���j�ce��0�oB���a��y�{��h��KR��@y�=}:�|!�&�KkS���D������v80ooK0�}���V��HSy�|�w<)�qc]3�!s&��0�C�l5T��t��A^)!��ѻ�a�8��c� mQ>0��៯@�B����\ �n1�H��:g23�ڌ���[ �<$���p�Z��A��K0~��A�}j>�>��,ˡ$r65+�Ce��
�
Yv\C
%�\� �ûH�}�5u��ka�P]��� y�}��fA1�RN�S�[�2T�1W�<�"�����G��l�ݣ��Y�]0n�6��xm� g���C-�wB�Ց"�ǣ�i{-5�2��u��@�ԸY7�jE^��q���=WM�NM�����0|�
�����ƶ&-�����2��/���'f\�K��8��1�������c��bD�,����	eKv��=�eNXg���k�c���3g����s�3� ��N_
�Zra�H�C�j��w�ف�劽����Ӳ��-G�6*@�5��mF\�u�Qy�d�g�������E��uTD3�U������[��H�k�zWK���sC 0�.屮�p��ϺoU�d�Yњ�A5?�K�*��w][� A��b(�x�a�5��AGƺ��k뒂��r0�-c�6�s�ue� JO�A����L��qWN �L�M��O��А�\�R��>�-�I�zt9�f?e�-h�K���c��Ma�����n%Y;��#�d�ag�:'�d�\~��-�3��b���C1l
�|l�ĕ|b���&�����U�ˋ��s�%�h�F� �x����A����TuO�i�'���v��ӽ���<J9�j��h}B�d33dT�ֱ��h3\�B���u�E|�Ј8�zh��J��in X��:+�㳠�r����<!.NUͲҲx]K@��o6��e��^JI������6𾀶�@;���:��a�5��Sgs1������#u6g���E���M�b��3&ݻ�z�{�}>����8^�F�DfZ%3�����_nx��6�����g���i�#bj@��H�7�����q���Idq�_!m4Y�P��+)��@�9Q��:8���P����l��"?h0�t
�]6[����s�?Z�"����������-BuzfR6��1�-�S�\:���_n��ۡ��(���$j�܅S\��vnu�N����@׽������]X�?1 �(��AZ�	�Nr��]�
L�[�!�DM��zZ���2���6i��Cs�ə|]�o��{������2�����k�e��n�r�aS�v�#�z���F�ږY|>��� �\z8HN����*1$ˇ������o��!s�t�`�����7��� �EyՊb���<vվ�.���3Gܗ�{R�d{C2�Ѳ����l����;�R:��B��=��hҞa�����}T6]bO{�t�ٖD�O(���&f?�j��Y�!zP���g�{aT7*Zz��G�㩮�����<1΄t:����k�ݚ��#:�HJ�=��\4pq��R��;����"��9�I�����3u�ߨ������l���V3�q�~sN��%C�pjy�e�Ռ��!�8�S��O��C�g��o�=�4�,��ڐ')�k�����d7J�?:jm!�X�Y~��S���iunM^�%���X��n����jH�P�x<:��xh媹�t����x�"}�J�1��G���Ƚ�k���������a���+U�>�k��f���M�����Q�t�*�x�v�����?�u�0c�_�pQ�� 85�������X�7uE��}Z�T.�o��b%�����J��X��0[I���X�C��Q�`��G�N㩢.�����&��p�!��~!��(�&[`�3���my̶��i�ʤjA�j��Bd��K�+HM!S�ܶ 1�t5�ҝ2$�pˍ�5Ա��t���Wͦh��f��<��c��1#�\���|`}5�?5����ic�
�����]B���~9fP��p����b!�������Rt��<�̭�)c���,���,A��8��Zi�*�`�JC�����%lDE�ǣ�[��+5�"��+ơa
����E�(yB�a�	��t�zz��Js�6a�Ez�Oh����Y���юA�o�'�Iw.���P� I�����D7܏�,˔$� ��f�f� ��>�p��A�R�.3kʪ��,� �Q�z�
k���ѱ7riP7���n���DU�����B�Q�V
f��[;��8jb/�;��vj�	0�i��Oe��ܧ�S��@��l��O�$U�	|��Hٛ���z4zɅ��-7(݀�ȍ(�m�Hjt�{s�T�S�PQѷ��k΃x� Ǌ�K�To���^����hM|9�<$���q�t%������O� �BQ��s=
[ao\)�������nU�z/a���m�A��,�|F �
&����s�����g�V2���;��˜h/b
�,q`���$�<i8��:%�j~4u�!r���Ņ�q��:��$���/qC�|�S9,���H�Z�_�n��n���@k�UU�p�W$�vt��Vaa�Y�����>_���^�p�f=�򯝆*��=r�~*��� �j����
�]�������i�y�5�Rˮ,�>�@1������j���|k�ձ�fs��z/��҆32s'�y�0+��Qt����D@N��z}`KyfHCR�
i��{�['P�LP�Q�7=�r��ʏ��#��� u�A���g[�#\�I�6ƴ���`��d�Hn�g��K����-Tuv�p�9�__z��V��0C��S�Ϭ�֊4���M�7��턺���o�_G5�t�	����݄�l�g ���3��0f+����(�X-sd�oO�48V#�#�ĒS\>F���t.E��5n;��w�3�.��]�ab����C����� �m����r������~��+�c�C�9-�lO��G	4(��w *<)�+��o���1a1��-V�=;��
Bq�X=5�~��HӇv��$r1���*ᗅO�[A�m˼IؠM��.�bԃI@Ή_� ay�e�Z/@��"�T"t�fc¨��� lb̂���"-|(�c�,*��GH�	]���al�[=E-G�a��gJ/�\2T�/�WU�D����4����laL�k ��I��j��@[R.&A2���ڦ0K��5.G�O�1b���D,��.�K�D8`9��:Ҧ���?���o%w����be{��O�ۣ��.���DU14�F�}<����w���g�P�A�u���?�]v"٬a��˩����!�>/W���逋�Ғ�-������>M<D�: U�_�3��E���e��ըW⋳�1#ipK�*E�����Y0��������m����3����,����J���nLsJ��'��j8��2ߐk��0�3����-D��O���EWa��XJ��D�S��K�c~@�d*�>�ǁW�X��.���$��֖7y&���1in��7��E�Ѻ���Ϭhʬ¬�Z(X`���r�h,�NM!{����[v4��<���O��8�c�X�**R�'.�� n�Sgx}C؆~dyQ���4dɬ	��:,ƭ6ZN���+�H5���a&��\mPY������������U?���T��cU�P�W@b�m�)��4���eOǄ�.J^FD⭖�Wj��`��nY��W	<8��,�&6�Z���#���%��3���w1���u����A���x]���g�9�8[��j-�UX��\ _IP\);�����=9^ƗC��p��৫S6�b@=^IyV�ٓ:�&���4M�[�� �s�����t������&0�ۀ|�\-�EQ���v����\d:K����օޥ#&��.r���z�O=<�`W*zG����HF莋�}�>�)J~�%3�X���/�m�@�Aُ�5��qE�韘v��G��k�����<ckҟ��}����DF8?���-py%,��>'�:U���?��KsJ�4��O��$�gsU��eB�KL)Ӭ���\�@Z���U�L�z>w<���W�VXa����~nA߷����%и�M�&EYY����}f�]y^@�:@{¾\�ʜ;v_��5R�5ju�]�_W�XF�ۿ��; �5E+'�����U��sƣ��Xp k�~5�蘧�K�Qf�H�U ��P���&oz`H�$R7��NS�F��$/��v���`Q�H2F=�W�BW�SZVa�]d[�$��5���	�o���?⹭k\y��� A��ed�:����e�+@Oq8����Ja_�H�#گ�o�K��n��\�,w�c�:)]zU���]i1����J��P}�R/m�Ź����ϰ��B�2�H�U&�~�b�H��vi���2s��`3�e=�����YO#c`~�v �J=��N�㑈*�6��\`ߔQJ��X���_^+�fuu �"',�n1>���O�H>�T=�&�\FzT�0٫�F���Cھ*mg�W:x����������BMuު`Bif���u��\{be��1kѷ�a�t��8���7؏�Yfp{�Gp�<�۰?ko[����I�O��\|�����2����[�nU����F���l�Tt��>2� U�P	/��v�7��?�b1Y�h?bl�G�X�swU��Lro��כ�-�<���}@��j\�}�D�H�����(���$ҿ��
�����̌Y\�խ���*��ī��~��Y��5Ǩ4�C�6�Q��QL��fʁ���$*+�X�͠0C���)��%�;u)�ݘyW�Y#0�Rm��Q�$3|�-��C��؟~�RQ�:������N�y^��ID�ttD�r��1����P}��N~�p���9�sV'���9Lk�y#����)AWG�,P�!�I `��E�D��-_a֧�!|�#�O����%�1�&W\���t4$}uc4{a"�(�3�#����[��*���{�y;��I��!- 1�ȸŤ��3h,��I��\�]'�t�N�3�ς�W�>AH��6��z��oȥ�t�:0�Wp?�������]w�9A��Sx��0�P�>F	��k����pA4�|雜�&�վ���s�1��_�09M��osG�>��O�	.O3���?���I�����>V�1��{pM/jbvi��#�W)���24֊�j՗�b��{񎧤��o��IlK4#q�h�z�w*ݰ�����YX�jw�1l�����0wĿ�q���)[����a�)Z2s?���QǛ7�	Ө����M�v���`ȿ>�R�Cm��	F#LBɧ��;��1�z/Ɨ<��`>.�p�hgڝ�`Yi1�?'(՜)vW�6:s�i��<�����/��P$��.���vvp�c<_w���!T��#�P�*�~{=��+��8?��k��v��O��l�;դ#,ۏ}v����.�0ݰ�,��hnrH���(q�([R����!p<0:r�>���E&Bt�%�-<�ϝ�ϥ��`4��
g]9������FqN�ᚏ�����f�g�CP@M�lϟ���c*0-���D.���Kv���������h��d��L��I�I����ꇺ�����WS���)�7*
������uI��-e�I>W��q؊�"�dS�/?^���L��g�3L/�j�欬O�¢��Kg��HE�/��<f�߮���B�3��
S��ԥ�,b\]1�*����=,�/v��Ym�4�jG��h8X��xfH�[~>��#-��c{��b�Se�G�i5�
lQ
�#11�����C@��b:wf���K�6P�5�N���I&w�O� ��& 䞪�O����z�rD��^;���iƐ����Y=��wY]R*7t7����X/.��Jj����׆T�ѫd�}��(mN����8|����¤��+���C�%Zb	b�6��W38�AW�?Ь쭀�1��)�+w�n�dy_>��o�]��.Ig��-�=������L���B������=��-	M�Ev����M�/T�	��=�)c`T�&8<���W��_���������P"�5ơ�\[,Яд<���6f��$�#��z��
�x*w���`��4�܄46��6�j1�#�s �N�kǅ/tP�ɛ�g�� ��V��N�l� k��p����o �~Q0�o��cK��H%�r�,wn���*!7�'�0�`���*�O�L}-0	����=b[�Rն+�6���Jt�M>=�C����U|G�6�͕�!�!���C��F�I�mlg����Ҵ�4ݟ���yzAu��|2uJY��&ܝiko�I�pX}�}�&��$(�m�.�Ȅب������#p9O��ۑi����*�-��wf��䙛��0f��V7@�Q�~�I������$�@X�v</}<�WñF�E�J�!�	I��h�Y�ʙ�Rz�Wg�{��sn�X�{f��5�me�2�=^O�i�����Vƕ2�_-�����]Q�2��?w?�y:��n�#]�Wf�q�ަt��Z��z��N,3��)�JZr7'����R��1/�l�˖S+!X��!�/C�5�=�\�J[����B"w���p=���i�9���n�_�6
d��k�v�<���:+;qί��;Q�� WY��e�E�}N֨�X"c�&��X����%���J�K|Y��i�5 �P�]\� O=¦�n�s`{S�q�� �b���Z,\#����8�c�ʷ}�d$�e�p���£��0q��7�yX�$�$�w�2CPe#ۂ�o�eH�IG� ���_J��_㐟������à*,(�d>C&[�)h�0,��щ[���߾��]q�ߍ�>g	�4���8�YB&�q7;���)sW�' c�Z�<��U�hlZ
\��,�c0pQ�r�2C,���x}�γ�w=��SRl���ݢ*Tp�+�.D[�p.��Q�&�Cgw�B�l���b+6��8������\٦p�r�qCRp��ze�w2౫�FR��p/�[�:(�IĢ�
�gw�W�X7�9s�CC�[h��~�:���qf�k�#��+�ڳJi�/���p*5��O��?�G9J%\�3�r�j�:^�ꤽ��ff`Q�}̯�;�u�g��d��Ϝ#͗����J}x]|�5��:ڵ�T�\)�s�Fݹۋ�.	�wM���=�-6�f}�ȓ�1��=���0�5���1hog�Pre?|������鷇��M\z�����%\yi���d�r��E�!�����Z(؃����p�U���qi%'d�_u?�d����րU,��}H���5Elp7���OY�_�u�i��L~�%�'��o�o�<��
�����҆�(G198�.�cRK"� �9��T�,��i�Q�sw�3�^����L�f��k�lA��$�]��q�[���T�0�����A
��I���R4�تW%@��Z���6۰��:�c\��L҂_�n��;��6���SЈY���<���*;7�&��iGB+҉�VW�>��v��&/���\������Y�����\@����{�9ـ���g�aEg�(�ߟ��������L��L���t��c�w<^ɾ�>��QU��t�'c�@wE��D�3�`l���[*R��y"���o�2k	S��Tk�"����I#F?�u�s�lYz��wIy��|x"��-݊�0j�G�	���H����E{'[�*�wϿ~�"�D�4�j�s9ew�Τ�|G������:<�Z4���4׼���Ϙ̤�=���p�XN:s�\��7�Y��H�(c���%
s#��6�>閟���D��._�����w���hW��S��i�b�%j���;V���d���eZ�٢?ۙ��rξ�����7����W���@��KuJ!��A�|Q�=4��%���PėʦAy�l�.�<�?<AI]
C��Z꒑	�rNˇu.��N�Pck����B*�pΚ����Ʒ��W ����<�]
~�D��V;���I�T�����K�Li��P�H�r����䧎�,�B����¾���reͶ�h�W&H�Q�[�P_6�~��rH8�W���q1KA���u�
�+%���.�&��Lw̖ԕ��V1�x`�?��:E��md�[f�/�Ԝ��e����c,����g����LJGڻ��0҉님���jM���֙E1{�'j�R� �+$��B�e���Lq�7�ңZ�5�Qs�g"�G�����qݕR�0 ���R�y]����#)K�V�1��q%�9�@2���^.��=W������VQK�B3[��GC3O�.c�W�Y��J^�d�@�৻+?����_�e��s1%K��G�����V�5$��h���A|��
q�0[W1G���J>w�y��W��=����ҟ?��hE�TA%����k�4@[��g���ۏ���O�'�Q�^�@��@EH���q�A8W�ӈ�_h��*�L��<�������!E"�M�V��1i�G���A�����	��E�6G�:Lh_^�a��8l�{Je���<�L����>��Ի�-]��������O��'���9ݴ��C��
���R�*���A��U�q�y����R�G�}�������z�#_fCT�5}����9��V��s�����^��'��**����k~_r��.>��6m'ZZژ���c�KKw~f�Q�/ieO� �
b3� �ys*��'ڈx�;e�#5C�Z�)�f�$Z�z���Bj������ŀQ�2��J����눫��������+�� Gv2<?�f���EW���O�H��ȝU�����bÉRY=��έ�'����tg+�5��:�aRZ6�����e�b�!*�ekխ�F��8�o�N5�/y.*E������-�f��@'i�>���dp����_%�E�
̫~���Q�o�`�Ԯ��׉_�Fe��C�U�p ��O��9�۷o� �@�x,	�Q�s�*����8φ]i�.����'^]�\V�f:l�n]k
�/w�R�k5c{��>��p������F�(:������>��D�Z;��'��HLw�;-�'��N�'�H� ��U��f16���yj�vyV�����r�����UW%�����b�M�!]h�=��`F�(O
f�EQ��8c����S�N��{�,V�^"ԩ��w6��7x�Mg�C�Lh�g������Lȑ����3���tr�uj�����NT�����w�{�q�X��9ӫ�*�?-�*�&p+����dt�uY_�.�q���q���X�����,��j�(����#�J�!+�����~�'�Eo:�=���#�����X��c�G�K��"��W*���Ir�]ŋ�0߬�r6X&����S�C�5�p�w.�O�Ի��V���U�
�&PG��_+�o����,���$�W�EY�>�r���M��ͻ���Nnzu�E}K?����؃�M��:��>q���m��0X�¾�9���Fg(a,���'�b���vI���-䢴A�94�U��d6�.}��v�vjD.���e5��lY��FY��qLs�6�̽����Xj]���M1"��
���v�v>�.���	����w!fqf�x+n���aK[��U�oZ�o�-��
�,O u�������7r��zu?�`ϙ<�"�T�������y�Z���#Zb���t�gv�V�٢�_�&.��Z$nږwKӎ���?@���޸d��O(�Q�a��37j�0���\�$9���,�%1�O��ȗ��z׻�)�Gl\�A�C�a]6({5X�К�+�"�&���e腛���W��eԱ�*�D>P�1i:�g5��(*y��#.(� =y/��vF*�D�-��N���˭_�mUEM�����`��T'Qn6J��%�cןZb�/c�hn+�^�+���/�ˆ�uި��{�y7�LH����VUŃH�:c��3��sw��y�������)bIK꟪�5A�̤E�K{HXtu��R d0��z�_U��b �$z����hϗ3��#>�0�o)t�y�j�����f��H�KӤ�:ʣ`i�H�ϓa�[r��;h?��G�Tx�����ܟ��e��2kmJW�]�~��� ���db���r1���-��ұ�MQ4?蕶`��O�S�2D5��>�bKUYT�Kn���)A2ś�6�к��߉q�lc���[��$��!�D%����(��Q�a���uF��xMU������_v�.g�ｋEpQG���f�H���%t �.��X����,9�����dV��'4r�T�j�f�fƎ%,P����-���<d@)�˟���������އm��lR�@�y��k�it�!p���T#�]�sTL\@CC�j%��Ĩ�:�N>�n�s�_@�Nr
3��]�P��,�6�
@�y�D�ly2�pS���U�޺�%i<�����L؉#N̅և��>P�eT��Ŗ���Ε�V���:�G�ŋ�U��;q��h/���b%�x��P��Ә*�.5�i�k	3�ךi�7�����|-��E*��]�8��\����C�{.Hre|	.��y�8��bZ8!gE��Z��3y�{�柿r�c�'V�j>�_a.��~%rk�e�7�M�k^�(��ݑX1��g}�]�'Mq"����q��B�V���\���UX��*��߂����B���I��#Yj���MdK��t�#|��bm��Bq�dܹ��ɑf�7l�6>���L�,n��b?=�pѿ_Ê���U��hɂ�M��̱�[�;-�x6���.eh�F^T�f�6ğ�#�'���	S���a�U������	��(�Bg�%Ӈ����~2m۬/����O�����y"��w���Q�:W��u�7?ײ�!�,�}�bsg��V��ā������PpZ�c�&v
�P�c�{{�� ������$�{0�k�Y�/�jq�U[�z�@�gc�MMV��oF?�/-�����g82ZTl<�lU�֎-�~V����^ɂ^g�ǱD���G��\q�!(�0�k�3?F�NI`����@�,C��w�y�\�� ��NP����IcKW�d������v��IE�C���c����|kG����D&�Y-~Da���;�F9���wޡ�ާ�GHJ5��+�H��1�#_�׋�^����X� ��-F@��C}��PU��Zy�#���!6^/]㖰Ԋ�Ѐ ����[r�8��J��#.X]r{6�R�`j��p$�M�

ji^�WA��_�K��復iR��������X]0��Xj����G�0Dy�D�79����W��x,Rȸ����A�!�W �x��kDd&����Җƙ�K�4��.��������,Y�+	�ʗ��wDA��"9�6y�r#� ��Р��k~Q^�ܸ��T~=��Og�"آ��Rdb����1�D�k��էE�쫨q�kdu\=1���$��}�u�!���&�ȑ����B���`u=���aS��v�N ��k��;4T`�qTarn7����q0�7�6�Ĵ���Q���L�?Ϳ}w?V0�����H�Q��BF4�ı�4KS���1�;N�?�؂ �P�l8%�$���꜆8ި�O~A#�p6���t�ߎc����0�l��	�������GN�j(g��Jop\�$�pu^�ad�#��<jT��b��2���//���ɲ�k��ۭa*n�]�l?	A��I�=~���@KZ�:���ʂm3q���گp��'l��{ѱmp��hC�xO�Aw�Wn���OS�%��L2��QИ_�V�8��֛Ԯ�����͎c�r��60r���CUpF�}�r���)F�v��� :]5�A���a¿R,A�xG���?�af�7Y��A��͚����y+e �"���V�R{���^M��c^X�ƔC'��m�6���>![�����^��>�Y��U�g{�-[Ek��6բ�]qb���VK���5�u��`��(j�9Zß��yԉ��l�+�+\�dn��,E���v	�wQ�����Mf����=��yل�M�~ɯǌ���|����q$ ����;;K�j0��&}��d���h�nZ0/!�K���l�b��� �� t�ΦBH� i��i���΅o1'b���|\À&}�����E}��]���zikvk~Ct)}͒F�)G�/	�NqvI���_�?.�_e'�+f"��A?���A�Sǋ�q���s�:tt5s��@�XZA��(4h?��p�*�?bE_����,��	P������f��q9�%Q���N]%[~��,�����zV#^���*c��I[��
�UM%&M1662J~��Zwm*_Uu,|Z�Z�w�b,��ވѠ��������^�ooI� �q�o٥���m92��2�+?���!�������]�I1���1�:��۔\�7�E����fyk���>d
���3���g��۱8��)(���#�p��t:��b���d���+N�7,ƫ��V��n�q���Ah$-�%�H
KJ��n����J-���4��}��ۆZ���q��Cy+<�
�ô�G��X.ؼ�qȟ�ǧ��h�1(+�����{�7
RnЄ[i����p�e���Eᡁ��䤜�L��R*�g�~9#H%i��<��H����Oy)����.ȵtx|/�T�`:v)m�>xt*��=��,[�J纘OO�l+�Gn�1�l�����!8�ܾ��(��z��;m�]�A3qX��΁w��}�/U�+�:��k5)�r�9J[vxK�Tf��ڬ; T�%2J�U�K~��y�����%�����<�d�Ǒ 'P>�����2��2�/lf�I4k�Zx-7@ԁӊc���t��M�c�\������U�������z�HnP�^�����?OH�cN[1���Ꭶq��x�E�[��Jl\���7�oC#��I�q}bp��G�H/`��~��s���[;_Y�[|r��늌��
W'YY�m^�t���
GX��q��5;�\�k)�cI�P<_t��D3%���!E�0����K������7�%��j �o�AM !=�v���9�ml���yaKC01�B��g�U\�V���}ܨ=���?Ւ��"4F�����{�~x��S�Vr�w�_Ä���U����P�bZf����zNz%_��
+�J��9äZRIx�٠y �481�ya�����+a�O/4���b1(*A�R#���N�o�&��^I�a����5%�5���]�+!<E�7�D{��ǻ ���D:�:w��y*�IJ�P���/�J�of�uTysӜ�*��Q� Gr��m~\i�6}dd]�*�PE�>�+�0����@t��f���`�u�$h*��Z���C5�i-u��H�$aP
R��z��O�+�O���s�q��g4&@�0�=9����[�����>��أYa�C���%����#l�~�Q۞nƏ�+'��غNS��~�z�=k���C ���+J!�Ge%�ˢ�<H���9_.�����զ�<��pq�*7`��Vg~���$����͚���$� k�. ��b#Y��&T~������h7?_\�(w�gI��[��1�`��᮪5�8`nh���������Y!<`R�5p)ƛǼ��]]pCC�ƋC%]A��nK)
L1�����恩#�܈H��\��,�"�ޤ7o��W��XZ�#!�8cjЬ�Y�G��{�/��h�Q:	F�f޸�V�/�y��#� ����̹P�S΂�����Kk8{�5W_�1���Y����8e�OI�ʓ�e>�%��/�&�z�H'�B_��')����V]�DO����"DĨST��e��yF}�#�8 DKfo-	���Dz)�c�/,�������з�+�S�%��?v�w{��zF��u��;H�際���:�Cɚ�h��g�D�xs�V\#�ؘ���L�4G`F�y�3�������C����6�&"oq'z*n&S��U𞮤�c�Ct�K~=b�A˚��zL���ʳv��b�}/���9�po�H�[�{r8.�9���CI�\���b�w�w� io��`P������ݭ��0+�cp|�T�j��BZ)~ )�;ʪ�m.nG�8�ٰ�!	V�X �vaY���!唐eb��~Q���]A��F�97 ڧ��uG�om<�g�!�l��-��?]]-Tm��2"ⰲ�ޠh��{���iY�m��Z����ǭ���ѣE�ʤ���t��b�{���p�`T��yZm�Ĭ=2%a���#������X�B�����J�;���I��P�D�Ņ�(H#�N|�}�#�.j�ك	��9�hj�ܶ2(U�{�;��v���K��v�ωI�$xnӗ���n/��̣N�KLL�&�U2���i֥��gB�8*у�d��"��Mu�U��M�tgl�i�bGnU��{�ϐ�`G/��OS�g�u0:·���i8�F@�Ԗ�u�h�o�-w�b�Ta2W�H�Ѥ���D��!�FZj�z&�F��W��X��������0?aƲ�q�	�'JԒ��D"��X�fOt`f1z����JN���.'7&�9Qv�$Y�'u��"�� ��ʨg���#�#j�R��������q�?�X��6�<]V�g����:5Q� HL�/q�Z����N��,`���Q���Z�^��r�#"%$��:����1?J*��f�R@��ۉ�(�:�:acǒ'P��*R�S���l\F��9h�1�
���	����>X��,$@� �T�չm���E��j|R�(-z%%)���>M=���.��Ⱥ�,�Z��f �הi�|B����C�WcӪbr��{��E�Ѿ4�(r�`?OHB��hč)��V�M����N�#�m���s�p�NW��.�Ԓ�{��X5��dd������P�!L6xo�� �����źp�RE{�3��o"��"�����z����%W���h�����Ļ����Q!�J��Bml���(8VMX��m��[6�*���G�qAz��T�M�����>4�h�(�>~B��K�?+xԥߛ�'���b!���8߽�ь���^~�B�ui$Yv!:��ϻy�	p���ܼH]�v5��lg�.�o����H�E{�"3ʺ��C)���^$pa��9&��S��觕�!�6�(��$�mjB�Ơm��k�P>w3��a��z٫���Tg���ؕw�G�p#��\�"�x��2Ǎ����w��7D���<U��4��2|k����u�mj����Ft�J�-����{K���I�%,ے,��4 �WX���%!<�b:)5��`^g�d,g�:0\>	_�Z�͡넡�EM�X���4�0�Q�M,��v0�@�ۈf�=��t��� �|�.s�!�s�u�G��)���bFu*�}��o��ohAW����0�~N��b T�]sy��IOdJ��;\�)�b�U_Ζp(K�������~�I2�L-C�hDu5k=�W@����G�O�[>��II�VR��F	ܨM=9C?�R��&Y#� �T1J#��JӸ�p��MQ.����9H�7��7�afM7^<�j�>0�%���"
}�Ӗ^L���`��"��ĵ�m&ǵ���W+��y�7?�K�]�u�f��S�w)6�l�p�A�(�lR���J�+^�-�]��)zkN�阋�L����!	,�-�S0rY;�D~!?=���L���B����A&����� ����a���E
B�ޡ��m/�4�N�V��Z�9���#��W���^2�'&_����H[�
��p ���R�k&����4Wn�BU)�5eU��.+m��#�v^�2)�)^�>+@J�}Ž%��T��X��.�a�M,k�o:E7o��,��M���]���2�>�fK\p����z`k71�ҙ{)i���M��m蘐/;:(1l5��D�=@Fo�sH�Q���ۣ1�P+���zX!�� X?�H��!�,��GֆU�n,+e>V-�İw�h�e2�!���Ȫ��#�7����9�{t1��S!^1<$k���⃈���m+I7��3�8,�MS"�O�hy�������@�u�x�+*j�	Y���-h�U-PMR�L�M4�k�!ʼ���B��3�3Aǟa��NT+�M��k��A6�J������f�/LA��W��zG��^/W4�CH��u��ְ�#x�F�z6!����W����?<4lL3g�ʾ�C����k�qF�������z�q���M�\�;���@}踐t䋭���g�������Z���ZYZ�38�PC"�0�8-dn$O��3� E\&gL��+��'�?��M�6�?|󬺍)o�|�X9^,�N[xB�T�����CūT/R]���c��k|˘��Q�&9���Fd�l�؜S^�k9�
��3�a��H'Ȭ	#w�	���V�=Xx�!�}O���&mq�$�8��4 u=5�4Nۙ�xo��}ٍ|?��V����_[{*}S��!5�
�h���x$b�0�<]�\㭫�Dڨ���,c�q`b�
��5ęe���jN�5�Y�a�ޢ���:�#�4o�ȅ�x�ٰ%�� ��(KݢyIR�B�"/�����Ξj���� �\u,�(G�vn��6'��^>��/�z�94oMYA_�$7�h4$�9��ʸ�و��O�ksW�/���Y�pV�ΐ�Ju�t��;�A��GKF<^���տ�����S[a}������x�8/ds��o�Д�M��H�	��T��ю��Q�6n��'�9�/71lhޛU�"���8�=u:sB��)w*�^��v\�9�����C.�Z��ϒ+=tmk$T��OE�C���ՙ=�D�-L��Kd�C�j�gT�k��E!����Q����ؖ�����9嬙�7��J��Ew�܋��<�	�M���e�>{ٲ�d��l`h���&��;P�o�ܛ<o���N0�:��.�з�ZлQ�bG�mȝ�(�����i�JA�S��'�2�̿o�N�\�ȨsH3��.�机��gݣ�7k�o���\Ϥ���H�F8��)<~�k�ٝ ���="\���g��O�Բ����a�>��$�U��z&,X�X��Mr�~4s {uK���R��r���M���q�҇N�PY�wп�XQ9���A�oEJ�ϸ�w 4��<�T�)�:��e?C�r�u5��QW�kHP�H�]gt�<�*��׬�d!�c�B�<�<��,>MMX����&aC�S�Sa���iS�z#�"&|(Wr-E2K����|yN;c5.�F��ݹI�d���UU������N��V�m��گd��Z�c�U�T��9c6~r0쮋R-�rK�R1b"J$r#�ajS�ϒLM㦭��=�_Wb���~^�c���ಉ�+4�U��N��im�y6�F&���6�?5�Ho� ��2�����N8�|a?�6��4}�����-�"|~�:v���r��y�}H\B��N�ԓr�@6
j�ϫ���A���:8P�Q��]�� �O�Y��@�������i����2��@R%�]�ߩ�$���^��Q<�p��3�h@I��]!F�AA���JL+�ɂn����B�������| -�s��ꢨ��H�+�tZ��4{�N�����>�TP��=��Qcs�&���,�CȠD<u��9�\�⦦���<#g�[}�Ia�L�4�!
�b3�3��tԔZ�f����v{��(��C]�+ ��,����Z6�K�Y�
8m9�u_Z��G%U�!�&	I�+ �FC/��6���~3�wޅ2-,��>�7𩲍S/�H��`����t�7p�M`�v2��Q�e�s��'^L'�͈g[ԧt�h�H�����d)�â�����������w�eO���m��y2��S�Ω���&�)��)"�Mr�����_Wd\��5��د�L�����q)�_/���ޱ�6�l� �*�G�+w��� 5�N/�'p�lZ�#X�**�B<<�X�͇T���4P�����]<#����|��RO h�urm��/���x^��^q(خ�g�k�Y������=�{��!��-_,�r$|ۣ��C��<Ύa����+#J����˦Ȯ�i�oj^&� �|��t�����Z����������E�h�F.��!����.Ǵ�;��b�ě�:��D565:2t�,�R���0�_�J��vZ�2\��~�|q}��s12|,-�dr�(X[��qb�Y	�3��J�Y>���#���T�mʱ���sw?��j�=�rg�v0UTu�~o�^kk5?�� �=f�Ib�2�P�?zK�$6�\�5_8m@U}�]9�%Ҏ�E ��4J��Ҝ^��[�)$y'����d=��p��p�Ѕ�1��t�cI{R�r����J�f�#��LB�1ڔ��Y�[�}=;)����*�m�N�������P"8��`�G�f
��4v"M�歵��h��35��=G�G{��#��y��p�68ᗘ��JeGFQ����P2�C��W�c����;#�0lnUh��g��z[ObT�������lp�����oA�6�Ľ�UGZ��LN�g}^s��� �aieԕ��>X������bߑ�nH���H*��V��yc����������L�n�7,�auLļ��")�b��$�fr���)�j/ �gj���7b�1\�y�9MpToP�_�Q�7d��1�
[#�a���`Ë����RϬ^��+���7��:i�mꂇ+cM�P���+Mq7(���'3�0�����D���x}���^�Ŗ4�6�\�9/O�ǹ	��>�5Q�|�&5�UJ���-���61����5����@,ɟ��r�;N4�Q���Dc)��vl�̲P���7���� �c5��r��]���!IW�曶'">�r���|dD��Ƚ_iHMM�_���(輎ᙑ+o�#؎�%���;�	CA͖W����Z�.o���
�p���2`�B�)W����;��<��ĹH���`�'�@�4�c�@���B���̻<1����A�fu��ޓ��GFT����Az�g���rg��Y-{�b�8����� d:[��9Ӱ��X�Hn����Rz.kZM�D镕^II*H�,{!�ȧ�\�nVI|_�J�_������t(�au�H��XST �
�[f��������!ײڑ	��C\���<?o-?���U��!���r��� c~�$��Ǌ��{1À�"�,S�"f�`��c&~��17>˃{}�=c�Ke<�)Җ�xɤ�=va.�dQE<f����]�
-C�=�����%�m�]�s;k����Lwj/�f\��R�l��/�&e��Z+�Z������Jm��P����<���c=����8gZ���1��p�W��� ����
ǵ�������l�0� "���~��N#ެ�л�d?0����Ee.`��Ǡ��׻�7�l_3��VBv\���s����i)���FM��<�c�������IX�O%ԑR}���y�u��j��C͛}ֿ�Bi�R��򁕚�����}{(����m�b�n���׃��]���:]��nO��5��&BLl�H�(�;�^��o&��x��.����O~�o|��Y޻�]4����W�!� CCY��9Y*z����В�5�H��Zd���	�?�r�إ��"�l�
]�����TG}�~�i�=�
e[@@i}��A'�W�&�L�D�w�h~ S��K)��e3�WX|��QvD@M��[�j��H&ODR�+�E-��)�]{�#Ò�Y��lA�%�HϜ�_� U�1̓�����@�e2���h�n��G��B ʋ��cW�6�[R%KӐ.�?|wH��d�{�W<|��N��*
��@��y�L{#�)���d��/ �'W1���X�� ����|�A����������}��vK��;69O��s�����F%[^�G	[���A&*����A�>����eҀ�GQ]{��������� ����?�\�Bt5��� �q�uپ��g���Ԭz?Z���2}%�R��sKω���]jMg�o%N9t�aP��R����b�9��Ȍ1nql9,D�E�6�ֆ�c�5��S�'�v5颇h��%�}/�b�׏���������}�bwl�o]������{�!�Q#�H�7c-����� �e�*��Ɇ��3t�v�{�N����8s�)���_;Iƴ��N��t�;'�ɪ�.�t�N;�C�z@�~��;S���!�� !�(���� S�y��Tw�Q�O���ri6  X�H�3ԑc	[�T?�=L��*�?�k�O]�ĂO�k�S3N�:��{���U�4]��\{@���h?�`���#Xϸ���إo�t4����
t�OĻ���Cl�	�M@:�U�i}cC:��+k�9)�AW7Z�_N��:k����Rq�dA�kR�]N�k�˾�	��ڤ������00�K��h��]k��nep&��N��:�iX��ב�g�<~D%�r��Tl�S3�p�8lF��P�e�����1JKxG__�����b,�έ
�f/��bi֣��"�&wQ'�n'�T<$<5�\HlL��h�AQsQ?��\��v<A��R5���#�D��a�L���U��뤈���|��b�.��������Y߃���ۃ�?w2��F��+xN�h^暚���YV OK�^U���~�N21�����D'x|c=3����C�|c�4.%R4 f�©���9�b�}RZ�Z��� �_��d1Jx�m�����;Fsr[�s}��'=�B��Q��۝����9�Y|
|NӰ=�h;�$V7܆��L�<�>]ҕ�����/%m�w;"��т�>q;t�c[!��E[�)�ʸ�Q�@��$�ϟMq�q�ʛ(NKŤz_u%�q�ʧ4.!���/:��Ik�r�3��pI~y�d2��
���X [������JF�ظ" �^Bo�c̈�g����	WQ���B݌z�"�]xkYr7����cFkB:1x�~�$H����[Q9n�h�#y>j��q���a��ޙI��ğEua'�zm��Ad���I���^���)r���3�n��f+	~{�ُQ�����4o2ޱ��H���}����:E�`���mͳ������sQk�L��U���p��i){��T ��M}����۲*���J���aܭ�'pl�"`�k@��Ai8G��LIt��B{/��6�n�G?c��7MZxY��ª�{��F^:�4���m�pdKN�s����x.�F�n� t��Dq�i+�0��]�]٘��d����2p�c=XQ�4=S���3:�JX!�K�,���	�qs'�����Ͽ֡���*�d�b�*��E��c������'�]�r�-��|�K�И�U��O�q�]L�q�%�'�t��?_�0�M��>��i�O�R�<!a���"0�1�� �X�_��� }�����~��R��&�V����{�Ε�K�fEX5˜+k�������	I?����bH��n���cq�'�f3_��`���?�4燅}��%G̎�?}K(�X |`�������Z��l����?��܇#�ɷ�� ��D���un>Ud3rxh
�JgNt�&?�r���H��ۅi;��As�=���%�Ӭ^�3��<��ڂ�<�ᾱ��~��퇄���j4�r�52~Mt[�Of�)��/u��p��hhO2����Jph�$Tn%��@���1G�@{$d�A���ȇ�yb���|���3��g��r(AO���?ɤw|(?�F` f��o{�����Т>B��%3��?\�����!�̟2a�<s�ܕ�.O6")�߅Q���P^�<������c�w��Ks5�m�4�NHg���C�\C���ʢ��&E��3��i2��=<χU�����I���.|̰Y�n��Y� �� ��B*u�W^�#��%q5�]�̑�KR�����Z��%��&�d:`��j�ق�G�� J"O�z�6���k/)��~��)��@Ѣ�Og�*�G;�CTM+(��ë��A�gX�(#�!΂�����E%�9_�|c#��B �Y)�K�VZ 5��.�|�CZ;@����o��c�	w��($�t_�w�`�89Zv�S�ݬL�Ö0� �5O��G����/`5q{S`��	f�汌1����e~��ު xV&�F���͏is��O/Qu��$x��/���z# �M4J~9��[�%�~iœ�@ ���b��l�WP�:Z.������<�8.B�]�^�Ʒpg� ��&����
�9ϺC�O�w�Z�4���ew���W�6�. a܋�1f��x�A�'�Q�#ko��R� $e; a���<�
&��QSL��j�����8%uZ�f���%+ߨ�gokEhM
ܙʃ�ҫ���F�Z@k�qӶ�8nS�[C��9
�o.}
��&9#�^w��i<P�^�46_} �C���O���K��\ҽ~�m�H��<*���HQj6\Vm�U�E�K3�ұ7���k� ӂ�H�]P�?�)��&t���]�b��CT�+�P�����f�p��c�,��P����['�?'����y��p�k|�`�xL��L�)�����ٓL�A�R9GN���	�L��[n��*[��kt].�{��F@��{�/+���5���ת�I��ʫe��K|��$�}cD�E`΍���Ǖ
�����]4��PN
�u+I�4>G��;��o��J�c�f|�7�pPd4��5ֺ�Ə�nh��>t=X<�g�|���i��
�Q�X�lrF�/�����K��a�'��7_#���=�$>�#��ڍ��A$�^�R㔪�d8/��M�
u|��I唈���hN�C��Dr�c��5A��c��g'a;%���+���"���K�J(z�uf>�l�jX�V�=XI �Nǐ\1w�S�OT١x�M1���C��u��Jv�=6aY��ͯ�&*�L��/ajaٗ��H*E0���P}#I+ӷ��Vr�+��g�V�@�������v�����[w�׹X�������~���b�Z�8��q�G�����4�v~i͇�ȅ��e[��D��?�Ӡ'LTT�æ�����Ǒ���Yn��խp����c4;=�｣�~n��t]6���^ΝQ}�ߙl)��H˅%����C�z�b�=��V=����X��Ċ!U�ޅ�q���|x�����xh"���G@W��	!\!�˲�τC;:�G�d��
̞FG/ߓ�L�UC,��8^ј���� ���A�^��'�'(
��m2����R���r��+!��6l�s�����I.���GW��y�*��fu [y&G�ɟ
G����&j��j�0�2-1�S:Q2��!�P:�K�(�m�n��sE�D+L�B0i�Ȯ�]n�tW��2���0�r�Ûcx�&M�{r ��"�j�����P���8�x)fhcѬ"���#"�R�~�>455��ﷆG�/����:���q�Q�����VW�:Zt֍�/@6z���[����U�pI9�Qv��R�5��=<���@)�6ժ�y ���������>#�ͭ��R��mΐK�jA�a3��O�D|�V1��U�jT���i�S��?kMq����%G�c�<zJ돠A�sE�N��G�6�2bd���n��(�=u*��Y���o8����fI�bNz�z'Gh1>n�,�C't��?i������1�vX}4"���^�Q}/;^v���q9s�~=Kl-��x�6��:���WZ�o�+5�d!��AH��;�L`!k�4h��9�_�7���b`����0��a]z���ot��.d! ��Nc`aD;�$!�bZ0@�q����q�����/ift"��><���1/`8�jXj<��vע�xk��Bk�7`�𾏊s+�8�|{Ǥu����G���u�ϩ�9"3�[�*�oa3�1�r���Z����S���T�X�y���]m2)��j�o�go�!�Ό����}��t
���}�0��r�l�m�گ���wu�@ w\I�S�~��� q�� J.ݔP���,�@X��v1����ؤ׺3U�E�rچd6������A����,s��k��.�Ae����xW�V8舶׿�l�������k8ş�����<���O��	�J*�c.& m�IK��'>�>zs�����,���PV�M`>�v����o�� ��>,��患^��{	>k+>��zX��q#�A�%j4�j��[�\`�dS���#���O�ă��)?Ӌ� /60��{sY˰�՜Bx�0oC�����D0Z
%k�%�CL��I1�*X��'�o���q��SF�2%��3��K�֎#̌��Z�A(`�0�$�ڋ���7ˍLQ��O1��-C3�؞�W�T�3\ԓkS��*��xs]��-��rY&�Y���|���(��9߶W���ԝo�nɲΎ7&5,�\���29�,��c�����}uHt�'�d��b�8�	�L�a���:�LG�|�T!�L׮�_���¼�w�;/n��=�>��}V6,�0qr�)������˄�0�dd�S��f�F?��k�77�)3�[�9���\oO���X�#Ћ��[@}�ԝ�p�G���o,j�*��a��`@�Y�����cR��}�Z�?.R~�*Ψ�9��񑸠7�fI�b�2��_H�"Kߥۆ�k�|u��a�@����Oa�x�G�����ﾣ"��m��C;�n���XGѸ�i0��"{<'�VF�~u�N`b`��#~}�	��[r4"&������iT���H]6�p2���u�_�9�Z�'���=���F��t�E^D����k0P)����=|^�P��������t���3��9��X�k_G��`�`�U��J����o��Ӏu�ʀU��w�et�O00�
�OJՔ�^����9�ˆ�W�,f_P��j�Ԧ���]��H� �eyޝE[�Ҳ�&�8ܲ���.e���X%��̺��`9Y1T>�.���]���#N�c_>��8���>y�U�+��U:�H�۳*`��I�WFW�ȽB��O������n�q�1=|^JT��
7A��j��',LC,�F�繭�ϵ��٠���R�F��ѲU*+�e��
2��zk��9O�'A,�_.U*�����-L����O/���\i�>��'�6�G�?[���Q��Ql�C����lT[w��kJ�i���/�dds����O��x�N���J���Ȁ�*>��i`�|�.&�G->���Z:c�@�C�O��\������GfW��>j9n�btZS�pّk���Ҡ.70�[N@�$��3&�8mH�Nh�P�0��?Qp;Aj��B1�QH�\ܳ�2�<���=����)���jޣ��<��o�dX���3�W�V�z�7�8��Q�\g4��w��ѷ����H�����lCji�q���B[���1<F�
c�
T�G%����w趗�=ӫe����)���]z���ͨ��Q���P�5>����J���5	��Ӑi�8\�{�Ǣs�.דđޓ�JҌ-�穻��9��H�wo��]XPG68��;uC����ew[]) ����i%DY󹣂Ab�V�=��;�֤����H�Q���7A;�����:�>#k��ў�Ϫ����Mx�d�#Ba�4�Ƨ��VK�����������ʹ�Y�$��ۨ����.��j?������;������h�}g��V�5���B��s��q�������Y�p��\^�(�����)�
�L�1ȠuǬb}�+fb4�BQ��������G�C]���$RS,�,��k�J�RJ\�@��#{5����j[����/9	���%��i�������{{�K�tցʫA��݄��}���H�mk�EQ�k���s�S�L�ő�K�V�ߦf�MIC��F�$��v�ğ:+�%0�NT,3MjA�����虶�q��S�h��²�9?^�`�)G�@�M`�;r��\�h"�A�߯ @�;��M4��oy�<�=a��Jު�W��U�l�=ݲ��_����z�c���#�� 誜�j/B��z�=�W�؎OYR�����`K	f��Jq/�:�Ȕ�ϳt�����a/��d����,K/��eʮ�Z� �ևZэ:�^�lH�N,�^
�==�|��F0w�=:g�]]c�T�����+*k��b�����2 �U�tb���zx ��q�`��,�=k [����!Qk�4|K%���5�^�2i�G�U����_�I]I��r��(جd�n�&N�JU� �N!{D�?���[�� ��%��B:��>2�Cﮉœ�K�i026X�I�U�R���]\w�j�1����h��c�����'W�h�J���IC1�t7۔�to�R�M�?���T���dĤX���	<h�h���e��5�aF���I���i;�Z\)�E�*t�w���<���
[�	D�$^1��W�u��D���q�f�"���D`f�#zuE�����Z��-Z ��B��/��\�9�C��VOǕ;V���;ؔ����Fb9%����`uy��Fߵ�CZ!w�{Ƅ�o{d�[�j�:ڎd��?��{�쯷�T�*t��I�eE��]k+~��>��X�ԧ5y�nSM}B��B�T2��_�]$�d��]O>�j���Ċq�X�\�����h���8X�w�@1733�6�DC��xf���-�&`� Z-I��,0��K�8��7Uֵ\�>v 	�\}iE�p���X���Sق7*؎����'j5�SF��	|P^�8%��L��M��J����Q�w�=Uw�f��P�k/if
�@�5qӄ��rc9�9���ҬK����r�M��}��p?�?�3��;����D���N��}�>���~Ҋ��	ږ���:� Cз�o��4���E�|@>bG�D�p�W�[���{L���;�C1��<�=�GE]W�؝=��z�=ڇ4�U�v�1�R��s�a�y�9��V�����!Ё:݃�j�*��#�m��}L���.gtS��,\�]�BOk-��,0ɘ�P��ȃCʳ��M��}�r�u�����{;�ǻ���fY���g�_@����?��%���\1�<�i�!f���0\�%��BL�*J��8rs&���p�UB8��߶��ڽ��f��ׂ$��g׬"��j������C� ��8��ٻ�:�?ss!�C8�lyU%2�1�6lP�0�#���i��H �>�|ǣ��s�q�9��M8ɒ�D�������2S��>M�Ŝ��=1��G�Q[p�ϿA�8�@cX���b�� IEt�3UD@�qY���?,���e0
�h����`�R&(�*`'��Ɉ�[,I�ʅ9��К��Y-���2޲���$/ѽ�c����+�7n�L��NG�����ľ@7��b(ȒV�>��cC�{=�K�.�����sE�M�$툔tFm�?[����eT�.�	홱3$��i���v�3�MD�TLԨH���ў{�&yJ�W�j�K^�'�X��7�r�����º�G7����&T]AU7��+a���^C��/�!ɗ��"�cL6��<N��5��&/KQ��	�0DtXG=œ7{�N,nZ�� �����ͺ����X��U
���Ӛi���^�#�K���%3u����U6��� �(eWiU�D,PQ�u�ޟ�g����e��0"~�����o�(niNK���|Ma��,n����{�1X72��T��[V��b�IJ�;����U���O\;גK�R�#\P��z�0���	cGP��!*^�<�iy��x��!�O!FK$	���"#���j �,�m��O�g2�\�XL� �����2C�wOrq�b?�%�)7�c]M�)V��/@~�����=1�+9�<j'WC�mx�/|n��B�}�[�)��?O����*^�}ŨN>o�j�)�0�#��e�!P�}0^d��7�C)O��2K���}`���Z��2┗Օ���=�2XZ��J�ڀ�
�>�]-Z��>ڽfA`�(��]�M�<�`��"��/NcN�Y�J+��k��q�`)�1��݇T��ļL�8c����
�v^����ZXʆ��FP68�����x�X���f���a����eR�^6�)8���I=x��� Օ �P`B�*b�&e{��z��	����5�ځ�*�oF�e� ղA}�ʇP�|듌�!lФ������N��>�Of(&L���j{DG���[|d�%����=4�a�6��ya�Ё�->_	�d�uZ<wK¶���^�GK�U: o����m5�x���P��T�!#��h�v����Ty���ϧ������ V���/�&�BV>q�]�U^��<h��fD�� è��҃�M��=߀]5�/�1ƩZhw%)I�zL�@hnXSS��e �vf�|��>�@�p%�C��̴`�u��~���F����
�h����?ոn뺳�Hg���8�jd��`<,�/�W���J��� ���L;�P��8z�D
^��S�yhN�Dhq)����|��S+��BC��^��(ɕ����sei�Ą(����ƀ)�ZmV0�pq�u�Pt
�'�GE��p�_x�+}���3it��y�����k�P��7K�yɾ:����͞�ȶ㗂fU]ܘ�_�`�H>�×dP��@y��onFg9���Cg�tϕ؂2�c�)���	P����9��p�$�W�D��D[�g���o7L��NR�g��Q�W�	}�����2*p�ư'#�T挕�HJs��m0�]Ni��^i�+lױ�Ԏ���	yԃ��n�~�J�n���}莐��{_�v�;Yq�E��Z�Xp{�>^k��)ڲ�eGڢ�i����f9Mm������Qd�7���]f�9Ul��H��!���t���r+�ߠP^��G�p�����MY|Kbȝ��s{���T%����Ǡ��o�J�$
�ؒ%ʑ��0�Q�ha/�d�,f��&�V�!���t����\���X�W��Ee>�k��p��Ue}ˇ1H����8�Y<����#Ў^QcL�k�=��L4lv�FR���y0&���h�a{ ���r��)S�-����okC-ё�RB�s��Kx}&7����#���2Ƭ��ae/��+{N�0v�eV�y��k�A��`��^	��W耷�5@��t0L�r�zt��ԏ1Qp��ͳ Su"����;1x��!-���q�B�+/L�>���j����ɑ�C������_6f�\��a	ګ3�t2��
M���>H���$p%������,�Eq:Πa9j���kY��,>)��\�i��f���0謟&6�'�n�)�$2M�p`c�Y�L��=hZ�M 9�cf��S5���d�����3�T�w��9'�\�b�0�gB-kwϒ�Z/�m��"���*��P��z�_.gE�����P��ԖN�<�Q���k{hh��G��Eȷ<�M��9���啞��'u��d�l�����&z6�[9�`7���_�k���͇�-�t>��,�b��
��E����8��5��%�R��cq����Q5;frD���s]�T1v6 �S�]k%�U��A��x�@��|tjw�Aɂ� ��$j�1mC���&���{�c��	�y{=�E������$H��	3uXH�7�l�f�i��1f����>5x�:5!��4�i~ ��x���ӑٶ�y5)�GƐ('�^��L��g4���@��^;n0�L��`+���U���7��DO�0��0�7Ɋ�&����c����!��8��{�X����}9`���������>`��[)]DTҗ�m�Q%���.u=�o�U��bm3����O���p�JFA�F'R��xQb�:Js�糀�w1)^��NBj􋯑-�b�
�p%�-ǒ39�,p"����c����y��O-`��SR���+�٦�{#�i1K��MB&ޅ󑂦*����Ϛ�va�$K���h23ip#��U��3�����]���	ڮ�DQ�TO<��瓫w��X50-m��pN�?�ǎ�ĵ-{�b�
��;��6����o��DE�A,j���EO�͙�:�xP�'���%�b<�p���$�Y�6*&uF��2���v�=�G��V7���T�\���+�3p2al����M-�;�a��\�bE�dC��Oq�����0��c3|�[i��|��I4d�h��o�XMk����m<w�L�~��y_�C��Q�@�GFn��0_>Mo�ӎM�	�
��iz���nҌI�U�Կ����ϲ�6OUY�s�w��v1�H3�n*򚎹�V+�X�R����T�g�׬�P���*|ueH[�om��/� ,��N�\\�xP6%/9����O��#���}}�ԝ��&\4�ə+U�'� J���X��E�r�x��7K*�����{tI<����,��,RO*�*~"a�3�{5���@T�ZV�2S��+��J��/Uc�%�۱SA�OUrs�k�Y��s���G�55�T,F�ep�4)b�_�D�wgF��1q����!W�W��+�q�6�e��A)�B�ůl�f����`}k��tߑ��H3q1W(��Ns�Ut۫�2Z��C�����gL��,�`)����$�iɠ��&	S��ty~���$���C㢬���E�F4aH�#��P֓U���E+y\tu�O�qI Gv��B��{���|=�f eh��S�n9���&%N������(�T���m�`���Eϑ�F��亮~8I�p���� �g��ra�J`�=��!�?�l.T��,����9�S�»	��ȡђ��%ܗ��/�"��ލ=�<
)������u��l���A��:�* ���U)�U��;8��S�c�i�xWF�*;�%��3�K�>N���8�p�t��O_���u>��5a�we�WM��3@�(r�uޓ��`h>a��X��靨G�����t[���5N�{i��@/p�9���9L�ϙ���A�U�t��S��!��-\&���j����)��O��������޳��U�UO88r4��4�-"]݈0��8����|�5��J����>5(H��f^#�3�u���H��'�h�HR���.���'1dl��`e2r��<
R�wi-��9�*]����dcqH;6ʡ]`9מ��M~��-��qs�x]�Ϡ"�r���Lo�!Cq[�J-�� 0!�t�
������ɡ������,��Z<�0wt��p���R�����>�,ͽ���[�:����L�o2��^��ǥ}�󏈴��9R��`bu V�f���T�������Y�g>A�I!�w�"������)Ҏœ�eH> Y=48�͡$�������>: ��y/��3ה@���Ծ��%����j8(�1Α��p݊W���λ4h�̮tb��Pp��.�Y��v�|K���Y�j�\7�.V��9W������J�w���'�*Uz�8S,����p�0V�T��>���z��?Q��=��k6fP��t�	�r����fWr%c=���x�C|[�I�F/4�z���;0�� }�`��c���ș��p����`[.�y.���=��y�Y&������'�j��>�M�AX��[�qf�g7��Oz�t�;"OB���]A�Sd30lK��zD_�%�n�
,�W��~?L/U$��P�?�R{���ҙ��QZ;��	Kf'U:�`��?˷�xp�&�"����8�7��kV<0���Fq��L��@�X��g���J%_��o��|�W=�3hE�A{����L���6�as��y�>�O����$�6J��pa_���F�q��>22�ТRb�s���C�Ԟ,=���q�eu����%ߖ�sFO<S�P�U��]:㔐���P% s�������3%�����!-M��@�,�1<d�Hw��n���\��7������d	��+/�mK(no�W�u��k�%�{��E��+�0Ƕ��"N�8$t�)<�r%լ�� ��#+�o��ShT����Oԟ��*�v�������GA�lb�k��d�a�o���M��Xs�����7T�� �����5.11g�yg�9���3x�\[�J�ʨjKC>��KX9���.�o�YgG�"���{��K�;�vA����Y��4��c�s4����x0j�9���o���hr�Ccn,*�P�~\�W1M(g���՘�G�c^{a�Fh���mTB�����p(��K����˦���S����
\p6/�� �ƐUN0bmW�#��Z���m��o%@��t�Q@����@�ĤqJ��޵��tr���]��u��a���p��`�+�j[���6��
��vkB�G�Ht/zs��H��^:����s3��|�G'�W��v�Qnq��X�/	�+f�Z [�ᦎ!0������H�� |�B4����ry�������t�C�X��g���H�� � nK�[/� �NW»#=��0#0�E�
]�tT�����=�G�l��ₛ(�(k3��k�Q��$�����/��Q�
z�Z	Ms�x�W�1����V\��Km�"P[$���'�G�2�.T�,2����/�g�P�ʱ �i��,���^o[O�%�<�}̄�����-��w8w�r/:/�v��#��Fx;k�Ʈ]ѥ��'�-���G�%�#?Q����IlM<Lַz�B��l�����A�!]���(��{ɥSg以�>_d?�j<�u�Ҟ��S"��8����&_0�:�� ���l��O�H����#���X���R����A9�ҁ��B����x���fʂ��LU(��yc6�2���k��ġ�'�=�2����V��Y��S��ߩI��b!^���<��7���X�߭�0FC���n��i��@���� �3/�"��Q#n��w>��琾��f�-Y���������M��m�>}�1�c��T��0���S��� !��&�"��f���Mu�m�>�qA�	�͋�L�%��?��2m�yX���gkjJ/	ʡ�)�6淞r`�܀�w��]9�ۈ?�A[�2cgBc��a���+��&�)�
E];z��A�̑���d��k^�^��أz}�UٓA��^��/�Fh|��D��ex�Q�ӱ����{�n2 ���ޫ��~ ��Y ��� �y �
��{>�5������iwIH�]"�{Mϴ�����]I�@�N*��O��j�����>/?�`#����('�!�1�v���/t�j?�HȀ�Q(�Qe��d�"F�b�
d�ov�uu=�#�p���62��P�ϡL!�i�:�d�e 	N����S��|��^'x��Z����QyE��r�\^ZŅ�`�����.���P�����l|YDj� @)�O�� <X���/p�R���n������$>m��9��R����ڈ�eh{(@���䇓���Sy�x�Te��@T�n��	m��ǡ��E�P-��lqGR�T��E��Kq	�ÚeK|�Δ�P��~L���o����S����&�<���N��6�}��!�Hy�ĭw3�N!u"�hC}�u�TTwW��p�
�����8y9��h�+ZSz��ꄄ�Ϗ�4/�E,�86��@��vPr�G�@�z�y�\.}h��ů,�&����'$�@Q����"��s�=w�E��|�^�y3M�H90Wm�j�?D�8}y���g�5���P,2�0���� 3}ooD��#�i�nproG''M�2�C�n�,�^ߵnjFb��&��|Ѿ3��pV�8��бk����{� Ԡl�D���j�G=�-�=��WY�e�l�۟��L�4yQ�qL�
��/��f/,�����<�$��iJmY+��X��ƊVU}�(��?r�	�(��=E7�qs��]�E�S'""�K�K��"�𾭏:��;}xG����QO!�	-�~P&뒎�F��ؗ�:����\���jUl�]�X)d ����:"_�o�%�e6SQT����X��'����O�ޣ���������o���S<�ş�L� ,V�M��j���\�6t�^�L&C������4��Q�m>��^2NȲ���fn�����s��P���ϩ{ҕD1B�R�^����RR����z���p��M�6\6g85ȻŽ��Fzk�x+
�� vC���Ln�&����D;$�R��d�3�k옷"�%xO��|�]rE8u΅Ș���ߚK���5*|�ܤ4������!fN3��36O��w�\�[��u��Vf���kj���h�=Bg&�R�r�u���[�;R����c�cg���H{Fm/��o�\8��5���E�\�[���hb1e�?g���|J�W��խ��,�N��Gp�c"R}��D��i�Y�cX� B+�Kx��7`3�2�ݎ�Bof��V2?SR���mwt�%��&E��#�O* ѾO̜���3C���p�ɷ/� �O�}z�W�1�gj��JfړS�k�`��C���s�����2��ծQd3����(^��J�Ś�&@3�X��E��ɺ�]�|���<��O�%�L���8�8z7�qs&�}�>����M�N�<ɲ(�Ô�Y`QA|��<����Y�g��A!A�ϱ��-65�$�d�Ԇ	,j�2���`�J��Pf�5�Z���F��.uG9�ۏ&w�<$®���Q������mh��@:�Q��ʤ*��O�'�szC�B�5!��h��{;"T��#�#����Q�j�-�mT���4z�����ڊ�eM�]Y+��4�<�����A7�I���1}�-�����P	�3
�H��z�І�Җ����C2�-~�][3E�W����6��e��[Ghɀzi0�Ut��Y���_	����c.��Vն_#��	��y�Rú�"�>m��\
/�)J����6k�_���^��9Z�=�) �t ���*!�a�V��es�!A�g�}u?���0~0D�z��IO���ޖo�X�f�h�i��n9�f�V�_���x��7�GZ�d�Yw��&|�p�/{����l@��9Ov�- �B��f��EFǰo��c��B c�DG��2uȽ����DhvNGv�W���3��,�X��#�T�@�8�L�W-��럊t(D�h�(s��%�s��<�ݱ��i�ԓ�]�fv5	����QMS��nrz�H�z����)F��D�u|�S⺺yP����=�Vs0�W[n�|]�JcoW����q<��*R��_�Ԕ�*��9SkI��o%�X��� ��c�i+9 Є]7;o�I�oG��_���L�;�֑T8B��ptPn��f��d��V==r~d#��N�n���pmF���Ҡ%C�w6?���>����a����)�zJ�̇����|��=�oU	�CQc����K+�I�1Ӯ�8XP�D�D��u[u�T8�~�M���)B6CS���=/��1t>e��Mߺ�"'X����J^;y��s��s�>���ڟ�z�� ��N�X�p(�$x
�7���b��^�k�ֱ�I�4 @)�/���>��8�[��BȾ���X�x &���F�����
�2�V�y\/�,�|י#Ç�����m�i�:�ɶ�j"�o��J�B�&����WAT��k_;asM�����y��dbJn{k�����$'Q�����+�פ��i8�K-�.���~b�M� �2<Z�_^5�뱀��ݫ��qȵS����mQ�B5Q= ��&C�U|�y��7�*3�>���(�S�I$��3�9c���}Z��6lM��2�c�� ��s�GG�p~���-.g�7��|}l���_d`���~s�������U���<_܂T[�o��_� U䬊��cg�]�ꊺ�^{�Ø@K�r��|�@*޿�D�^�_������a-���ܥw�����Ѫt��F�j�C�'fy��Q(y6�5&WF�0�p�α��qJ,��!p���/��n�� l�a�=% W�d�t-n��$/�Gq�NJ��0�٭��68�I��[��`O�g_iA�	�,�����1~���?�b��D�s�Q�xԇK��$+Qs��,�X��|
M�8
��֝<�-�>(;y���F�w?4���u&��Bo����l�<�4��ө!�];��W���~_����ЪNs�C^ܡ���u��bM��T�Z���<���\�W��,�� T���C��hm��Bn٣�Ä��r�����g��RM���l�F�=4�_�\ϜF7�@j�����%�tb�֜�֏[;e)O� �Q��2d��]m��v\qc7�|z'�)J'<�_����be������r�_)9��@��cb���w����4�C�ՁJR��p��0RzBNєW�u�X���K]S�5^$=���(fz�����x��� �_F����Ȣ��[ѵ��t���a��!�U�<�i��s4�O��"��L����%���i1��?�f8�P'Ȣ�uߍ���E�}?=�4����i�C!~,�� �Ld�h��;�K������k��P�⩏��DQmr�Ť�.��&���U����
���D��+���ϰ�5���#�1psf�����~�.H��/gy�-����w�H\����F�F��^�h�A����@��bt��PL�Й�䱣I����tݏZ�D�8�CA��|t�,Ɨ��ޠ�$a��=��L�ɢ|��n�%���Ph0�H�i�@�N�D���V�C��fm��Aso����Eۯ�����P�����͎+m��f�{��{{���m�*�.��x�/���v21B7w���|�Y���a�]��d���W��I�<|2��1Ϳ�Y����)�1�	�1d;�XI^��ɛ,U��6���g�|W�~WDlЎGK�)ש�;D���t��M��Ȧ��i��y�נuVY���3�6fk���z��>0��e#u-Ϝ��"n7�K���5<�*�B�í!;m��'�u�����m��)f��_�pg�n���=L�Ȇ��;9�a��sv��մ����f. ԋFd�M���`��U��i��q��]vm��}�u��r�C=Z���~�&�*�b�0!M��Ǆ����m?�R���aVV����޴㺇��A_�A�Ib+:�q��E����;Y*�ڻ�p��K��ϯ]d�2��dO�k���G/YCKV�C�#(R�α�Z#{n�x���پr�O�a�3�6Ar�yX�h�vt~��F�d���a��u-�����B,�y�I�c���qams���wƟD�N�����	sb��Φ��S$���03�_w�hY�����[2�~������w�p�^9EkxI�z��N���O��ߐ
�2�-�C&16(˱!�D�|�͍d����F��XdV��T�%[��?~�u❳���Kz�~�|I�_�w��~�.���w���.R^L nU-D�^
C�:�+��L�?�씬4��D�qc�j�ါ�G�(�B=����-R�4.L�e2cm0�k��Z�1:�����a5�����o�#A�$��J�vdZ���3����������������n�qsy6�@�(B�Y>����>訕Y!g�d����'s$rŀ֡� ��B��g@0���D[}�ˣ��IV������������
&i6K���	�~I
����ޮ�ڔ��h6�)q��_��a�����{`���	8���:�bt��e�* *,6�)J�-�lf��-+�X�^�Vx�����H�5�OHY
���d��.-��,�4�L6)w��ы�.\)'�@*�&��l��>e����Fs��Qu��1��l�Lx����i}̼�,zL����3���&Ͼ��=��[$P:��mo���i�Y�U���L��w��<�����[/D��s(.
���4�����ŢrG��/�ޡ�1EȈ㿉HDv���v�����?��#�P��_��N�QO4QWn%�eV�qG��u�9�3���X0�Y��yiY��#�U'��c���>����Yz�lRx���>^X�j̧�Y��&��.����%�Eh�GO\~Tl�#�հB�YM'U#���[���άK� =z{/e��Zz�0�8���\M�]d�N`�K��C�co�MG}��B�/ߥv��O�X�~GA�(��ɑ���e�-�?}{�7v��ht锳L�r�vO���y��ɷ�؊��ܷ�h� �%l/A+�t�5�M�ۖk6J�^���G�e�5p�*�� e������[UU�_0pB��Ǥh27,�����G���Э����R����})�J�5p�{Xr�.�E����p�I���ߡ�CYWL@����7&r�Lt���+A�Uq�q*z�*�$���}���H܋�M�[�C�M:����n�+3�L�u�-}�Ϻ�	Y�lB��5�3�A�B=5�$/84��+�9�3,�T��#W���6ɕ%;�)%�T8r�C����,1���/�xE��F$.�c#�&5��u_��pY(D��G`_����	o^r�
?��q�D�����f9:���c}�7yf9]��R�hä(Z� �`��GA�"��Z�\|�:<�,\�\G5�Ȣk ���Id�P�E���T"�u"ړ����	Fn�C_����hO��_��F��2q��}�݁�Jr���]t��:�r�k�O���$6�gwR��.@a��^�f�MS\-�h�Oa��8���;VUɂ���8?P�Mp�Ӏ~��ۚ�b#y>p(����3�P�_*�3)]�u�:�CY�{�U���La)�@i"n�E�ߣ���n����A�^����{'�~��T�QPaЁ�3�-�O#)Q�:�r�^�;�ɶ;y��bg&�i�����!�G	���.
�G<�~
f��r�p�^����'JM��� =S�i�X��	�D$��=�ׯ�YY����ۺ%@�Z���)�Z2}����+ʭ��H��= �}sf)r����to�ΰ?5���M��A��t�`�5�M%�JC��I;]�nl �J���B�4	��*���SI���f"����~�[
� �.��'�?���d�V?�<Ǘ>{^,�.������0M�<��;W�{5��\��z5�P��,�0���]����>�u+��hG�x��n����ץA�a�GK���$���V�T~u���^���36�5N�����v�}A\p3�_n��S:�� ��h+!]5?�t�q�yh����Q�~Y��e����� ���'c<�O<��	�=j��M�o ���<���Z����K��/�?��K�1�36�4}\��p:P�]KQ�}�&J͝�{$\���c�S�%e��R��=�s5c�� P]:�����Y���v�;�IF�s�P�t�O��,I�J\�(8F���
:7�vA_���z�U�ޞ&����*�X��/.����`�ۙC)�u�Wy�pH�ҟt0!����F����8!�!��Yx k�l�k��޸���V=�l �T���.�=ͯ�V�P��aX���O���U����D��Ux옊�����:�����@�yZ �W���C��hRԻ��X��@��3d���W̉�M������~����L�cL�"����7�\|�\��W�F�:l����s,N����W�8}��D��kV&�c�&l:10�BcI.��Dr�=I��!b�G{�yi#���2<�N�l�u�A�<CߒJV�j���y*S ��k#�p�������N~ݙ�Z�`�xj��qp]�������x݅�����`�M��u��6 ��T�H�L�4�+n��8�l�=�X̎d��9il�i]?(DS��k�[��y���?�;�p�ߊ�x�/>y(9�75$+����D�-��:}3K��y��y����4k��{)�pWΒ�3M���8�GT\ ��X��Z�� ��V�� �� %�&-b�v����Q�}r�.X]�5/9b��#�����Lp�|[8v���l9���aԖfW�����֫��V,q�;�3X��h2TFM)5�e��յ�R���0o��ԓ���4C��NdqE�^��QC2|�NC^�;[{D��WU����l��G�E"]i�h���V���;�N�Ɓry3D�m�j��.��"�0_��Rz�f�k=����G��Wt�<�1i�B�z-`0�����z<���U�D�5<�_x��̭�/m��ە��EƔ�Z��ҹ�K��Y>��8�p�
D�RL�
뤨�+�����)�q��Ѝ+�K���XձIjA(�HT�����k�o"d��xà+­��KOhF�Y��9b�7w�yy��ڈˌ���{�jN�ˋ��g$M#I<��m���J��kf!�ì����}�/���I'���>ޕ�9��*��M���綻y��Vyt�D�G������]Ԏ�FS2�*��]bõ�FB1L�]S� zib(�n�f�n}X"�46n�(���R�Lw9#��͔�(��آ����ЭF>��]мF�f�z,2);{&�M�44��o��ZN~�۴50[������"C�qv�+�#V̈́����g�,���y,��;�H�OK�8�Z�O��E�(�(=G!e�d�C���.��0�l#ҸC��/Q�Ⳡ�N�V���N�ċ�d�:v�w
j�ul_NKfoԘΒ�dL;�M��F�A�3����MF0m�3�Z���r�S#������^+�P�����x��tq!v������J���+�hy�=#�|6�y~e��)������N�s�n� �ڠ�Җ��/�Xo��4]sΌ&fZ�%�?A�		�tĠ!�-�eY�=�R�kj���zV���9��^��D	[Фc�րl�nֽuǭろ��M�g��c�\C�-	"�RX)�%1J�1𮴠��
�'���|�=N|0_�����o�e�L^@҅Ğ�"���(�����f�L���<]%)oi'�+!�o�p�
J�B+�!o��4cOn�ӿ���C��{ߨ_��)�:�qh�z�6F���[cjLNޞM;����L����a	�E%v|J�v�E����6)8���+W�m��������I��h�U���vٸ�l���e��)���+�0�MŜ��w�����<��.����������p����94f�1b���ϙw�L�W?�B,�2'��L�fh�B�^�w�4��^��[LK�������L��R)k�S,��X���?��Fe a���z�L' &�LUJ{99.|>���т�-�ެj2�=��W`֤Y	������~���M� `�����H�C���|M�["u���=���(>�}�����̻( �u��U�h���zS#0$���"��'Yݬp�A����zL��)< Xj%�#�a�z��uV��&��3n�qS�`����}���7:�"L�I�3YMQ�N�+��TT���^�� ]�&�wތ\���+�U�-��Mb7L}s�� L[�M��r��~ζ�|
���{�1�(�騉G���t]r�O��rZ�x��fϯ�S���殈��c��hu�Q�T�n�6��.�_�wX
D���g#K'�aZ��?�Y��tP��WP�c��-A���"9�$�y?
�<��O�����F>�B�{�Ђf�J���ܠ�@�r��ʹz �v���5�"M@�<_��4*k��;lZ 3K� mE�jT���cccJ��`��{�>kr�����Ά�f��7ƌwg|���� 1%�.#�Q���0W&���!���;.TWဖZ�v�ڰ���fdO7��)��B]~��8���2�?zD�R����Ѱw+��������P��>��ǟq�J	l'(� :�Dڳ��VfS����wH3/5�ҹZK�>�������WW�1�[�;��}��!m�܈�#��m���d���߮-�B�G͢��u�>��<�q.��7��ՙ9);c椺��ոs��@�|a PkW4���냺�j�U��J��8�1�Z�IyYs�#�Y��nxG�UM�%� ��2����E�ҏ̅�-��]�g3 r���4pً��7L���
g��JY�ϑ�/��S�U�|��n���'��2lHoV�;���W�z�/�n*G2(�t^nE��3�-���i��
�(f����M�u��4�1�w�*��d���]��u���W��L�ֵS*���iC-$� ��%~d��if���u񽘹(�u��#�� �}�y��Br��*]{���da��hiۗ1K!Pڟ��9aOV<h�n�c@��f�Iӄl��и��L��ї�=�r�����®8�Y��R����a�<�u�������?�c�4SN�8+V\����k�x�^��RV�o��7z�n����Bz�iq��i�3V ��o�sm}K(�'M*\3�R��-�b_��J�m��E��#$���V����z�^�r=��SU�z
�FOj~����tc�Ɂ_KxW��	@�,J�������U,��+�X���0����by��/J��B�')�^�!���`k�S1ʺ �O½��-η��k��f�U�����3�OV��d�.5`�kw�JL�Q2�d^:���ws���t��rt�@�4dh�s/*�������yjG����ץ�82z�^\�kͺ|�I�D���qhu���~G��=��{߈�d���a��~�r�h�o�u�J��?K�H_#�a�5�9p�-a�%�S-B�M��a7F�1����
Xn�̷~�#j�%���[�?4����Kc��>IC�j�9H-�U��
Q��T�Ïu2y�%2�6:`�4��<�؟���	ڠ/"�⺅7(��wjp���������(�:s�#d�* @�LZq)��5�[-���.���ٜ�	��q��ݠ+���&�ÈaF�lv��J��^MK�LP<b���P�ǦX�N�ח�0�^Zb��׉�W�\a���x���Я`�����vR5�/y�ǂ���>d��Ҥ����G��6W!�$�U�ʱ���ϿB���P�7dG��.%����_��l�*5|�.���°m��@Ŕ���ǫ5h
�^�A=a��2��5��h�̭�}��Ei#9�z�~Ĭ2`]Y�^~x�;���]B�t�a�<(bK�ߍ�,�U?/٫,�g��g�8��nno[(>��M-��ۼ5��lx/2-�PӔr�gki��f/K�!�M����_�:��ε��6�'L�����q	�ӗ:���l@����q�<KU9��<�Sth��;�-7 �ه&�Z�g����!���\B�U!�=9���e#����n�/|}�LC��V���]҅����K V��x�L�ѳ�v��
�N=cE��B뽸o�^�,߷�m+A߉�]�R6�!���t�zb!���A��S���i��,��k���\�og�����M9{v����~�؜�Gx��q��h\Y��+��J�f����AS���/
d/)6��_��VB�byQ`���T��Bnn�⥵>�I�l���-�������,��H4��B�X���5m���i2�dWiK��U, .y �������4��d�e-|@4DrS�A/�����(z��s�G0w�α����j"ؙh�{�s��7w��FT��/3���C
'�)��wގw���K�S+@Q��&�o^�?ژ~�i8�t�C��+��!�4?�+(�j��:۟(o�*1 U�g�S���wgg<��O[3.f���l�<��jH{��0k�o���ԐD��6��m�L�h�Q��כs��5�����j��9����l����ԯ���3�R7&�T�$��ˬQ��ludQl2U1�Sk-G>��Y&Ӻ��p�l��`޴���2����l?D�b��q��I�D�|^�b�PE��Tv��tZL�,��e_YL�If{���Q�{)0~�M㟮bS��#���0)a�S;��W+(<��g1]��Y�jx��w&��+*�%�d��/��l!�{j(�r#+�![��X�P��`�T��}����'tf1��Z�!�;[��Is=��������Y1��{9�� J+�L�׀����g	3�2 k�6�3XXi���z�6`�ON'�u������&e��'��V�lT7�ʢ`�(����ܥ� ���gu��O
}��|�L���C�ËA�+��,E��z�{q�[&j=ݒ���d>�_��o�C�o�蕣3��o@�T>��������)�j�<~*�V����Y��֙O����N����z�}���<���ڊ�D�w'5R,�}\�^�O���g�S��MEO���)xPK2W"s��;�9d��8 �t+�E�O�9���W������ �N�1P�hq%�PQy�[��}�S�	�F�+ͦs1	ic#w�����e;�7_��� ���r�zN�a����a����0�]���y$N-;�k��A�d��;H�A�12�XS+��sHx]��5��꥝T�&�V��(d�5�b��X��~�[���H��^f�y�.�������H[�������%Ǫ��{4��<��tN@�>�(��t��q0��x4�MA��9R6���l�in���Aߊ��x�
�3ﳞ�������E�ΣT7���ܪ�?�j�ۿ���9���*Kx�����̀U[ ha�sS�Q7H�_�Y��(:4j?��!w�[	���������ыw@��f:���d�@��M�r�dvKэ~�.���3�-�L������7i����2�/��z��(H�%�vX9H���I~�����m��@^n�Aɷx�f�|��k�qk<B��%�.2a���%n׾>e��9�=�41�Zo�<=�w�Fk�/Q�uh"W2E��@�S3"���Iֻ'<C\	��95���y}�Ͱ��K��Dv���A&�����*�ֵ�%h��T]��ϖ��]&��H�A���.n��ԐE�*q�n��_8*`�R��aA"���bicu_�a��l0��(����0d0���oP-���Hw-���i�|�f�ѐ�Jv��lъ�J���c��FCy�ĽWx�v�Mv݌��a<#��a�����̖�cn��m��!C�p���7���n��Da]|��%�a����U�N�"�I�#�LaW�5�yO
v��2�9(*}���K��_#F9ze ���8�Y2d�B�'��z`G���[���!��{Vr���;�Ϝ����*��rD�cnmƊ���8�Vp� ㇀���Tr�eV�v~�y�^����3)á(�$Ι�#fxu�k�Ad�6u@[�*h̘"��)L�����TS�/�.��/F�9+�7o�	����ri?<P໓�>����>Q\������-uRX/���t���-r*`�kcu�4y���:��Tm�B�wy��9	�7=�A��z�3��BLd��M4��/}@���*�zӖ� �=���`ZrN���%�\HVɅyc�S1��!'�G�h��w1i�1=ޘ�����R�5�	����`#��
+r�@@�V���<�Wh����j����]�`���>jzz×=�"f�̑���	/�+�T������FP�Гy��d �A�C�R=6A��BN�]Jv�؜�c��B��i�[n����t2���Y��s	����E�e�IITY��n:X�6��\�c���yY��
�>�\����C��G%@��Ğ���1��E�p��� ��F�t~g�;x]L D*e]��u�fN���1�c���.��!���K>��K4�@;��}?%�~;��hnL��oe��J1�0]YvZ��K!ō��W�)�=�Aue,`�sk�nԁ����v5�Q��s�T�q�Ka5�����E����[�Ѧ��|�����	�*��T�RI��K�JQ�⭿'�$-c��SJ��ˌ{�6lK�}��p��0�Sjb>(�/gZvr=Ndc�z�B3���tJ�"`�@���r�}<��!b��9������҆9��;�{@�ߡ�";�	Q��:�a���+���=69���f�E@ ��� ��N�RT�
'�Ux�L��&����7GC�W
S��n�7�p��ا�@i��M��A��"硎�O�Z43
	I�Xʞ�^d��=hThЌ6�)�yQ�J'?]Z��P����`A=H�u�=}�4r��A&ktP��2
���y�2� ��QJ\Oc��OY�K��8eo��o@n���L����q%+�#2\F�����
�9Z\�2��unI+���,pJ���
�ܼ����_��^���������ٕ���k�Q�I�͚��Ե�|�h]���W@�'��Q����6��j�����\�@��+4p�ʗ��î��Kw��9�aQ��eěW�f��$�� %��O�=��ŝ/m}����3���F ��G�.��Ȩ�k�����{��e�j�m͘����Q��h� `D����E�=5�Fu��K%O[9�� 9���w��Yc6�\�c+�r�6#V���p{��rG��@É9���å>L�nf�s�{늨�1H�G��U�"����QO�D<��Yc�3�x�`p��?m.TQ�
@i����  ��\\��7���N���|v��;R�|�h8T��2���q(�k.՞�n�]
8��q'�������qoӕ��b0ɑ�C�����+�X��y�D���[N����
�;&�6_���K��H�x^�l�=S�|��ڈ��~�~|���쾡�
;��u��#,l[��%һ������i�rFo��΄����k��fP|�c��)�tk5o�c}6y[�k�#��C��z��~_g�8�����ŋr�T`rɫ�_eP��=t����u}����7�Rj�:��z8�lu�U*��HD֠'y����]η�C�!+0��,����
ێӚPTs�S�.d�j1��-c��e��Kh�Y����$��YԟZ����:�m���8�6�5&B\R���HC�I樧�'�Q�+��/Rħ� ��y�=]���Sc& .�N���!*���������8}�vĺ�>U�⼭�k�G�H�� `�Ǟ�1��̳�[R�S�t~����	r������ސ�迠۱N7���fB"����;�u�t��c�N1l�?��3]���i��5;���ot�RS��îM<�����G�}S2ne���*e2�bc�ʦs�<�h3�y<����5�t4RZ}�#���d���|��U��k��gv;?P�<��_ߚŝ���i�� ����X@u�7��T �p��㪂�u�D�b�:�bʵ�R.�ۢ��+���b>h����"jU̘����_���]]�z��k���S+�#;Y�B���t�WS�����U�ENl5��P�ԸZ�@ƥ#S�����`.1|G˓w�U��{qio�4�G�L��YƤ{�y�	���i�Ŧ;�zf� �@���AQ��h�Wr*d>=$)�o�E�!��o�z�޳Jp���^v�����!k��}�*=d.����P�xE9�D�U(��y��Д�'���������}�n����:��A��u�Ɉ@��(>��(�g�߾��ɞ����fe�ĀfG��_hѬH�C�yF��[H>����
�����
ULh�.����>�5�D8ţ��]���}� ��\�	�*G2Z,�����,Ҝ��6%�x�Mx��@�+sAf�#�u^�F�e���~�g��iw�����5�����ϩ��%�{�_x\�:��{U�Tx�����o�Y�8���Ӕw�)a��i�"8tKBS8N����ж��z.�N��L�ЫX�`��ƣ��}�7?Q�3�g��#��vۛ</�2J�#Oc�ݟ6D:k�Z��֭�P�D���C�p蚑�ώ�U�|#�����|:���@vix�xG-����� kn��Sa�3'�B�M�+$L�R1�a�Շ��ܫ�{a����w�/���W�����y�EhG#��h-�na8�,�����j�A�a7{Hn(��B\,�8����{���(��06����()ڥ𧴇Ca$,:�%��ER{����y�5N��i!�	i�6B2���9SE��Cs�E���kXcx�m��gjE��'�GBK��[����c��A	k���B�����Z����TZ���|$_=��\�{�Bp$&Q�y�Z��jJ@׹��l�>��1Љ.�:i���h4�k�S�*��aY��zY(�->x��@FE����dw)���yoD�d��)A7R�@`���"灏C�ٮ���n��	rW�Md�3��P��۵x0�ei1��&�"6����x5����b�'��Zf1+)l�Bǐ�;�C�lǜK��a���6^��%���o�@���,Kh_&���6�0����3n^4;,�g�����ňg�Y�*�'�\=�C)�Um�>뗧�G��0y�W���yAt.�'��Z��/:�����7�;ܪT/�J{�+�A�x��O٠ޝ�OE��瑞ֳ�x�wڡdC̖[���?��Yp�,��K�ֈ����5%OE5�!L�~�V��1;�\oN'X雨N}�J��5�ᒣ|�h���.	�7�{w�I��A�m���e�0-:�.[F�����>��V,���p�U�и�
5���sS�p~�g��Ӄ?nxDkG����&��e��/�<Af�s�����h{��Bkf�G}�	;b?��Y�/l�Y\��-+'&�������[��3���FM��{_�T>DFvM�@q����F�P��$J$N�(��.j���y�>��OW�D�lt�-�e\��8�6:T���0|'�U��*�<u>Ȩ�7�:L��+;!3M��j�_D�5���`�x�doY�f�)ciw�e|�m�)��3�cng��=�bz��TW)G�F� 7�׼7p��p�ǅ̣7�]���&�`�� ��&���/��q�g!����"���$�B��B�����j�з^���8���nM���&��l8җR��K�"zP��I�W���3Ǆ����BLa�ieͤ�Ƶ��j� �H�'i�4仉�/L�%��c<4sί ��4Ł�!M1h��C�xnB�o����h��E�Ju����%F�AFC�5�_��r)޷G�;w��7K[FPg��ﳑ�rBiϨۊ��U�gP7Y�4�@�?;�0A��[��2>�,e�I�Մ,�#�}]_Ւ韑½e���z�ϼx� _�6)N����"�O���,��/3��������24܄����,4�:dt�6��C�� T�E3p�{��;�@x� �i.�f͒$ G#l�:��I��S:�[AG��$��q�|���u-r��L��h�2����̖�����k��S�]��n����զ��v�Q*"�/����]<����q4���[B���j�L0#���3P�g�cE���S�vn���.k�,�o2��!�̲��00�ӿ�5��/��E��Ĩ&�DX���θ�\�tvqd�vw�(��R�ǽҪO�(Q���$��� `��LPJj�9/{�u}t�o��o�?Ԕ�06� c�Y힕�?5}\@i$��L]�QZ$�y��*/�L�W�+�٫������,^I�G�p���-�%�������|{��C~E|����+Ț�{oQ]!�ኍ/���|�8����$�Q���Cb�|Fb�������*�{�brf�%�