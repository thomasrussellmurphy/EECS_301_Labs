��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\���V�fnvx��ÍG_;�ȅe�~�>���9�>��Y;�0GT��}��E1����E�[��G1wSd� ����z��5KC�J���z 盳��t\Xj�ۺ���V+� 9��G��BOێ7������u��t]x���f�y������K9&�쫐y�ݙu�I��h���R��XN(��b��äo��T.���B��˱�{��!33u+�❊��W���IiY2,�o,^O�}l�ur�oJG�S���Vh��90��й�^��Q~vYO�Ԣ�画d�^c��g��F,�xJB\/�<��K��[�5/c�� 8ED#;����������\'7Xx���u�>�A�|��	Tt��j�WF��`��>+� mt�F ��5�G�.���~N��-_y��cc·����O������%��%�����+,	}���8�r==�}��d+���r~2�d٭�%�	�`�'ɇ�"[���	L��oMzǺMw(��ė5�U��`�UH�W�g�.��E�4���4�>C(��EK�)��-$ة��LBO�[��9`a1�T�XF"؃�@6v���/�����	p5�Q���hÃ3�P"� ���c,��T��J������g�5Ћ�r,�{P�|�)���o�)K �����Ǌ˒V�Ph��f�pog�:xQ�Qc\�o<b1>�'U�H|��@N��~s�>��F�稴倣Y��ZaƔ/dY3ߠ�63��kĮ$m�D�Z*�����d��ɪ������' i�]������V�q�*�=a�?SMc�ϟ��z_�%�C�$A�	e�b=�Y=$��eD;)�u���6jNǋ���Fvs��h�2&'���{���E�jn �=��6���(�p;S�6
�%ٵP�-�3�wH��2sKڔ�7*q���D�"���X�$�]Ʈ -�:F2�NgBƿ�C�+�Nt1����0�/m+'�����3�ft�4�}�fv��ϩ�ớ��&:�x�$ 0�"HS�`D%O D^W��ֲ/���Hx���a��*=lBgX���6.�G3 L���]�
�;�n�8?%�.n�S��Hy�)֝baa��� U���J|B�j#Ȗ�7@�36ub.�8ŭ�Ta[Y�Ӏ��xH��{�_ee��0q3���LޅPYI��U� }��k"�G�"����d��6B�Qo��ԕ�Ҥ!��=A*©B����nj������0Պ��*��_I�V>L�i�g0�)�ׯB��#��D�M;#�ذ!�;>�\�x^���_��aY�4)�˥�9jkLyg���.��#w"ܧr���vT�ǃF���ġ;���>��6�$f9NQ��d�p�}Nڰ���࣠s�C*�	���#-�<L\g%���۱1*n�Zqz ��}�3B���������v�ܞ��Z���z�z�5�@BI�nz�Av��fVA�G����9�DB0t�i�%���i�B�j�~�B��D���?�L�y���Ta�K
��؎��j �4���P](���!�0r������Q�U� �$Nͧ�Ğ�*;'����R����$�:�iC/��A({�8Ҝ��v�*P���L�q§N5�����j�?�9�7Qq��x��},�
�A���۔��.�v����=b��l�T�8����n>��Ziw+��B���,H�r�|�m�/���7���6]��.t��5�k��:��T�R��
БuE���+vG���,�?!��@����x�/f�O���@�r�>�2D���tP�%�E(2���u�����9��ǓԴ�+[d���5O?�p��UVL�����[t��z����	�\ ��٫���%�<����OW�ô��@�[:_�}��Eg[�`=;v*5K�_��zJcIV��o�p�-dYL\��#�MOp)ن�����
�'�=��*���[.T������$s!�E��E��	����:�g*P��o��!˨�_��k���n%���0��ǯ$ч����(d[��π0@�*<�؀��/,B<1��%I)����� 
� ���F��R�q&�X|��(�=�]JFaK�G���1H���XV#V�� �w&Pe�_�.4���h#F�aT��hl>rlA/v�Wd�W�H{�.� �A'Gv�Rm����E&7�W������ߠi
�ݹ;Z�����Iϗ\�@��(�M��}�oX-0�pZ�K���j�DޛK�`ؕo*���e9��~�����C:S�α̬���_\:� }���@wfj{A������$�|��K�n�Rg̝�;S������nڦ�mu�,݀�tJ�p�7��Dr!�yWɻi������!�~D���6nˣ���!�\h��R 2�7`�?���bV�.�Ǻ�4z�0����w��hA�9Ra{��	��ǎ'�2�H�V��i?����4۞�N�d�0ǐ��${��0�!�@��)E�C}��T,��щ� ���3" �8��r �Qص���k��&���q��3g�~l9�qY�G�'�����$�D�k�ӆ�/;g��֮�.Z*�=�%LT� �bL���2ޮԼ�?��((����N^J�Ϊv�a߉��a�g2,�R�\�2�v�+�rP�\��;Ƌ�g;3`����zw\�J�0%o��ևb���aoD�8G�&�L��w��b8�_���4�W�_ Ԇ8?˺	 ���*t؋N�M��yG�([�M>(MЗ���b����G�l'�\2z)܁4I�D�&_F?r�W���ǯܾ
����P��T�TyF�k��k� ���ۂ��tJPɩ�@��kBs�	d!1���6rM�iԧv6!g����G+MW^��Cߥ;��Ӻ��8��5��moO��2㜔���W�璍b����DU�D���Րr=~�)��&٬8o2/t��`�C�5Vj�I���PQO��K�����-6���_l��aj:�s����q3-л���5��9�(IA�+�-��'���s���Dʹ@�����j��w~���x���䥜b���|�gXv�N���C��sD��~�v;"�j\_S壐�\��̡�	g^����"ny[ {���3a���|}���x�{�)!�g�����I��<���96�V���X��J���f���
��6`<�0�?�/X�j�?�#`�����s}��ٙ�bL2���ڭr����vb��H_��h�����Lxi0������2�n���ܝi�i;���dM�X|Z�m�PIݟgz�,�@�G��T�b���Y^�[[�'���~�6��(K%w�]b�ce?)��nL]rZA����_�-�����k�m2!�; য�A��<- �'\T����Z^%���#z��iT�8}6�Ï����E��cj2�y/�)i�}�Mk�Ow��BQw��Q1��T*)�Rg}	-�H�I���eh#M*v�!���Vr������М�J�5F%˝����r��n�`�L��2ًT����,8R�Rݐ1;ބ �����4>�yL��s\Y]ǼV�&�3�V�%y���r���=ޥ�ƎCsM�;�!G4P�8�4ȗ{��������հ}O�|;8c-�����W�l1�b��rF(�+�
B���<��bL%��9m�3�}�˻B��0m�_��b	_OF4QN Ɋ"ѫvĄb��`���7Z
���%�p+C���|J*�
�G^�n^�(`ko˪I�pJ��)����T�+���'��lx��o6�]j̡�ܵMf��@a�^t��Q9���I���w�b�������-l���Xt�@���4�������VC&���#����ߚ�?(r-o�s��t)��+��6f��E<�v��X��ݒ,djOU�[ t��z�ʁ	�4���m&�j=����~��[���"�g9x�n�����*���kش1a�S�^���v��\vL%��8�CuA�_���S?l�T��[b��5ɏG�qt�=��$X{�\^�Z�v�j��b�JLS���y�x�6x���P��	�OES�І�}�4�3�L�.���VA��e��e$Ŷ|���/�#Rx�(�=���ikl��I�������뇲/]����LeǗD�N]�H���*�8-;Ǐ{=o�o���r���Y��;QD�#&-��Y&"4J�D����6���^xcD�m��� 7g%H����bK+s��	�2o��{��9���`�_�?�ub7�1����YË��1�T�j�r�aT}O@��*^�]&��$m����MI�O���C��j��&j�m^uk��R�k��z��VkV����(ZhH�1�����D�n����K���zk!�L��+���G; �ܝ��~�h�W1�h�c����z5mi�I퉱��p�)��T��D�+C�bF�9��fdr�_�-}�m"b���=�qk٧ �{%�jq��8���:��(�øL���:��JU�Vʞ������^����a�:F&� �uo���J�{�:�P�g�Z$���ztN��ae�������(!2ś���O���n��9��~*���_I]�yk�Y��7�%0����;̙d����ԥ����,���]>��K��w��r��a�֟Q�������\	��Mob�>E2Fk�Kx�-G��b_��@�1='�isk�������(TV9��?	��?�	<h��Q��l)�30V�X���E���