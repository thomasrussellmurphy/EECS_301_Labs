��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8SjfSު�U���K��)`�(s����2x���̬ʐ�QO1�?͛A�~iSAUo��,��Ii�F�_#�� �K)�r���I,6l����6�0�c!��["!#��jS+���u�]}����AZ�R��fok��V�- ���U����L��p
ZYW�9��1R��MAԪ��P�K%f)g�[�U��^=>��AJ8���|mn�������\��uJ��װt���K1�;����͑�����S�H�~Y�ɣ�Us�!z�����cH?��W0�ք!ɑ>���4����9c	`�%�23m�N�ݿ#��wt,Hp86v%ͺ`sfr.�(zEe:~W��/FӤ�a�f���t�2���$/E9�"�V�1%^xp�nx]�>�ړ��XR�T��>���5B�g���G<�R]��{UF�'��b�9b
Y����Q�
-�=!�o��:M`7���ϝ@��Ok��s�/t�Y�u�_�v�%�����`�7��x���>�uIi���1e�v�ou�L�paϣ�,�Z�\�qr�iTp�0�����߰̾?�^�"�GXe����v4[�R������`�W]I����@�4��_c�L����O����O8�=��}-8�X�%�QR����;Q%0�7ʎ�z�X�1��#���y*B�nŊ��Ni��}񐀺H�r�Ek Mtr�XsD��5�3p�qC_kǟ=�N�����.���dW��ѓh��T���t�^H�n"��T>��G�Q;�� ��Z�d���e�eW���a�͠���5,������[�.rݩӓT�B��S��"�/�d�vC5��E�ڭs�zYf�J���n�`.��ap9���
Ƭ���|?�v�X��B�@�$���6���a/����-�d�ϲ�pGůd�Ѓx���ځ��܃��^��h�Å�mG��������˯*q@�����o�񹇙�՗l*k�3&�����۬�tG�}qޓ-y��Tu��@�l� �@���8A�/�~g�����"�r���d2���@2K�A������@2I@�O��?Cj�^P;��a���n��NM)����������j.�����2¿�L��Lk����\��M�Jv	�̤�Ƅm��
����}ym���J����T8�H�4�h���!P�<���sJ�(�B{O�o�}�%��E fFGg�Ɏ1ـq7O^����>�*�N��d��f��#0��Y�&x��K�T�J�� \^2{X�}PSe�[�Z��B_h�8@5���sr��]g!�<,���Y��U�)������S�BA�h�9/ 1:r������8.�R�#Z�z#`׳�FT�m�S���b>0@��l�Z-�l�As�!0�nώ������PTT�:kV�{;|�:�U8��z+��aڳRv'���Kn '�E|�e"x�rz��_pF�������F�ۅ'0�3-���g�����eD��1y�f�{���a�]H����
��B�����2.$'���I/�&E�2!�oj�2�.Ο����KQ""�"p��?�l�n��BY�%���x���������(20�g��L��_�2� VҞ����w��R-5e����7A.(�˵,�6٠HQ���<,☦�V�
xx"��N�c��e� -�;R����Δ%�f��	���~|�(R(�	<�F^Y�s�ǫ)O�N�Y�r+V�Qg{�)��D�Ҟ�W����;o�6M��|�����"iP��.}b��XU>�szDg�}#n9s�k�7ͫ]�P ��B�;�ī3�txq����U  5�&�����讙NE��ݜ�7z��![�D�Ϧ"����&�NG
��'�^�C{}�?*�{�l�@5��r(A�?��RA�s��x��W:��e���ӑ���)�|튺��!튃QD�r���
}�Q�H{�6��G��puL��R!�NLq4�&�%�0N7Pr��y��{|>��n�]�r)��� �1����:�K&�û6❔~7(Rx�_m��txHĐ¯��lb�w
�B�IS���ܵju�Y�S�1���W�\3N����{ \�2�u�d7��*�w&�;�����n��sL�t��gJO��E�Խ���F��᥆���Pw1O8H������`bb�M��x�/�.k�*�SIS��Ά���̠��`pE��e��"�Q�j�qzKgD���;�O��oM^Z̚��5H�|JE�~���*���<���Asx�͐7ǻ3伻����OD�-q�0a���
 HR��:��j�����	$5�
*o�=��#�Y1�Q���Ra���Il?`�fd��B�i���j�
�d�T�����
��^��ysS�%U޴�J���Xo���ټXp����w�G��y$���<���:3�ܼ� ���Ŋ�ޠ��%��]�-8�s���w��q�a2}a���0<m�m:�{:k��7Q�՗�T���jLƊ���V�� �3v��D�����{��G�qְ h�/P�@��ဵ��j˵JG_���܌�&;~���J3|�A�Saq��[L6����1ck�j�H�J����y��/�˹tG�Q��d��V��d#Y��̾��|�l/]P�R�����D0	l�t�آLe|ea���^�j��
2�C�8��yPF�޺ӟB1:)o�w�����EB�1<�b�@w�����dv]���)
D�*%SO7"ߊD��ׅ�?���櫺���X���Y��Buj���Ċ���e`�S��m^l��Ew6��n�~�,?�P�l�a�5�q(�w�ȧ>szm�d����k��V6�:A(E�%4c�\����q�y���а�HBL��D"k;��b��Gf�a
�����[��7����d� �V+B$���N�M��4�X46�5,R�k�>Z%{��i���k�(M�}tb�sCnI_�y�J��W1r|���6���{IL,��KI�m��k���4^u�PI����I��Ƒ�|x��C'V����_LӤܿ���I�9Q�<]WVԜ��*�9������P��s+Th��*�ѡ�?��h��b��~-X���2�e���7j�
N�~�����7�l��>K�j�nGFMD7��}9�aj��N�.x��^aH]@f������|�U�#,ō��!/�������A5�ûik�n�����-]��<��p��{i ��xTR~�v,n��;��E�(*-iP��l!Q��wK��~z78�Fm�.��6�۸�5�X��Ό�q��������vvTUN
�����F�j�1<�v���r�R�%h��
�?G����7���D1���P�D#ɑ���>A���{w��JjR�c�A=F2��$/�Zri����f,v����/ЖI����HiF�MO�NX&����U��DM�M�:c��A�V���� ����#m��)[1��5�ˈ�f\�&���&�q���TCl�1����l�V��f����#jefA� ��q���m�n+��^(1'$XE�	}g3���»�sm	�h���E:&���6��	���i+RrE���y����C��3��,R�9�	Oz.h#DY���?ȧ�i�^�����J]pA�"Z����Cw)D�/�lv\4��CV���	�X%U�C>��f�TLB��n�����������9;vLv?<�mYNr	� �vq�՗�j��*���6��Po�O�h���D��wc�:�G!3W���s�z�5q�"*^�Ou�"�*|��pS9��>�XV��u���˟!{�.�����X�昃�V�))$u�<�݇j���"�B��a��8�ۄ�?�u��j���	�r��'+��DGȿ�1�y�1�����~	Z�J�y��8�̒+�g����*����`��F��Ҹ�7i��^��7���yi0��Ե'hm��ģ���М���^k����&c�	&���'���-�D��&��jva����Y8g0*eS���ѽ��>���%�$R6�=
���� d!�p�e�
��0;zn��.LY�����0�ը���������ײZ��S�Ya�C�;!-#��R��(���������);=��G���}�
�zT��Ȑf��}䬬1aQ<��܏�%�ln�B������f��9A��ўv��w_,�G˖��j���X`��"ӔGIŠ.���i��v�>�}
��-q�L��k1�0��u&�����1�$d��5�P-L����p������1#��nd-�C�i��ae�V�n�xy+Y$�S� �F�LLW�:��� S�nH����;�Xs:�w����헐2�N�J�xx��܀Y����.���y� Ⱦ��mf}��go߄��Fy���.
�8�I�1�?rB��d��/<)�G(fr�#�fb
�Q"=��\��PP��gp�5��O�=�%��ޡ2)���Z��;F��U�kZ�r��}A�L5�Q��߲���K�!U����Y�6�A�i�'���`ؒ ��k��(u�۰�QF��~�[��!��=o�/�<�s�HA�c�)"�ěX��Ews"�u��k���N��g�BFf�,��8:����Yo�nƍ{�呬>b5��
u���~E9A��T��S����&d��gs��ţ,�,�5��u���E�&x�'��MT8��}�>�d�8�ǿԙ�~cFB��}�$�J����8��GLq:΋1���������^�d��.\��]�RCg&���������^!z>Ht��������H���F�p�C�9�2��Y�G�5RF�m����o<Z��<I��e8	�U�����(t�aIu#C\�G�K�*�]U[��0
�oǿ�>�l���'Ԅ���6)G�fa�~�����S23u��%*`�6Ե���iT�
���5n�c����~����f+��J��{�H=��
fZ�SCn'c�P_��kU����뇑n/W��	���{'��*���,A.nךþ���\���S��&�Nݖ`��|d�;�&~�O�L3�x�~�À�D/���摖����)��AP�x%��W(Zҿڱ�&p�Mܧ�F���SEk�P-�U�ڴL��%�(�b�����$�^��hi��<�,��n[��(3���V�)�%�Ett����T2Izq�oNƪV[~��u���=P��Z�S�3t���^�=�J���p"��p������O��.�:&^����H(�=�̓���+Y&}l����ӢN�&�O�2z�&Bl6z��H��71k[��a�O����.'Rl	�Jd�}}`�b�^�,n5�Qp�za�����F��3?���M����;�
o�jܷj�QM�˨���_kS�d���Fb��[(<۶�s�T��C��Ά�+'����j�b�}��V�F��x��,yAj_�|��dL��澲�����W����f�8���x9jf<��K�$�t�W�:�����e��P�\f�s�0���)���A<2�%0	���w"O@Sh�'p��G��z;�\gD��B8�!�:��%Xf��c��ƴ=Q��RK?��ϐ�^��I��,? �n�\s�x����P�YͷD��q�c�\�Ș����%��r��^!`����  c�V�F��k"��[��[ݗ�l�
Ua��T��q|tê�>-u���B'��j���q�����է�sDlƄ������viP�~tGG-H��|%{e��wuD-�6�G�g�{a�Y.�|(����|(@q9P�{"��娏T� ǅI�b�G��r�1_@�@���No�6T?�d��bz>DEX��
�{���P0���ݚYh���d]P��I���D���C�`�U]�:�3�>%���!��,��XSbm[[=s���@7�{NcJ�O�"F�Dmq��cف�fr���!a!�����b:����T����2��.�?Qm }�z�����y.l����R��'TΩ��;g�1��0(�G�r�����4��N���
dC��Wo�e�4�w�O[L�1TG|�R^�T7'�������T�G��Ra�����<[�1-���CM�n�����05�uB�<�)�~���bf�S�+J��"M��#���-�8��zݥbY*�(^�<>r��<��Y�U<��!<6dI�¡����$"��^����Fg�,Ϙ���;���t��Fw�P	�뷮,�~-���f��z�����V8��r��c.�${X<�yH��&��=?CY��`A�h~�G&�-��[�3�Շ��h\_�~!rB���I�ڛI��zXo��z����y����8�نΏ
��E�;�4��{�.���{�>]��ٺ��9�����}K
�@�㭅����~��P�T�������\p��i։p�����K{��hjv�h9@+�2���[�|�־~r�30v<#'�x�ViDX�T0�����.<Ǒ������.Ň�ɯ�&��)�Q�%�(]�a2�ښ+��(&
1]t��)���#h��M�('�{[����{ZJ��~"ݜ�ˁ�
CX9���"\�(]�Tf'���7�� �--�Ӿ�����:� bu�F�]Ǫ��C&��%[:��)����B0wIg��0Y+1^��^A������E��q����c��&�O��,#l��E�$t�1�s
�X5m�#�w��1��.�����ev&^QF�KS���t2���W�������)�Ny
UU[nL��(l�x,�'�^ZJl�[�g�aF3u���s��-�Ԑ�ĩ\�q�g�tV�����P���0_�h�b�[6� 	W2v��i�iZ0�1P��g;yy�����;�z*}X;V>.W�E�hۂ!".4]���V�on���Zd&8�i�:²Z�?�s�K���|e��Ʒ��(����`Y�0����ݯ����[$mQ�?��}�Mw![̬��<���n������M�rQN���rR�c�(qt��Ly5bBe�;���!.K�\#*�fAA�.��j%@X#��/���	b�A�Z���t8�l�U����f&tw�f�ο�߸�Q>-��8ޏ=ql� �5gN�
�1���鐠_o����qT��G�8�.���D�Ct\~��'�D���rÖT�,q�HtP��� nn>O\b�^${��k�d�ƿ�͸AlH�99���O��=!���9��'�	�G�rm�e�(������7���X??{����ݤzg�4n�oZ�d�@l�_�E���3�鉬�t����e�?�4�b��Q�P����|�U�]%S$�C�����ҁ���!��ǝ�ڟ�~l��ls�kLi}�TxD�}���^ף�Ї˘���Eĥ�lta��"~·����Mi����t�lՌ���ɰ���A!�Sx:H�k��w�I�8ގ	n���k��C�"��٬�M�n��������a WR��Z��į(�x�^J���?atmi��D�$e'=G^Q+����7�]Sۧ���YS<�5��R����%u�	j��=��:a�"mR���Q���'�ϯ��).��-��ξ�&}A����{�v%f���(?��vo����o�� _�L�����4�|վR-�QD���#P�Q�	�v�N&�Gg������{s��֫q}Ev����b�I��y��Kϭ�蟣"�U�M�W��Y]|���I��NEɵ���-D���9��(;/�p��x ��{����}�Hc��, 芋n�Q��3�O
���~��34�b��Wr{�@��{���/�>ޡ� e����㽨�t�@��w*m���:�m��2�K;��)5 �?�	�j�A��grc	~
G��X�EW�w��|(���o�rd��8�G�&YH�H��G�nKN.��ќ������=,�?���J�Di���7=��ժJ���|������F�P������S��jiRѹ���<��lf�M7��Q�2�>�|+D�\rZ��'�?����I�9����E�&�g֋P����
�kK�Z!�Cd�_D�SŮDa����]�&�4�',�0`8�ٞ -]d��ǘ{��������.H5�D{�.�p�T>�߅~ܔ�����20?շY���>��3��N/ƿ�؁�����y��l'��mC!� l
�>ԴV�6T��#�� �"*矙 �?����w�B�5���i|����-o�����A0�7�o3�\�γC � \�3�����*���m1�,���oH[�N�:��Ӽb�6�j����Ȣ��3w?b��V%�\q�;�'��Z,*d�1tC�vMD��z�o6�]FUr#��>�]�P�7�$ ���x�hU4|2ZB�F�PS��4�����4�C�8��ʴ �r-�"���� �|Iq�.���rQG["q85Kf�{Gߦ�3�l���=��s �%V�� b����׍rL&�^6�.D>���1h�_^}@bYX�N�e��Ga�D�Ƒ�Z��=����=�M�Y�1�t1�^~l�lQj
b?u�8u��ܿ劰�ǁ^���y#�c��ӄ�蟥�B��b�XK�>}Kg�6=_���!D	�l��2�\��o�ϸ��Vۉx��$�����Os�6{���NQD0�$ڀ�BW���M��]��O'7 ƅ�
�Q��֛�+��^���0�GԳ3��Zrm�>��VӁR�������d��^&�0$N!�<�z;�`��5)�G<�1~W�5��*F?�� ��
�5�N��΃��a`^�4�uf=������6V*J���-:ᴔo��E�Ӄn��޹t��:��N8f��C�ꉼ�>�b��� '�
�K3eUW�r������K���:�һO�ܾ�@�Im�n�F��@ރ�|xD���Z��} ���/
Z2Z��-���<~ � ����y���m֯��#��o�u%��KyrD
��<4�y3߂�}.Ac>�����H��P�(
_��QA�-ss��t �{�� �;3rؒ]���ӵ~Wz�	�)���9fbr�dO����|`�Ld4uJ�U���cɜ�Í�D�[w�H(�_�7�g�#�rM�zl��@�#4��<�b��({�=�V�JNn�*��ֽ\���*�V�XKm��*Wd���ۣ��ӊ7�М�h�|�F!�Lpf�ow����MRh�dt�wJ�hY��1��3��e���GuIt����D0�E�c���n(g�F��������ų�V>�b�^���ةF��ϿoT�K`�U���PSh�R�ڄ	�4���������­H�w<����B���p�����s�[�&H�L���3�-k�#%���`(����ؾD�d}E�$+1�އ|����0ʓRe4Y��]�('b>�����wIQ6Jy�qXK�g��.���3T��_A�kJp��hyI/�ʥ�t��b�2)8'��9�;����m!w]����"��%'5��2�����N��j(?5ؼ����d=����a�?M�N�C�|�L��>��>*#�_3g|��
 ������)I�$ b� ����Z7�'�p)�{��b�,C-"�"Y�
M�߂d������@����b\n�0 Th"�>/��
�\N�����Xh�n�}<��6��\ċ���3�S>�O���BDZ��=`'��m���= T	��P'?bL�_;��)Y�Dn��,�m��Mx�*Sf/�l}j�N8�;�[�0b�M�4X���SA��H��iE��@��?��1���-�th=�,A�?V�w֖�o;/r�YeǠ��l؟��5���3����P.�3TA�����(�5bNֈ�b�̗ u6 sΥ��:=K��i��AC)] �s)9$�J��h����|�I"1�Q��y�<�������4��i�o�xv�����-J���]8����ǻ��w`�f�in���d�fZٮ���^W��8�}��E�۟(%�66�(C}����<n�J\���̷fz�ㄏFf6��>���x
L�+^e�����]_�i���v��t��1ٌ}�$U^�SH��]�c�HA@c@��lC��l���Ũ�R�f�L]��I�5�6�<7} $5�
v���X� �������)�����y|���3Y��OF��;�1=Mч������Jӱ%Q�p��ذPߓe-S�^��,$����I�f]0�E�{�����;�O6S�}<����\|}���-��W�N��?OM-�KO�x�$��-�;���]��-�ZY�L;d�r�ū���v�	;J���:	PF��.��Cऔk��e��>�hw]��F��p]Ab���{�[�	X�/�=QP�R$Q(tE"c�_��fY�mv�f��Gy�6�8�Gq�@t�jh�gNc���rh8�o�A�ϱc@�eo�p𹝦��vz��r���GC@��$�x"~P[��M6���])m�/��7FT�J�n�j�ߍO�Q�݇I�s͢ɷ]�ɏ�H�J],����.?�a�S�H��K��Ȼ��c#��T�yn�:59���oN7��~D�a����2�����̎�mw����x2ćKC�(��-� ���~�q������J.��?�^�XS�I~J�&����d~�����/�>����aH� ��AS�̯R��a���s-|�2����~Z�SG7桧��+˙�Gq��yጇL�8"5�����������i;�#WB�����6��6����H���ݿ�������v1Ud�K�G��[W�30�{W������;��z�M�B��j��6�Y��`S�Uf)����<5�Ӳ�ix�_K�G�"��`�s��0њ3�J�,�inᇩ,��C{$��r�'��2*iUR�Oy�����\k鴫xe�)&p�b� '�tr��{�T��M�c�"
�����]`�u)$������a��3���ٻu�$���`
��KMr����`\o��}�7X����pu)��f��#C�];s��?k!�WIm鷜lz�!"���Ѽ4NGwR��6;�ԕ��	
 ]��\#����N�f���˽?�lE�[��;�VzvE�g�9b����h_�#���@�QJ�E�l�Y#qRqr�'Z��B�ã?M�O�5��% ⠥B����:^X��_�]/s*,#d>����>W �X�ƞP�� H>D@��>�s[D_��u��W��8eY�D�Yr�b%G��:�� <V�����SRo�uE�ʈ�R^����$&�@Z�7΂Ѡg1:���?m	ɚ�v�6l*��L�O��z~�ƕ(�s�%��6�KaE��)4�enm�J)ݝA���L�����1�rK�㪬ȇ�� �2Y��j]���J�2�Ug��G-�V6�]���q�K�B<����sj�$���͈�5�>��{�Np�p�u��o��E@��.y<��)ѭ�\,gq;�`�I�Y6�%qgZ�d÷��x��(YUm@�<|ȣ M�*�8���}?ޗ#�W�̸�˂-%gفˮ�0��POdl��|U)[�)r��g+����d��Y���*�68^$+�5�Hj���h���W�3�jJ�ɝ�H��x��=�X^�F乸7�Jq�W��_��C|�E��Q�S[Gz�"c�TKr0r��ei3A{�#�鞴!΁?�#�p�^⋩?�\x���1�'��y����{���Jc��J�埵8��M�)���	�$��o�V��'��50��ڵw�5��\`�[��Z���r�#O���'2��iC�+1S�uJm�S�N���RxgC�p��;��P���it�x3o �2$ol�pF�DW����&-gcH�����/PI$��J�������!�L��<����w�5#���5\��$Ug�#��̀��d�<d64��Y��Aӡ̷>ZI��Lv����Nwy�0�i*6�N٨I!"�-��<>g����c����5"��R8qB��s���~�6���Ɏ�u��@�PQဖ�̗�G7e�Gvb;�L2<���H�������ݓ?m�%��H�,<�ke���Gˇ���+*��S|H��
��X.緽�Z�d6��D(��:m�!���}��t��Z�b�s?E�7!_��d����b^x=���AA�1pMQ���c�۶��c���V�8�����2
�/��H
����j�ԍ���p��$t�n��Y��i3����)���Y��a�����w�	Ƴk��V׽S#p���/����\�r��:�BpO<�[�����x�%���zSLU��p�T��)��%��d�����M�����W�e��LJUU���S�c��"�4Vgt��D���z�@)���A�M���v��8�,���n�u�����EP���v�|��?4}�6 ��������bF��?dַɮ�Fύ��=���|�;�t�J ��O���l]59����ڃ��I�a���NDgA?ubp$�MC���5Byl�L�F�2��t����&%-�%>��� �J��g��];�ƛmؤ��]"�����wd�6.����5%6,$!Y�iʿ�C\M�S��.�q}��9��(
yO8��"��FJ+��=Qoi7\�+��mۻ|�v��} YQ���wa�5��};����>%m�~�G3�8dE4�>�N��Ck��_��׊.�L��M�DF�`�dJV7a�N�
����0��:��CB]�<�$���A ߈�z����v�M��Cظ~Cx���D�Y������-�N�&�V����c�9���#�ΰ���%��,�ϋ�!k��x�����p���� u�ռ@̑����WS���v����́��Te���=�i��U���ΰ����l�zf��3��mG]֣#E*"O�������ޒJ���7���2
��=H��(�M�ӟ�m��교�70�D?������� A�+�#�o�¶I�]�9�R���);D}C�_֦�d;�u:5";&c�3�H��I�'<4	���6�����)�?y�QS�����L�CCu�D�i�N�`^��Y��H{ӛ���.�셱t�K�҄��a�p�Ny�^�:̵e��ˁ`W9�Ϗ��XY���$
'���h��ӈW���S���:N?��X�~���C1��	 ր�1����'KJF�@���e�HV�'p��i��6$��\0����9$����X3�AFs<^@�F�>M(f�o,L#-��A��45�@~.�tڨIȶڅ�������n�H�Ű#��!>GB�؛)b kIE�;��0�A�/ɐ?�h̲�i��h�t������һ�Nv��o�6!�L���������\�?�Yo��#ێh1n6���b�k��Y�m������,;��Xz96X�=��������[(�1�h���?ƀ���=�Oil'?���J`��t�|�Q��x�8���xǲn�JCtt%E����~��*��w��U�T.����~ٱf��dTaǓqp��
������� @C�2論y�,s�ԞjT����u�Fp�3�"Wt��^U�LhQ�W�C���Ҝ�SyHq�ۯ߲M}86㷞�n��iM�J �ߐP"~}����������TMRj��̃@F!?B�9�ck�q���X+0;/�x�����&�MP./�dAȟuh������?�Zj���iYx$U��$Md��X�F�L³^-x�GZY��Y5��(����H�{U�Ιh�+�Ah-7��W2'�$l�
7���P�{vc!���bqr�l���Gq�Gr�4�J���z�̏��z�Eit�&��~al�4�-�4����|~�v�"��",c�ɉ$I!T�&��ƀO�ğP�)��,MF(��`Оv��K�F�������*�
d�Qjn������0pU�u�#F�+���$�k�vH�eo�^O!�Q��7,
���8�8����/�ԶG)�{�x�o���
��}�,�xΝG�3u,����y��Tw:-Eaۮu�dm�	�����i���j�8p��$A�����&eEY��f�c�)4l���kļ%C�-E��ɗ�kOh�ytQ���k���|!��eH{�D{�7��s*����q�"I����*��\빖�17D'��4��u�
z��-�Է����˂��8��'�lw_M�E��0���}J1�X�.�/q�dc4�"��[Ye�3U�X8?6���?V��	�s�g��=ԫB{A\iYv���(Pw�4���~�q�+un�3��Q��C|V<V+sy��G?S�a�p��\~n&>�����W��$<��գ՘��