��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\���V�fnvx��ÍG_;�ȅe�~�>���9�>��Y;�0GP�5����ȳ����#�����Ѻ��VnJjv�y1!�;��������}C 	��vqq�����mp��*����t[�K~7�d�|�k��d�3�ϩ�#w ��p���>�փ��S�3�Y�ҋ�{��
��1��TRpn��&A���ܐ�Q��P@C'�CH��3y�6Ҝ���'����� hh�cg*>�%Q*
m�ؠ����ԓ��p�_lq�K��Ϫ��E��kh�V<�O��+�M�ͥ#�1���Z.%����q��p_�~&�3�@�dG|ۇ�{udG��I�(�r���J����o�s6�Ä���QO����?��ی��Aƺ�Ou��dB�`�wm�B�/%j���C��T��­�[��d�a��B0�Z@���Q%�J�{_��l����D���(D��Jxo�='̪��~�׶j�J�j��S*	01� ���ʞq�����������Ƣ�u���!���ln�
h�4���� X��t�q�C��h�֡u����XHJ{��h�|�Lѻ�g�����cs�B"αRzx�S�&��_�F�S�}6�����u)�{�X�h�Qa�4ު(hem�4�BbR���<²_'���93nlيe��r�B*םUu�fr��
�#���4�`�p�^&�0;C5Ղ��`��@�����Sz1mC�U�������ӑmu��w5(6C�����%�̒�\vNx�>؃ݾË�5e��9W���vЅ��I��T��D�Λ�$+������-���V�h�N
�'gm^PY�(c��`Ⱥ�zO�ò��*�lw��W�_���p�B�.K���^��,-k���Kh����@�� έ�2Ϥ��a����mC|�A�s�xG|�9�7_;�K ���	�����1Ek��@(� �a�"xI�a�!-4!�\�S�N���9[3�MT�e����M������+�÷��"���������RvEm�q$���:w|W�l*�8�Yڃ�Q?�Xꩥ{D1�=��I��(�:60�LoL*����-J ���Ǐ �ْ�c�Y�y3��lV~%�Ui@�咆�*��W ��؉E���F�nr�4��3*\:@�@ҳ��	�0wǖ��;���\�^�����.�AU��`�ԫHPY0��}�=G��B-fa�:LgU?���,��	�CQRfҁ��/M�/�Q���$�vt����1P/|/�o���?�!P)��������.|�p��Pr
be�U�м3�����K`ru�-?X�T�����b�׺��	�'6���HȠ�G��ط�b3���ߨ�������B�ΨY��]'~�Q����@���
���A�6K�{�N3��+#��*bN�(�P��C@�;�ctE�V�����;o�=�Y��i)��FS���G�bc�)$����
�9��V�����J��߀�P���H
|�(7I�k�5��;����Ӏ����*�Q���Q����`(!�>�$���%����Ee������-�ʋ�I}'3ڌy#�oıU�L31hiq�#���X5j������TsNs�n6=��閎<S?.s��,?�Wۄ�q�����{�]A'_y�Ľ�B\W��%����1���k���l�h��6�}��	μTCgd�uc�h�J~�ҵ!���kR��7��3��M-n���x[��('��q	-��u�Š�,� xΓ�H�S[�0#�&?N���.-�����'��9�B�?6�DX��[����ʿh� ���Uf��x9��d�y�Kn���L���k0.���^���/�f��LB�N�mj�x������R�{���
7�kj�C�\n�RM]D.7V\e�1��ÍQ����pv�`�1������a���M;�k�d�S�c���׷i]꬇D���?,��Y�b����;_o��z����ê�2< �t �\�	sZ:46�9G��
ѹn5�#��&G�9��9�iC�}O���c��Y=����!X%���	���r[�U��84�J�.?�w�G���#t�:�i��3?�Ll*V��$&$��ɬ/��o�8_tn��ۢ�C�M���pN�S���KÊL�g�'��\��H*P�ͨ��2�a ����`�oŗ�+$��gs~
��`�/���{+(��F�6M������Lw?c�O+��X��Y�hXv��m��:z�J�C)��eڈO/Ϣ�)8�� ��w��l0�����q�#��n������(b``��N}tה��rop���W�I�֬?���X2,q�g�uu����?��'��i���y�7w��u ~�a��8��v�JsB�" ��o�۬�Yx8��6ho�fp�z:�tB��]C+[~��љЗj�p@�ێ	�x̀�	���J;~-R��X�{�I�L�I
+�ZfI��g�zIH�=	��H�  �A 0n �G��$;�����#!�4ŭ]�F�4��}�V�qt:s���P�����OX����V!CI���;��/c�K\����N��as�phr����vqz�\�c���Z �Ѡ�_w՛��d'M'6��!k��<h�F �|j�$LD0�s�{[��oe�,CP����+:~	~T��x)�N��ñ�!����)G���bǝ��y�}QÐ�jvﰑ^�9BZ�:��tQ�n;a�93��o��Q��|��ܒ�3f�/�-��F�H��d��L[�2j��㶅�#�x�9��p=�/�}�����g'��|d՛)�z���7���@HS�`gT0��z³����#�{Z�� l)�c�L��-��lL'gb�+������A��5�8<KֲѲ:���R���G�}����4^�20�!gE2�n�۹���J�AY(5w8�5��������<���KSy���D��8t�"8�.�Ւ�eq�C�Uz�I�����O� ��c�'z�������.~[8�Y���'n�I�%A�Nxt�~:?s_V���+�����+:�]Z�O��-4�%;��|�$H�kC���h�?�;smꑙ�� =�0���j�?��Z����1�>�6+~I:�c�ZBB�k��QnzV��Bw4����^ϬY���Ms�y|�8�M݁0�ɍww�~�����sv��k�R�x0/,��nD��x�c�)���$u�M���礑��G�5�i��֧3Ljߔ�F,�\�WF�I����Z��w��j��þ��KFI�ٮR�N����e���l6�R�l��E���{I�䴼��^xrEM�V�=�!c��_n�I"K-�#[�����{�(�;AΠ.�| �t�?����c%�,m����f���S�7���|�2IԼ5&��pI�FQ�����[���+W�*y�/M�X�2��R�*pk���K8���CIg���M�rO���@¯��4{�*i�;0�7ر�0�.��p!����gF��}NNTTx?�*��eh�"g�j3j�QO�BkM�Z����Uw����{�R@�F6���e�A�.�%0-�fk����N2�s��dkG3O�t�p31'�o���&�͈��L��6f����IM*��F�Ӷ(¾-�泤���Ahڊ�x���x�f3��7�?�9������?�)�@��X�X9��-�E�����}�+1��n�Jw��*f!{���tO�YwӸ��,�ww&���-�G�f=;����?<�:���q`���y�' �\>�r]�㩥��.[x6�����U^�l��ԃ�)�١:!?֥J|�K�c��N9�9�������'�jA�y��ܱ�R
%��Ԕ���0�rڨ{p�8�J�z��Օک����>��������m[E-�K�xV�~[��^��RN���E�O�;�\~�S	�|�#�1�N���)򜷙��q��9}�����԰�\n�2��B�X�y?�ۢ�j/�"<���P�����%����!}C��Ѡa5��=+u���Sg�t4)����gib0��͌�Gu-(� �����9q(���:���>�8�
�e'>ţW�J�{��AYr�,�^P�g8L@�����y�p�*�[Ҭ�w}�9rth�j������1�*a�U�^}�\W��b���b���d�<م���s�V6���8��ށ�tF�׌�bL���H��%t̜���}3���g|��z�4���s	�r�j�i2\�rG�4;���3�����3\�@&[ dŚ����Ծ)v����Ĝ��3|h��%��Ne: ¶��!?�J�z�֍��$��F1��m�TL�C3��"��3qA�	�7��/q%�i��X�$H�|ʴ�<���eG�uwW�B�p��X���y�t�6�)�7� }E�rr�j�&����Ѽ���3"��b)�tIF���s}���	F�j0�)�-��!L �A?�(�6��0.���V�����BB#q�^�Ê�j�϶ 6����Д�����Sk�{c���`B�5ݲ���ZR����I���H�9��K%�5`҆5���Տ0۪�>&VA�r0��XڇOT��z��=�C��U9�S�t��ju��$���InRzu	�G�Q��g��j	v���Ɋum�� ���
>H�{+�*f�b"�Y���mj��l�3�^R�OF�����$��<s�	N��t�M�������
|~��ׅ��O�g��|��oh��Xr� �H� �������#,��G���z����avc�
�FF��h���n�jg�:�^�°$Y���	j�^����4_��:�f��Y|#�s�;�<&��&[\�nz�y�O�M�DH�4��\�$0>V��N*2�
��[~$�B�E~ӿ餚�r/�WH��''�=1�����ZIQd������p�"��{�؞y4B����~�b���3�ou�_�[�� �֭Ae�Y� ��Q��G�~���������7!�O`�|;1�t�-h�?푻"��m�g��jƆk ��b�&�+�@iq�9T��s>����oK*�m�-{#*�4��_Iu�:֚aӍu3��<%�A6'�>�O�;�sU�`K���0����t}N>��Nɑt�2>�4s
��?�!�?�҆�٠��N�t����P������"F�j,>�ǻ� ���e��S�#��!B Q�~�7*{�`2;jO��p�忪�#s��c�uv��?���]s4����PzWV�:�=���\+ LOl������V;|
�_����VR�pƝD���b։�6:/�)�m��i7Y�s�+q����X�>}q,v�����WE�����W�-�$l�t��Fh_�����}l������;�88��֮�rK�pT����D�Ę,^Uy�K�P	�� �P�y{J����.������@�'��e:�I3	xTi���7��>P`v��ZV�\�ݟmKt��o�l�L2lB�M��c���2��K0�֚�>���k_\9;���ht�L��ưG[6��s��;i��ym$�A�08?��HQ{�f�!�N�<颾���ݻ)��86SE&U^�+���0d52V�`�	��R��AG0���l��XO�ܷ�Om���f��� ���Sjb�)7�P]�߿N����˒����F� Od�?�D`c��@����%�C[�S�` �6r y�.g6:R�L�ta��"C'��ߑ�q�]u�۫m䃒q�C�
ʦ���G�"N����h_S� ��4[]韜��B(PK��I�*��P��x�S��:v.��T���u���u���LP��Z��9=��n�i�2s����v�3�4Q�0�d��C`��_���̂]������?+:���T�)�Ջ�I��"�ߓ��b�U��d���SϤ�Q��З4�rMNR(�rs��!��+��1�!uYj�\�w2�}iCy �G�d6�<��P��4���Yp�����ᗣ�<�gœi��/�j��@ݞ
]��t�ی��ӛb��=���ڄ�;NT=����t�qp��'#�e������<���Y�����/|�'8YW�8MX��-p�T;��"SH��7�]��q)���)tca���1������j	�o�������2�_�#rq!�ɸZ�������È��:Z��RYc�:x'���)�."��<x{Z�`M�(7٩�z�F)��
Z��c��h>��e4�.�y�ZO}�:�����I�z�[j[g��>	#l�.d�oK�x���m7�Z��$gi�
��6UI�O�#~uj�� T@�&�VU#0(�;�_v�Ic�����\x(I(������N�s���Ȣǰ���4� `�?�r�V��վ��^FY�g�b��SQͭ�'|�}���K�ƺpM܁0���΍�v$m*؍�<�&�foXT��2f��}�-E�q�"�w�B]ϭ�����h���@ژ���v`�+2��4s=+����v�\����?�.�%�*�OZ7�%��_�blF#���;8y�r�|��-�G�W~�u+a��a]�%e���-�Ɓ(}�P�/׼v�XU�iI �!I��\&I�_)�q����[3�D%��7�q��YtƆ������;߶�Ox�{��Ի>�F~>'���jtc���	z���Į>`Q]������>�M�#���2x�}���z� ��bQ�߁���v�ͮ�|ޮ�4���"1V�=X�虜!��/��״1s�WX�R
���F��,���4��!*i���za��,e��T g��S��ܨi�]��@�`h����R
����[*.��,��Ɣ76 �m1Q���P�������gF��Q�خ&�f������WsHVdA��!_C�@z)<�F��dKdE�����[�9�J(�0py�+��=�����,���bz�����^��<���r�N5|���_`mL��.�{��vQ�33�VRG�)2���x%̋�o�Zw��n�5�F��q=n޵�K?��OG�m*PǌH�;��hm�B��x�����Qn�[:L�O�L?Nw�"Ƙ{�py�t�`��n���yA��`�*P:�^7q�(�9i?��B�QƩ�b�nnE9�z�I	�fr|�b�V�t��N�sQb�V�3m�l�UDVH��8���Ű�� ���˨�E����Ƃ�2jЩ����49M�ߐ:tG'���(^h�v��,�gCV����D��1���� 7�L:�O� ��B�1.���q>�۴��YaƋ�,�%�����+�z^��������F���,����I�����YD�M2|���<�r�u����������X�d��%��/�eޘ/Kc~�_gkb�Z�VV�yA���6:f����ה�'|?V��P�f:��g�V��Y5���.6�^�j+W"s�������!��a���2
���G7��(ka0uAm�Y����Ѷ���֯��2Ƴ��S`�.v"TT>���Ʃ�c6'i�}�oyNMs�瘆t��Va�,�6{�X9Ԛ1�6�b�Â ��Jb�F�'��Jiw��>�7����g�,�|}�t��Ĵ���E��GG� )P�#:S[%O�J��J�I���{ze9!"4���@��a�*�mZ����d����3w�?i��,�7`�aM�T&?�ܡ�.2ث��A�u^�SeX��v��'�&6��^)&u1��؈���Ʈ>+ �������)���=�E�G1��<ԡ.��h���9H��~JV�2���J;𤆐��S��{�e<��O�L4�І� ������K�c���&<�Q����
��F*��K�삋$V��I�r�]$P��.�'���J2�M$`)k�>���_�	OSj���^�~W���ѡ������ɥU�)�,	����۠���.��V��-��p��`�%v��xd]����X|�<���+l�<�jY}e�]8s� �'6����(E�:�vF,��]�ﱋ����	 ���d��[/���3R�Mty9�����^����>"&��sY��>��j��`0�oC���2� _4�ho��:[^���p0�8���N��vm���!�q��'�61`�͸�=D���9�cD�#��_�&`�o��v�֔xP�[o�Ct5��R����m�=d��ܥ(��m�ZpRma���� f����{B�>�PD��$�K�]�x/Y���C� :Ɂr*h��7��7�]X^)߈��Ԏ
g�u�l� C?�[c����6��΅�жy3d�~��z�Y�S��7Ĭ�ac�P�Jұ��D�Dr�_��W�(nU���@u�P>�~͡U��Y�����T���R)�}��4���.��L'	�~!�7�� ����=�sD��|�	��4ķy6x��D�a�9�RJK���\]jzߟd��0��k��-"�p%���bZ�$�y݂�D2�����e�3#"nicY����c!+GXI����Od�f����#�J�ن��o�K*���|�['[�-F��6�ڸ��$Tv���%%����4�����IU�(�C�I��<�?tЦV�hn �Fòz��Ӧ�F�v��.������ݟ�ذ���>%!e
���
������b@�I��;u�템��9�moO�kA��9�|�t`}=����")�Y}���8���4�pr@T��4zJΡ;W/oe����$�Ē����Oi:���B�p�h���T�c�2�,��bהv^�Q8�9��mᔌ�v�E[�q�<K����t���Y�3�>}� Q^������˞��3���;6��z��!�j�T�r"�+Vks`�IO�A8���&
Uj�P^��Z~�Ksp��>�DÎ�3.�\�����X��d	㳮P�y,!B1l���CR*��{he�ַ����#�>l�Sa�<:���|�ࢻ9��)!+Ƥ"���Xͦ�j n�>
m*�P�Gΰ�4��u��5�P����?�:=8�_fM�����y�Y,�������P�4/���g`=�ڕ9��=�!쥣4�&�E�dU�cL�G�BkIf ^�a�H^��BGOh��ԛ �*{��cgk�1{B_�\��D������!���n���Q��qw��!�Pm�����|196�t骙����m$F!�ɷvyʰ*a�l-�i� gm�!f�<b�����V�2�|J��	�JYj�B�OF MW�~��[WC��F6,B����k�O`�33��Y���M�}��忡 
�o�Ns��_W)'�ޓ)��q�o�n�Mq,ڜ�0w�7$Iy|&F-�֥!�MP�5O>�Jm�#~��W�����Q��~䏂�3���f!Z�i��UI�ܮX�w�>�֢�1�?�-��ChR�`
�!F��4і����k��Ys�b�_݃�^�ă��^0o�`aBm��%u��9�3Tg���Q��9�Z�#^ ����P�mu�7y�.�����{?�G������
'���u��z�2(��$;T����X��OW�+���f��^MU�*�x�.��:ahtZ:mI�.�5W�}lA��=2H¾�@�?��YQ'!��h��%��AL��1[�+�x�?�,!6GͬyIK���=�*k�h��[�t�D~6� ��2_��{a��):�%5��']�`��f>+u�gW���i��t3b�_��6���#)5xi��s���w�/��=Ww��yR�5�^�1��
��U��f�j�VJ�󎡂D���Sxt��1�,E����1�2�_�4�v���ǂ1;봶F���8�I(��H@I�͹3��
^���K�����R�;=t3gl����:2��v�FK�>�(���я�V�Ĳ���D���z8���"��x$�:�_��HM���i2P�����>��K96]}�]0��	�l�h��9�*���+�bqi��P+ke��������ջi`!�qOp�ˌ-#lev��Ձ��yy+�U[v����Zۏ5ڸ��4l���|3�":LM"Y�5��fx�X	[T�<���I��:�v����F���2�~�2p�"���{�ܿ}1�_կ��BQ���Q�Nb��ko2	�'�F��N�������0�@�+^�Of��j��^[uyC��	�^��I [4�a0�����Ax�Ak=G����ȩ��[��w!tAa������
i��n�t>q�Φ�j��_�cy�]�P�zX�
:P	�����w�2'���79����]5�p�(,���'X��!~M9�ؙg���G^xf����;��=h��9|�>����ڏIyk�1�6��Дw�aM���WV���3R�jN3=�3�e��2�؊��l ��	 �=��Wu�$�.��[�����<S94�c�?���-'!v�4z������+w
#WE�yhZ�m�ʟ'��Cg�*�5G)]s�3A�N��"T���%��?���6���6rb���
�������$uE��0�[��/�}jO��8^q	�	5���_)۱�_K��ަ��N�&ى���v�r^�`�d>�2'�B =������� �?���Yf�Tk��1������:�0#U��X.2iK˱���k�ߓ]��� ��Ⳋ���˃E\�=�1?���U�$O���F	��9aTT���T��I?*���yގ"f]�Ƒ�R)I��{�W�`�2@E�#O��E�9�����vx`%/Ʋ� ���o f����w��U�����?rv�Q��Y����B8,,f��9��~ZN���n����HᰮJɧ�4�*^�h���W9z��c����uX�(�'yS�!@K�5S�:�(Y��v���)E����Y�:��Ȕ�ڵ�<�Ơ���C��qEq����oxW�m�ʇ�mFmZ�"���V]�����)K%+=����5���i�{�A�놙}�DuA#n5ٰ�Y�q`��e}�S�^���<�n�_���̊8��n_���cS���a��>�]�pA���Fҿ&F�#C5���>P#B/�)�����F+
,�դ[��4Q]�Q�Bx ���֒ f]641�(8P	�ڗ�2Zo�A�~��!�)�3�ՋNF��eE����}��t��\rR��m%z����bC:��ǅ�