��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\���V�fnvx��ÍG_;�ȅe�~�>���9�>��Y;�0Ga�%m郵�Z;R[_��cJ��j�F�l_����.I6Y�%b?�ʇ��8�1�?i�~?u�E�=���9�I��[dҍN^y�h%0����/��JTmWrmw�-�١��*�h8�r�8]�M�p7��l[p%Z����n�����+֙n9k�[����l|8�I��ºQ��q�7���<�-)�R_�MF'����1~.�!��8:/t�b5O��/P%9��t��Ai1n~n�q0Z�G-��S++�m���:C�m82`w����F�%�SKkI8w��u��5{� �Ey|-����DTL}�4���j�Ġ��_�)1������������'�}�\���܂NGZ�k�hx
G�6�C>-�K�B���vZ@ۨ���g���ڕǑ^���*g����)�Y�q	Y?m3�L��\�fKz�S���v�m��6�{`�m%L��/�c�����?�Y�=f���&�+ �,��	�+\����e�l��`���U��~��J��u����P�rFœ�`�~"��1�{YR7D֊�ߌ䞲�����E,�[T��cَ(6�����Q�[��	�t]�rT��d���鴗ꄲ�G���r9:�~O��j�Y�u�˦�T�M����e��k����.�e5�sxKE1�ȤO���U>Y����t���.k���xc%�o���>�A��2�~�G�9_�K�b�G�6�]��1'�K���MI[��9�¾��tS!!�%$�Jg}i���M����6<>�6k�Ě�:���0��Ǽ�W�^�}�A�����V����@=�7�%"�MN4��~?S��tt�{=�֢��F�w�Q�2��AmYe0I�W�$�.}�3���$�QQh}�s�#����M��L���'�~��x�)�W4ȟ����2��)(3�{U9�y1�Z���(�����fY[��.��x�x��[�Y_E�y��]��!� \
H�Ov�Z��ф�x�}��}X�(t�1��8Y���
���8�=�q	����\�n̼��E��ݹnE�.1�H��I�a@�+P�Ӛ����%x�4U��r�!��S�<�2��0��]T�v�d$c1�Vl�-��z��7�޶���Mݽ'��ǭ�`��Qd��դK�t�^s����[Q�(qW�ɗ���X�3���u4�0\4L�|��rZӦ�Ⱥ�K�� 4�s6�����wŚp�D��;�"��슐�!J�ޖrp^:�^V�D}5 Bf<��>[�I��f�=�˰��ZU*���O��k��(������K������M��F�f���n���qh%��_����)u���{���2x�5�:/K-�E�(��6�_��O��ڝ�ϵ ��=�+���� l"��R��V俵aP�Zܮ��ރtX��~������2%�s!�NPX^��9�5��������Y��R��4�iCLf��wj�2�C3�#u��|�;R;:����?c���� S7E.H	�T ���o��Α {Tc&~�u��]e�jx��>U���+�Z��^>k�
���۝��S�����	RR�hN,��,m�f��M^��{��Y�&��� �o��lNu��i;a�����hP���/��� �NݐE�|�M]�SBo�l�p��ɻ?�ZE�Ȇp���3̊��K~"^M�j���p/D�ZhOQ����ZXFD�KK0����аo�^(�5�j�k61�W�o�s���R=�+,Z�����%����5�*vQ ^E�O&U]J'w80`���/��`b���ȶ��]���k㽦Y���0:��my4U�Q�4�W ��s��,���55A���������'��z�F�>�A�|g�@E�#�p}7%�EQ�C�r��� ȑ�%>�NW�����39�ę/v�_����q|������I��i���.��쏙��R��=;��Y����vj�J�ST�>�뽇Q�R���Q:�jV��!�9Z�&|&�&��jQLg��/Ϸdy>��yf�I�$����A����݁�i�_�����j͈���h��!sA%�_�=f�=9�sINy��qM��+z"�#[�k�@z�ϖ3�� xg��e�h����8���w��B��RXX�/t�mY�`t0�[�Ɛ�e9�e	�@�T�J{J��j+��,�~J�ٮh-e�m�e��đ���6,�@ğs���;�W:f���=
��'sdJ��5߱x;��%�U�� ������� 
:@Z��X-�O޿��Pr&*hȹ�*����V�x7|i̤��o9<Ac��(=J�����P3I6'K�A�f_����ފx�*IX8� c&db�4<ix��R_��5_��LN�^V��(�Oܻ-��H�>2������F4Ie���s�qZ�*zi��bFU�0U��t����C|�Y�G��;q��ۑ�,c8����������a^_?�Lb �����g	�ƹY�`�-�0/��o7��7�(�Q��9)��$���
���$m����rc�Oů�9������}�N[���/K7+�%��.��7n<HL1&�,J3L���`�7�Z���
���LM�5�*]��[�ȯ�;�<�a)�訍z��� �s.x�0d��fF�j��um��f���)κ���e	��i*᧓���N�`�BB�O���:��yR~>˫r.&�#s��A��df�l��$�O������G�޶���y�+Q@W�)��G�J������A��I�jL�����ڷ�iQ�c>ñG�|����E��G��/\��>LI&�J|��D��Ƀ���SA�fU-G��/�|��,mq�݉0��_@|��'|x��q�~�rqB��G��K� ������edBB�ԃ]{�$�;�,�Ũ����!���F{���6�gIn��<H�����Q�ck�7�A���'�q��69��@�S���z��č����Y�8#��Î���0��D��-���G��LP^�97RU����X���=��%�֕�M�q�T��o�(w��J	�s�Ӧ�1F�3����^Y���l���OD7q3�ߓf.�B��:tc;{��{��m������^���t�~�C���K/,��~��-���FS{�P���Lu!��o���M�?�F�L{T��HQ�n+";�� J_�����`+��!c?{D7�_Q�*
�7C5L
�'��ۏ�A���Oj��m-)i�c�ZT�0���	��"��|Zl��[�h�j�;C��:�MI?�f�6�L�'�P���V`��u�%]r��Ku�/��Š�j�t��]ۥ��d	5<o�~�SH�T[��n'�3I0�G�8)���n�R�J`������0�n�������h=�(���������0X^I��!�u�̀����0�9�G�e-��?^�x<U�a�����G�4Kfq�ޔ�Tn��%Ʃ;%� �3�khi�r���OC73-►{�|�!�7�X�>�]�%̈́h�����'�;�/D��tw�'r)�v�������%�Q#�,�S�e��/3��Q^w�AY�GR�
eYi��y>�]�l�\�`<\��VP����xq�W�vP��I?0n���+���&;:)~ʕ�\��qٻ���pR��D\��O��\������(	��~����8�(F��Cav�jw�c��\_�,��}azCx���S���k�W�˅�l��f�6�SLzbP�������~~D���@c(����A���Cڹ������C��ޘo}� .#e�1�g�f���;��R�X�~-4p�E}��Fш:/��q�oY��b�s��U]�������S�����p�ħ���<]�n��.�*Pτ!�Ԟ���a���(�}z�o�8��G|�=@��4�*�FCl�&S��W�,�������7��%W-��m�Z
\$�'�D��!�b�Y|j;���>L^�E|��W	-z~��o��`�Q�ƒ���f�_Ng/n�Q)�����\�o�q���0fF���f�Ô�}E�P�g�0�VKnJ0n3�et��f�2����/�K(��[y�k-*�"m
��
���A��!���)��^G��V���3�ȟ��gۼ��j!�Og\A};MLǈZa=P�y����2���Tues8da���������^���V�n-�)�^��O:`nnB��ް�nU�m�����9�|C�aOQ8qf���_m�Z�ɶ|B�щZ�s(ݾ��aG��!T�I6�X��)��b����'"�'��)C�:�?4Sm\���&��
M$?��W�ܺ!�A)r�;���[���XE�q 9õܐ�3{����}�ŀ؎�����c�k�	t�-~���cNk_`g b�'i�N띞��cA�~�/^�>�R�r����պ!Ӟ�ݢG�� C7L�O)�`��B���Q�g��a�h��W�"CD�#�d�BC����0�:����M��_�
tQC����Zaa���4�SF���$$������&��Z������z�ݴ���Ȫ:���v��Q����ao�S2���B��+�����&X.� �|�2�|��	9��f��Xfg�����8v-
OE�n�f읢mf��FE�en��?5��)]ي�h@<"慃��Uaj��G8C�yw���;�6�fo���d0Gaa�>����җ�_M
Ƙ�H.��K�/_ܾ�HZ�_�Ib����WN��0�TP;�CW����Xa��V�r�J�U�hE�6l�;���L' �b�/l�͉9ǽAI}���Ӳ��6�߀r%�-�*G������#*�{��>�j�Y�5Q*~j >����Eѣ:�A�!VU�x��"2!A]�)߳J�@c,��Q-�����e����!?�])�p�H�{�Q��=��^�.W:HQ�4ɍaKXr��$�����%�c�DS��D~&�����ɦ���v�{v�}���Y��f��>��=s;�͆1QrQ�t��B�ڣ������<ts��� �C � [	�
W�\!|w�V��Q�m_��|� ����)��fa"f=�A� 1�Y�-�-�Q��r��h+ފ�j-�D,uD��b�?D���à��
�TU�E��rnC�!#RG��#L��V
�rA^G?��i�Dt�|V\��&�!3�)�	�u�[��<y�ǡ���3KF��Ub�~LX9�
�p_�a�@j����YxS]t[���<�w�B������h����^�glI��ꥯ1��B��]�Eb�*�t�-�eD`�{?aYg�yp�m�+DT��)�+�jғF�8(���οA���>č8x�V"���C9�yb՛̳һل��3b�3�������J�����u���Wiq��	��%�G��J�k��ʧ����Z�����Vy�	d�:��ՠ�(�%3���[��Aa�9�ѱ�7a ���3ƗEsEZ��\�\���v\�i�bħ�E[n?Aw�Q����;Z¦Q�}�>8%�φN��nUyV��$O��U[��.�f.�W��u�?��q���1��a�'ul�>n9�C^�cK���ז�e�^ؼ�Gߎ���8��!.Hu�[��j���HyТ�F�����|�<D#��Kش�5/�JeߩIS��vW�Sܪ3����u5��H,\��z捉-����ujA�O�G<�Vz� �8bj�{��V.�� !~^�`_ �~��|�$��|�Z-a"�-v�R1��x�J:�G��'�y�a|��$��i:��rir�]��o��,$��9��������\�໅����$�^�CN]Q�R��P�!��\��Ȋ^iA_$R��l������U���Z)t�#�׎���\�,=�ŝ�U��p}~Ψ��Ρ�O��Ȑr�g�@��X�Z�1(�@3���3EL�����t�<?�:S�@����((����o���t��$W���)��r��5t�"0pB�({$�X���
ͨs;��L��vbfdI.�5�刌��I0"6�a��	>�Q��8JV%[%n��3���}������~b���P��i�[/�Wqb��C{��K�iݶ�Hܮ�D�z�|��&�I���^�e5�jMJѽ\w�������^iqd���������H���_݌Ǣ�2.u��-��7��=�B�"i+�E������]��.YJ�,j�ol�-o�j|	|��5ౌ e�ꋇ�?i(�1����/p<�wȲ�1\��Ӈ3�9�+rz:����^��7UERC�����tBi����K|��'Ŷ�.)��F�aj�]�HѢN�r���9�m0X�;�^��L�d{��Δ���N�i	��8�����5���H��p߄V� &���RW�	/�m�-V1Y݉K5�]�l��m�i�ԫIU�q!n�i��I��R��[wj�#�\�?�,�^�T� ��^^�	������d�Oˣ�9w��`5�<�}6�$O���r]�]_��i�n�ԕ�p.��!>Z��֞$휟��=�mht�Y�dݒ�c)��=�4{��~Ф=eMG�3ؼ�q����q�r9�	�k�Y��Y���GW?����g^��Sw|��n)H���J�q��)�����M���Zȧ`�+�fz��X1₋׽W�����)�"��E�!����/Df����k��Z���z(����d�F��P�:��;�����Y���טH���n��_�w�iA�ö~ooͼ����;N��SA�te���M��ݗ�j�D��ҭr �;_)umm=����0F*��|�As���
�WBz��O���G�Y����'�}�pN��rC�	sRX-VX����U��jhU�aT|6�'���t��!��I�(/S`ň��YQ���~����AV�-�ి���?�.���̒#	�����wDO��|��xk��܌�K��0Y��Z���C��FvnN.�1g���(c=�|��B�P�}�����B����CL��r��c��%7h��*�d�(|8�ߘq	�/�'��2*�-UI�3�XX���}ݤ�"�� �1-����1y9����x�>�o��W�)T�'2��AK�`d�N	��,�����]M>I����ʕ�	y=%M��g�G���k�vY�P߅exPOl�K����\T?��`��w���:]��XhP�����)0o�	7���ό��1��ܒ��7_ �DB>�x�Fr!�CD��y�A���2���ٹ��!I�?�1nG��U1�y!�]�5���U�C���U3+��?���ѫ�s#6{��Ag#�Ia��[Nq6y�h�����Eʺ5{��Oӵ���sB~�}͞�Ѩ&�����S�m�1��ٖ4,ߟ_e�C��S����.4Z-;zV�� 2�cjk杇�.w<{"���H�*�Km�B�����U��͓�@�1�ʨ,� �-�DUc�Rx�4��tǣ��^v�s��g�j��/L�%��$��ϊ@س�]X�A9��y!D5��S���<�I�t��dMO8�:m�藾�fP�6�������40���k�k-� jPv �S��%	0�1�-jcr�(XD1�mӐs�p{6����Ӏ�~���QN���4a�q;C3A�Cԣl�2,�G�,� ��p{;��ҡS� tv +�݈e��e9����@x�[+��r����#JE|i�X������?n֡H�$�`�iZ�~�f�4����W�|/�mA8s�'/H�;'�vw8N2n�f�w6H&�����k]B���e֫�nҲ=˶9:4;� ��MX�]�ǒ"Wt�+]U�Z{�}�����k,�6�Ue�-�{��n��G� z�o�t-��t^]d�}w��Eo�`tl�r\�me�꺁��jc^9�( �Tj��ѕ�T>��
�RC�o���t��%r�E�4"K�����0�Njz{���j��^�d��U��D�"H7�VQ���v��S�Qm(A�WSf�]��1�a��T�X��@wbx DB����^Y�[���z���CH ��?%��ف:�ڎC�����"6:LH�"�Q�ekC���1���gϽL#j�:�q���R����\v�t�u���7<l��]�؈�@��,c�OAB�ņ�sB~TW�M�Gi�K͹�Xj<��E�e^+x��u֔r4��[0R5(��Q[��/�Y����[[A���;�:?�(�]>��lr�r���;%��{���l�_�����O���Q�I;\�H��9��>�^xu���boA�\�C���fkDx��`�O���lp0g����?^�qCH��yDȿ�<7�Y�%����~��Ow��������Q����t�ZhdSs��Z}�/
i��r�#~�P�GY��C�j������L;�KN=p�������F�Q�5�N���K��Ǻ�x4���$��?�4qb�/vʣ'1Sj��?5�׏�1�!�_�3BX��z��g�&kfG�Y:� ^��Kq	��J��ʤɘׅ�����ːB�X/
�i�Ǯ�/�{PW'�#+���N�?F��[FW��l9�v�.�4@a�#`l3G0�M��#�I�b��.c��_{�}c�������T�{�`\�JX��TRN�T�����N"3���Z���;�Ud6��o����Yȟ��;G�����h�)X��n�B2O�%��5���v8W�c�%�����FƢ�ݚ�X�p��
��J[.�q���ZK�a	�cB/aCHhin�h��ɡ�������[���k���':"x$i��d�n��h��5:�f�gKqۄ$�\�(��p�UD�����fÁ�N5b�$[��Tn�I�s�s����.8����9�-����]���@P�_ry��^_�5�:����3�P1~A����������B(�|����(A��57�)D�i��jQ�#t�����y�'��'Ҡ]t�n۹<�+QR����]������-I���͵�{�dX��ר��2^��j�W�73,Q��vh�n�\ݬY���]�/���dԨ��fw�,��8���	>�pN-�k�z݃8�;��&�q����fV��\ژ�PQ�˧YSw����ܠ�B}�)LuM(̠�4�}iK���k4;�%A�,ۉm�64�-��{���ð,���}�R���խU��y`��29C?�/�7k��jޫ����w�ד(`�ďm�'���s͟w���J�y��t��ȸB�ސ���SU��,�c����\;8	���y%.��?[�
��_k�e��aR������R��DD�:�Co"��D'�G�A8��X�t�́;�d��ԃ�>g&ཿ�ŉ�- t�%wɴA"8�f��
�yV��oi�����j�SfF%;{d�5�0.� O/�~CXb�נ���`�ԍE辎������NM��a�����B�H���鿄wt�<8%��1�|���Ǯ�nj�H�t�Ww#�ٚ~�(;ސ�T��/�3�ܥ���y�9XƋ���m�r�T'	@��<i��v�`O?�%Cg�c�k�D0��X$��_�ny��e�r���d���`�Ɗ�/��/�m|L�m�95 �
��`>��kށ�H"_qQ�f�`2`C����[��S�MvC�����o��M�g��5}�5ZN
���}�m��0 �Ie{S��3{o�g�S�y�1��v�a��aJ��+&ݥc�~�Bp�5I�G��>��� b��|��'f�PIAD�Р�a�2;���t@̰�p��/�Ǡ�^�lY)
��m��Yf("��\���Qi[j�8��yD�E�M9$�s'�j�珕*I�{��Q�/g�����+���Oc#��:�ԙ�K^�/�mUQn2�Z�-;�>��ZSI�ܐ=��=-�ɦ�m����W	�hBH���ޒ�  �#�B$Ѹ�~��Oi?1�����߶�H(�~P�<]�E-=)��út1�R�ڥ�KPB�=�]N��8��٫�S7�6\�OB�L�)z�q��F�%E�- �݂e|��݂��5�`�&ߜ���z��V�+\sQJ���R�i�=uӤY(
h�����1;��!�Y��}"��^�27�L�b����W5J(����lǝ��L�:�}��Rm������q�4�i86�yNeh�$�����5��Ⱦ^�W�OW@����Ck^k�L5�c<��wN��R���ʒA�h*�8��
@��L�uT�9�ɷ�8^�Ӎ��CNꉆ��G�;Q'Q��3�C$$f�`&�X��b��ę�d~�%E�jS�e�y�ֺ�H�:gF6���^qH,��ۻ�x%�����A�"���om���P�C�Z:�W���e^ݜ!C��_%�߬��<B��*��G�7R�+�ܚ�	՚s�L|�.|�̪�i�Vʨ�������x�t{
�����cK>@;K������s���݆�Ԃє,�*ªN]q?��3Ƥ����^�ڛ�1�E�ݰ�������,��$��
�A �Mpm������>�<Ʃ���?~�/��1��O��/_�����R��7�o������Q\��J��mߖ _Q�K�����n"%<��tY\� B�K��!�� ��04��s��r"���ov���)DS�������W�C��f=lt\�'����h�%^Ɗ�B�,�_����t^qj�cJ�yi�^7��
��<o��r�uYG�&��mx_�z���dׄ���0�5ZE��+H,;�B�hK� X#�)�8��J7 �ݺ���>k��gUx2P�V�Lᛘ
�
���ם� [���4���w7�����"XD:�4�j�}S�d�n�=����4�X�h.�M�&�J��7�f҉S6l�[/�5Bksh��Y�c1Xl���Aq&����f+!�<,\�nU4o����e�I_�f0���y\�h�U�6z��Վ������C�8��n%�}�	=���-#�K�dG;����7�V�<�Z���<�q�	���E��:�i%Vz�`2rA��H�����+� �;	����:K�;~��r]����$��M9V�Z����W����;3|ZL�#bbz��Z�:�&��N�S$�^���'n�u��!�[�����F���yQC�$��^0Io�X�$��	�"��׎/>�����GL���NO�v��j؜Lى�Ȑ��r�����:=4���iI��J�їg(D�����އ�IV҅��#�)6�Ѹ��m����P���jR�	�C��������<�U7+�y�w���Gz9Q[.�
2��f�?�M��3�ϑ��3ظ����W57ղ��ÕD�BM�����1a[Y5�%g�ﱾ7@*����S=���?��9b[���d�!��\��z]����.n���0���%�pm(��/'ӎJ�AY�I��ڶ���تM(\��-V�r��h�9E/��T�PR�ٍD����q������H���"	&�˨���̉/M��T���B��,Y�dξ��p-|���Z�Ve��{��n�2��Jr�C�/����׶��G즇�oY����S�
��CE��h�����!���}�r�_"��*���mԭP�G�Tq1����?���9����;�m#u�W���2�%-�צ�Uo���C��f�=m8k+~�Uf��O�sڎM��\�3���{n�,���a˸ި�B�b4�ȵ��t@�	�����˯ۙ��\�#ǋXS�]!H���m�����LA�.��� �39lmA>�7W6��w=�?���x������tFD�4�G|�ܔ-�4jy�(D3Z�0���՞pɿٛ�4�1�?j�f@����C�Z�d�=�[XB�k���l�Db.�1�ݬ/ە|)<��^ec|dÇ�]c�-���Y�%�}��t �M�S/�1Ê�ܼ�R��L�&��{�+R#(ծ��={{�ɳ6&��Xw�I��'��"-�,j����-������B����� νu��Ȥ�ݐ��-Bțh
��g�ĐD+�ɱl���dm�-)�$������!3���b6XaCV9��!�&y�i��h%P{�e"��qF���9�޼p ��.�d\��e_�B��ڡ���������<��J$ҨpVe���v��QE*�.����pR�z;�&%��&u��~I��U�ƓQ!d�����đQ�׫����F��Bq~�[��'��[�y"��Q�N���d�&n�/"�{m���T8� ���7�����s��P�i#��9	N\yOV	�.���9�^�`慗:���Ǩ���,��R4t�<M
��;�ò��+��M}Ђ��/�	p��#���q��+4н��c7~�VLI��a�2�liS-Jm hk��*1��,@�
\�2f��H�t����`t�� ���U��XT��֤�1�R��f n#N��� �=SD���؝��`ѻ�n�����MLs�ZU-�b�p'�g��Ȅh�:��	ho:�Ƽ*��4M�ԁ�(��O�%�Q����X�����؎�Mcsp)�]�]I�N����:]�L�Y:�@��L�J�Q��ꗴ�A�w'�����{"�� \i�6��U���'W��vPhH���\�����y�w�p^p#�-�uB��.7:��}��~�#�;F<��b_��~�Pu�ᗒ�o��ܖӯ$<c`�9&�|�TV2� +S���Ճ��<�[M� �[�A˳�$�Lyt���}��l�����?W�S���z�q���|Y�Y���Yf��26��NgK捊Hp,u��e�L�^� �
�dQk��xZ6gRQ�66��5s!Q
j�@yn1��ŮH������"Χ.V��'�"�95��3��&Ъ=G��8l�!Yߔ{���9��3L�ژ�w�Q��%��7�]mt�֌"�����Z��FuPb���5g�d\$�u<��}?�$��iF�s�^��ɜz�O3�cy�����
̔�6v�?�lI�8��㷌��d#��#� W���DO H������B}��R�Jj.���Q(����j�r�A��v�.��I.����R��_1ݥ+65i�a� ��<�m��Q&���J`+e'�L�>�d���;�.|�~�&�G"iq|Ⱥ:%�>�+U0T��V'>ω�����f2ui�B��u7s�e��k�Bw2QP�羴3\�)�F�E�_7��[Ҋ�����S�ο� ���X�B9�$�֝� ��,���Zn�{�hG�Z�p�h�hX?�c9AE�(�����Uaf*�Ȋ�3�<�E����e�X��{$����!��^�1#e�����l�f6 LCt��M/I�w֌�?�U�r����LC���%��I�����+	f����G�ڔ��j7��xK-~�����7?hV#���0�����\J٦����.�O$m�`�V����ʫә���͆��[e���er� �W�&�1A��ǣ�&9n���)oV�i�.�&a4n�y-�d�6{
6s��GV-��lh��gT�o����z�=R����[���haӫ�2*F�7K���sHߊY#W��U�*�c���P&�H�]�"0�4���<�DI,�;?�n���JA#?�Av��\0[�d=����Z[?���:U����y%��x���g8M��B�qd�0(@$����g:*Xn����`��tJ�R�Z�����^���ߎ�_�"��s�]/N��=8X���<鎅����r�v\4�FM/�$���-�-w�Yhl��QeO�� `i�`���t��GC��@)R
������[jUAZlŦ>!��@�i*���|%�B��'�D;>��D*;b3	h��6��dՂ_��Vэ[��Ļȕ�����%z\"��߻��H���E]��)���6��P�wc�{�3a��~�E��)F�t	�A �8��9/v�c�v �>�k6ms��ċ	.�q�?S6ש�e8��]��
v��z��%y/�_zI]V�].�pL��y��'�~��g��md����A�� "���!)�9W���mβ��wGq�!��W<�Fjh��3�I��)y%�O��i��ȧ%` q����JTU��o����q�)�Sӓ�Te��W�fhW�
Ⱦ�rA�Ʌ����P���@�.��U�w����ThKz:`��2����Bl��Qɧ�]�Cť��:1�L�	��L�n�춀���r��LH�y�R<ς�t�ꐍ`w�O��in�x�7k,8�'4N*!d����6�bYW��	��"����v.ƅ{�n��hh��>aC��&ˢ��.rت�2��݄���<�f�𑓆�Bg2]����@���C�\̫�Ov�'�ku0]��1��g��ȋk��5H�i�N�q�r��2-�?EX(�f}>���r�1v:� �=�Z��|-֊�|߯vz�h�I/�=[2rAdP���K��՜Eu�揝$gz;��� �}�w{Z�.��C������FJ���m�a�AJ�dPm-h��+b����ab�ך�����+�5��;Sx��p��wo�M��ڟL^�8�2� K�����Y��G~�԰�e�	��i�I?���k�	�3���'lV�5��&3�+o$c����vK<���t`�C64>� ��@�t�$z�ړ�kɺke,Uo����n��B<d�Z ������*�0��g�v	7���"X͂��5�}����
�_���S^l7������ѯ����7Q�0*M��L)�[���3��෨Gi"V�^����&,C��;3�=9v�n�:`��}٤� ,����âZo�y�)� q�Q�A�
H��D;�e��Mx�5#g��K��������sg	�䚑u��:~��)��z*�ﾀzf�z��%��hDt�'(�R�&�S�ՙ��~�����<R�y�}pY�R�؝i�:��%��ϫ�1�������p�4�8�R��6g���nD�E�%l�����Ց�3��xؠ��_~�ex*����<����BejN٨P4Mxߩ��}�Y���PP����ʊI�/HE�Ґo�{�6m1��$������h}L���}�|�iO��q���d��;�l�����i��M��E�t<�כĳ=>�9IC��BԾ_Řu�X�P�:^�S��)+���v�wc7�F��á�i��	����'��|��f�(&6��r*^}�M�j�'l!�W�ݞ�b�rF���Օ�.Br/��rje���U_���;����6[Fw�?���irj�|���Sy�YڧŲ�5	�c��������+���ȟy}��D˖�)N �~>|K��
&������EQ�m�?b�D�Q&'�ȴ�3���"y"�C����w���g�s(	m�����#�>Ɯ���n�&p<�P'1D9�ݿ�j�Tޝ]�Y�1+H�'@K��E(���6�D�tA��q����@��N������2�%�j64@筛(ܒ�T�Ӆ�}J
2e�����4��ҺēX?�g;Q���l��z�̽�A������[�2��64���k� �)=+�U4-�E�A\\�����-��* ���B#�)�ֽ�ldλ�Y`@F�W~=I�Q|���Ѕ�S����M����f2rY�(�llZ�vg����Q�
��cMTs	p�����N����CB0�����Rk�G:ʛ�(�r�9)<cXr�&�'^��"��;x�[X/��Rn�b�BJ�rZ���6���x�YY�Qk9���U�1�5�c�vT4ڈ��cx'6ͤ8�O����+�ASs���1A�|�q�S΄T��Gg�t]�N�����<O�L���R���p�����Dҟ��T�y,�,�d�W&�����_��-���\�2wC�0]�j�cF���i��P���+|��H#g�aYY݃��CO�^c���y�h
&h�3\t�0��鉌���lL�����SHl�LM#G�'13�1b��e�o�=���_�*�$��D��� ���1��8���5��t�~���lu�����~ǥ��2K��m��3r�!�z�s��F�,�j��3���E�s0D*�����e-�A��"�G���u��Uj��=��KH&�����Y�)`!�=��o� ���O,�lM =�!�,o�+�\�yq�A�緃�XlO1z���g���PP�չ�.� �'i�om��w�(���m+dςx�G�0Ak�L/��cs|!�����f쾕��l�����?�}g��P�5n�X#U+�*�\�ʡ�g�p+�֩=�ll
�?8A|"|g�Τsl�7�/a��j�ȼYM�D�OF��c�]/�a��~��B?:�tWr��6� -�����4t�y��	�姓���\�K�$b�Eq=,�"�^䛦F{�}��ܟ�(�|xU�<�X�9c�q*�N��_n�{u��d�<�VBG�*��C�*`9��Jh�ܠ�� ���k��C�!L�:�9C�z�{�ᨐ[���\:p���#��s_�H�ݫ�7�'H9��^跠(NG��b�Z�5ti��=��$�r5a%��O�T��d7;�������Bsɞ�B���S �bT|�Kq������f��ꨚQv-��5<�8�I���k�kѷ�v�T��i��V�c�:9����]���Ay����SR^�@5G�ԥqs�<ūE�eʻ�宙���[�rnI� ��{+��x?%Ð?����ʕ+8ЯZ�+p����3���*9�����ng�;�p9(:�&�;Y4B�2~�'>�9��Q����Q����6>���|߶og&��f4j�S�r������1G���`�i������E�'��3��P�_��!���=
<��토��������3��h�����
e�N����<��S��jԽ/�y�:e�Y����¥��LưK�3D��0_T�� ���v��9�_719�s@e��������_�$K���T�.d�c�_,'�3�!�Q�c�Dj�sIj.����!B��#���ntqUJ��=ނ��-�7}�t~�#�g�|�,�&6oT�l�Tg��T�1�͌�[^�3���k��Ӿ�Qٺ���F����^&ı�3fM��N����|c(��[�R��=)���	��Y�1h-]@:��?��a�����Tj�y���g�n�A'U�` ��e1��@H!8D������S@n*�	d�������'��-�g��W����.����b�$FxU�����`���%�1���3�6?����u.��v��h�Hjb�V��YU ������B��<�*����]�a��\�S�BؐP�'L_���]"�6�BƢ�Nv^�X���	�r->�[w�����Eل�27C����[��#~힤L�ds(&TV>vv� 8�������U�NK!�Kb�]��o��<�:�0��1�G~�s�]
���_�+�O�+�jt[���
Α>S�hj�iM�k�w��0*�]Ey�1H�:ӏ6��ID�3Lx� �`��2nH�0�K^��}�ã�(itf��Ƣ@�5�ߺOٹ���W9bȍEd^�{JP��</}<����>��!� ����;"vim񑸜�|Hh��ڈ��<�b��ǜm�៎v˺����m7��{0�j�Xv�m��nG3!�������S�K��Y06�n��r;o�m�
��h~�h�,[��GX�%��@�r@lY�E_K$��)��)S|�����Ce:~/T���4�qR��{OH�'r���eY4b��6W�`�x�e��T*�����ʿ���Yֵ�Ia7�Lé�3�H�4q~�<��V��g�qI��B�m'w��X�:��1��J��H�~�Mxq)dzLB2Q�xk�@�E	�ď(5�2g=3x	�I��:.��g�:7�:��Ф${�Jn�@��Lu���=-���Θ̵=�'y��B���4��dp��IG%�L����/�e�
`wy��P��uS(L�ྰQ�V%�����' ;�X�o�������f
��c�[�Q����۫�nQ +�B'���+���o�I{}" ��S>6f[�fv��,�U��Y���FW�o�/�u#q�O/����E�d������Vmq�[��@J /@n0M-��/����>��CǸ�0�ѓ'֕x�O��f+��۝<�`�� bi�e��j�彑=��9�:I���d�'�z`{6�~�o��~<#��R�-N�G�R9�����6-���n�e�R��lw;ʎ�"tiX7�4�։G�|��d��A�7"y�j57j95�y:�}{M���0R$��3��{�9$��S癴f
=�ÿlb��ga ���T6f��\țzZ�mazV����Ձ%o�+m��[O�����I��z�p�IP =���=���|*oh;-�ț�#�	{��,�K�Nw��I�,/Z�htߤ�9�^� ]�%rZ�B�����T�0�3���[�ݠ?�~hK�572
�v+;����-R[���6�?%��E��9 �>�N�r��B/؂^k�⑲��lsA��A�x�/|�&���m��MU�-_�~��i��_�/q$���	}�k����`��Nsoy]��Cq74Vݏh7 �Z���u� G0��%J?��k�c��~R$����Gqu�Zm�/E�\��8����Y�j_Uz� t��>���m�S��SRI:t���r���W�d$`�f %��!3�J9mV���	#X�ee�2N E�)����-���lA0�0ۺ�p��@�g����7���4hh$e�7/I�]��c��k+��Kp��p�R�j�7�Y��QB� gxu)���TT�J$�@���{f�5ʘ�_R�\�Q��5�uc�RpOqqU���6�����y�P����;0!el�����t�_�q �o����xe���GrRWj�����xh/��f"�`��,��%G��E4�כ��|%݉�+�M�=�m"�7X4t��D�C�� ̈́���B�R��C��h'�BgR!j��rb�#=C~����[L~\0��?�Vs[G�??�|Fլ��O��O�TCۚ�� �/�:QsSVT߁i��qϸ��V�ADj��<�����P񣥇��wM�(#�zp�/{�v]dF=�Ղ��P:��6�(�<�}���h�yM��e֝�}�o������R�8t#Ӽ�㏺q<���y����ի�6R��E��ǰ�u����j[�0�d���X�[��2>�+n��*�|���)�9ϟj�{�DڈF����d���;��E�Wx�8[$��
�N��"v�Rͅ�=;��`���a�CJxo�dՏ���>h�+�:h��LоR<��I��`�* B�&��ǿ�'>q�݀�t^/�]��h���u�+4�eݑȱV�"�ꊐ���v����L D�H�(~�0/�L)�p��=����nt�;�i��������ڂAY�v��ۉh�&���Xf>� �_"��d�f�X������~���:ԑ��'�4������`���
�~����U���m�|Bo�_]�M7��	G�Ε��þ���>��,�g�4�lV)��|����&���7j�H�qD��c��?�VƏ�+��j��=�G��D�_�� 4Կ��$ė1�>%c��t�����(1 y~��Ͽ撧D+a:>+�}���b3ߵěg+��9�c�0�C������)h_��1�j��`���fK������:�ǚ�Y~�ή�\�g��n�|�G�~l�dѹ��������s�Nс^�F�E�@�#�����KT=�V{�[���SVޫ��)���dn���L�hbN�<��
a���9cH+�Q��ɧB��������B�=�Ng�53����4;�U�����"���_���h��;��)��*��IL<{�D���shB�!����f�n� ���mL�=�<�%�Ɛ*KUK�t�O,H,n1���Q�n�Y�m�A���"�#�e7��K�T��}lumx��ь��Koe-����L2��H�ATR௔�o�Z�`)�A�����b�k�a����L�p˥7=��dɟM"�(�}�W���O䨪�/�r�4�``i��/����f�3���Q����
��r�r���� �e8���U휜~:^��0����-���d��V� ��ߍX2�ܗ��1/�M��:T�T.G�%R�3��F��'��Q�!m%D/��E�dX8�d4����Um����&�ș���?�s �?E Ճr�F버1��=H�[3Йs�rA�~�1s���0E���lO>#��f�z�Ir�֌J��J^����F"%�� �^��C�u�8����̥@��,���x��7�Y8�c��5��!C�1;��+य़���h�^'�4L��;�>\w�N|��S�C[t`�
��B��RJ�񑗓�(5rދ�34���=� ��޴��j�� 2tɶ9�ݠE�nN�Q�X����>f�dM\�o��R=V�f����b�4�����A�C<��*�^hثۓw���D�3��^����ď6{O
��8��p��ߋ�N�^H�5�$���A�9��ѿf����vG�ȱ���N��J�+d�J�9g�$gV�
 ��*b|�H�[�}9��R/��+A<x�5�����v\̽���o�M�b�)tc΀�^��`J�g��[k���rJ�% t�E��2�.Q�⌜b#J�DiCi�����R��0v���z:�VsRz��7:_NE�lT�"�>�~8�X�7����˖�rh1rAL}����ۇE���R��e1�pz�9�T���"B�B��j!Y��ړ^�M��]7��B�E���y���c�Υ3��8�˚��)�	�E���*Z$���\]�S�6��b�>5ͣ���su���c�]�˕��A}��Q��:!�V���Iڊ���g�ʯ���r���]í�L޶9s�s�ʙ��ݘvA���ܥ��!AT�N���y�ۤ�F�7�7z����@�6�4�w_��܋gg���������3L�3 �<���i���3��c�1��v��.#�i X���6N��:>�t���_��Ȓ8���B��xX[����OL䕸5~k�N�+6�K��c�х8x��[~���h����R�M�=����Kf�Rq��W���T���;��M�4rO�|��z}���ؖ%LI�.�{u<�E�yہ�*W�NUxH��6}%��i^n/wh���K��g~�< ��]�eFM��c�3�85?*��)��$�v@�"��٬ �u�aj�y+s�޲rY�I0x�'~��.'Sඁ�ce��u�1��X�G�q��Q�����R����(�.�W��w`��9�!Ʒ�Ѕ�EwR����Ǟ���&Ge�cT����~���%v��0����B�o/�p۲X0~���0X�ߊ ��>��qHQ�}�`aF�u �ݙb;�s@+5~���M�-A�݁bT���O�������Mo(t���&�	?�x}-��8P ZZ.@H�=�J�����k���J��2����J�O}0u>��g�;�H�G]YƜA���{�HP�X(��fn�Ѿ�Œ7\*�Sty����4>0}(�F|�(�Qn�fT.Co I+�@�7wB�ᐙ#�^�����e�."~M|���U���T������T�y��C����1X�^� �v��j@D�e��0[����,I����O�%n`E��2x09/=�z�M���3݆-*N�̏j�v[H�Ѡ�=w����ͥ���/pfm<t�8	&�3��H'�<����K�5L�Ô�Z��i��NG�&�ƨ8g���f��w)^��v��#h���>-[�ܕ�q?����&5p��7�@]�WL���|����W(D�����3¸�������Y]K:Y+�xa�8D�����F�d�Q���Ug�vӞ 0���b�"�L�v��1�Q�|��VvN��=J��<3-q"wJ�"����~�bݶ���4Ђʚ��="�`i����fTWE�F�@i^O����l}A���T&������j*v�~��"y�G�w���]��,٭Xj�x�ZΣEeL#�ε�ن�8��*n�-	-����,�'�t0Ͽ����2CA�X�~4bH"����8�*��76Z	�VkhB��J'
�k�0X����흿�<�s�^�����i=yloҍV�ז�������aI��u~z����B�+s|����IS�"X��r�/a�ׂ03��zB&�<N�qd'���Z�>��ʭO�]r�]�DφIh_X�|�-;�#^wAL{�Y٣e�ca-�{��Pp:�h��ְ=�x��z^��,�z�q�8�<��1��z1|d��+~"�5ki1��ؔ�;(@%/nNe*�wg���Gɚ�><�(
s�h!�8w}�Q�G�&|���QK>����������Rw�'}���V���Popv�]Mǆ~�۫E�@��tgQ\���p���7a�/�j�O_���g [5;C���M��,^�I�c���lN8����*����۠۷J�;�"�U�7a�j<`m/o�'Ur���7B�)���q(��!�Z�1����ݔ���Cqhr,��L~cmr���;�CA���\?XIh����\o4��B���pJ��^���Y��Od���
��.����j5*go�k���Mm�[����ǔP�D�FY��}�3�ME��N�m�o�,�@�Yn1X��N��l�¶�-��>$����"�E�������Mx��c�G����Z٢������P����Bg}B�Id~���<ķ������Z���^8?K��P/��$j���ã;Y�t��o<�sB��u�����1�<�.KK���'�O�}��9��Q(����Gc� EF���H�1P$��9#� �Iʄ�R�w7\;��9����l���m��������(�Gf����9�,�����UiB"��y��hJ�x�z�DE+;�;�G`q�st{|T�~ d��1��(���n�$��|�&��>;
��v�E�������ر3E^�I���Z����_K���`8b���Zlc���2r>��bgb��8�٫=�)�'="�����1޽{u�&/�GǛ+��ߛB�Q��٥�!Hqއ��7g<���ce�;�������.A˭�{$;��f�*7������[�*�n�����\'saW���턌�����h6�ʓ�����b	R�0Z&�:kW�����v�b��(��قl�I<UW^�n!�� ��e�e�_��h��J�R����㚞���@�K����*��Z�☫���l��a���
��yE1H-�VD�,�x��|;5S�&uڃ�����q$a���q�Cǅ$����|`A�<�<�*E]˴F�����f�ݚ�|�=ʝ���̷�֙�����gXi���dFI�<��ϣ�Ƿ��>J��f:wfg�F���R�,o>�u̿]o,���}��#�غ�8��gP�%)�����#2��BB����Go�[m{gΩ��]>B��_�M��LU�5�y����0 i���zad��3U�*l�m�?���j��a�Θ,�}>�?��4]T���@`��SjF��`l�O@E�L�5�X�9�J�M<�1}$�Ar����9�2PBuM�W��������6���ԡŅ�d�v{۽����ԏ�J��HK^�l<(5%"8�>�)��ј@q���V�?c��/L݃�~BܺY͋˶et��JU�7o�Ӽ��k��Irlok�]=д��7+tYZ)��=��b*�f��Y��#��n����ܠg/|n1Y`�/��]v"�����r�Զ��h�x9��al���)�,QJ�}���Wv�#�,�g:�"��R�����;��υ(���]�e8��R9��m��)1�1d��yMs�Т��.l����V[�}ϖ����za���]���L�sƘ��g��v�X����֤�f>�ِ���B`��$�1�A�g��W�r�:��r���2���.��ȵ�ꑸn $������0Ҕ������9�uY;Fl/�(�G)H�x&����e��B�~U�)��;˯�����Ic�hײ�5@��H��{��5���	�|[����l;W@/�s$����\71B�Y�1Q�ǒp��7�7s8QO,HB�}I�.�T��fK�.���J�'�%[�=Ԧ7N�v�������wgwS�"�>m&�������<yCZ@p�I� \[���z1�����{˙n+��� ϶�h-�I�������9bf�^(��HW�@Ĩ����g���>�*Ou��5	���%�b|�ˏW�u�d���S�;��M@ea9ލ���MŒ�Pl�|���k�K�+�7I���G$��	��7!;h��So�ϙ�ӆ���.,K��H��/�~Y�R9�ac~��������H|4,j�^I�EI�`�I�"�i��-!U�f��mۍ��ֵ�Fz����W�b����I�Ϡbz���"����Ɣ0*q��ܯ�y����ˌO�s���e,�"-��IU3�XN�{L;4��[�2���2�t�0�������;&}�MX��!���ʠXF���99z���8���0"׿��̈�ٶ��'�
��I��z�L�Lt�"�E�����9�?���t�uQ[Qm3s��`�g�����ݔ�z��:�Q��zBO�Y��),)��R5�=����Ҿ�Mu��h`��C��L7��j�K6�*Z#� �pi07��1kk���C��?cF��*�y�@��G=堂i;_!c%?D�}ђ�������(w	K�v�%`��<W���mOgta8.��j�~�zfG�7�J�>�
gPK<,\L�ѐ=�wQ˒�!!��^�Q&��C��;�zAR�[��l�9u�S�Ÿ�K-�t�|�踠� �w��9DH�k��4�t�.I�ұ�f`Z��kvgq 1n����w���7b!L%���7uU����U�����ݤ�]= <�p�V�ۗ2;��u��䒬���^1ʅ�� `�
�c���e�s�S�|ʰ�U�[h��y��q���7�g �����ީ~�.��]�9�r�	�o��tlL6�5�,��V
��|�e�A�#�<���Q�%='�k�����v99��7;��(2
�#��� 䞙�ƳS�U>\BI[��ģ���ѻ���&�ic20��zq��<Ŝ��I�����j�Ȅ�6���$'$,�a2^�mpy���ÕX���2E�r	���#E��ʲ�=���ߣdy8U�X����[N�kt��=�j�g���a�Rk)���d��W��.��$�vu�[a&���������z�/q�*�
�L��c�`
�&�b>^�4F��W2�YuҸ��ȎTТ��k>aQHf����Z!:�u�B0v���w7c�����y�iƯ�(�����yunT?��q��ڬ�$6�Qp碡�����2�m���ܛ=vxe��s��]�5������J)��~��YE�qI��f.���Pz0���߇C�_���mт�t%J�H?�_�{��)V�@B [�s=�8���8�8}���3e�;��s�l��j`w�|w���y�}U���獡��86f���Փؑ��������K�t 9Z�N�N�{Z`#,t�`D��LE���#D��6���[v܂XO ��(H`.y�X��sq�v�I������][�YH�y�*kxj=�Y�x�Q������E�O^�;/�g�w���ľq{��#`�<�2A��^��[��
�^�} �E#�S���O���wQ#3w��`s�O�T��E�|�0ѫ�em�Y:{n�x ���61jE���J"f>\��Dm^@�a%/d�2[v�W��l�ռp�����$���jT����o�w�.gQ��%t��eߦ�v�Ϙ����K�i'VEj����_ޢ� ��=�Y͠�J7`���#�4U}u�����!!(��-qdu�'�ݪX����Y�N����sZ�b��/��`�q����� l���G�p��(�����w�V�c�_\v!�qq:	(q��X�Ov�y���l~��v�� ֺ�D���~��0+(*.�l�PD�07����.ce�	�j<��$^�y��S�>˝�Ǯn&��K�5�n�KX��!W5��Y���G��T���1|X���1v�T	:�l�$��a)��'r�2lˎӵ�f���E:0UVYX�"vn�[�ϔ[�����q\��ȼ8)��i��Q}%���8�kvB�A	U>/�o  �J��B���ʻ���w
�T�r�8��N]����a<���t��|9[���.���G�F+��R1��@�FU��F�_w���o#%��}���r��	�7��aYS���IY �Sx�r�ma�%��p��>� *��F "34����E����~��T@P���o�F ��ҩǼc:t?�~��v�N�i���jJ�m���,�ҋ�D��7�H�-�4vqY�aݣ�&J��������=&�]��A�<*7$79`�/��klN���Mg�/q�M���b���$�M�^^ P'Gp���1k_�����5���� w�swJ �
�E�{M?��&�e���uv?�d���/�K���$%U/������};����W?����QP�2Y:���t=�f�~���Ь/{��7܋�}�|0�{S��Rx��Z4�9-�HΚ�}oz�k65�B'Bњ]5Q,|��o�p¦e���4�ྰ�g���O�z(� 15 H1߶J������W���7ߒ8(\E�.7.�}wҞXG�K�ں�g�]�*n��v��/����@�|w5]�y4Ĕrh��ƽ�r��d���H���=t~��Wv�ˈa�K)N�5qՉ��A˜r�����z�	�f|�͐�fC���!��<zM�?m(�O�o��T�<_��&͇��=�G����bm +�j��$A*٬������aYr1�<�(8Z�$4�E�L�Dv�`م�{K	=�{���Ci����b4����|r��q���jh�'~U8@Sެ����ߋS5}��.�2���E��*9siu͆$�#q��(o�rF����wv�<�0��{{Ih�#K���%�}�:�+[��)G�4�G,+���W�kw)ƴt�-�]�
@+o5�-�#N�l���!Cj70"��,O?��?|������؋����,su����1jCY"�����{�6ѯ���.N"�uH0i���,sV���*��a3�[6b@M4m�H�D.��Ba.��S��L�9�[�iāY�u_����l���HD�&�,ըR�dv8ky���G���:o�\�U����43-ZL���"-j��G)R4&��� N:��"�[]� #����iD�9 ���*J���R?Օ$[�D*C)t\ǰ��<��UF�)��H�M�]��|�v�i�-%7��=wY�r��1�J�s@Lv?���q�G�~ۼ�y$Z�:���[>�L�
�|~�.@=��Qt���� �J_8�S�HZ��̅Q���L����+~��P�l��f��K��^t���/���G�W[�Nغ�%	d���8-`�ٌ�J�.��b�o$����S�)�S��L�E2b�F���|�Ě�_��<���a��2p�K�ݝ9���'�%��?T�!~~-��HX���aK���Е��gX�0�%�5���-0��+�jMo���s#kɒ~����1<ڶ>�����#�U��Q5f�m>,�Q��َ����I�4�j5
���^��߽X��e�X�!x`��"�P���Ub�����0n�'!�>D׳��7�.� [�38�Y�_�b��Zm�$���b�[K�7�Ĕ�ԕa�S�R�3z�d�HUxRL��7�n��k	 �6���f�{���yV��y��kʐ@[�Xc��:����uۏy_J0�OqcJ�P���f�4EI�WV�9I��<�;ȩ�ƥ�!AMfjh�9��9���\#��4��Ν����̳$���A f�"���b�}�Kkqѩ�+a&�\�N�&����3w���<�T�x����q<���&��'��3��Mӿ�3P�g�IG�$�U�����4�G)X��k��=�4-�� K��C�0L(m��{��d�uU���b�eA'�P�L�~V�qV��A� �F�V�b�aQql�/��p��(<|�; m�.u�'PoW�b{�u��[Xv7$B���9r��a���(r�Ǔ�=3��3'npepǨ>���;s����h���	v?^�E��z;��"��B�+ڗ���4IU:��Ǔ�bA�+v%�9M�h�f�˖�h>�d�rt���=&���H���e������l�c(��`��W�g�V��淪�ײ�	WG{b �V��[4�O�<d�H��R���ͦ�W��/�G�PN\,�����U��s��6� �u�oP�R��1s:'��QaTC̠~���y�ʰ�A�<�����E�ٰܟ�IQ���BN�Zd�D=]�b��G�˂���2a�@�q��}��<�f�!��$�**��7#F���V�nA;�BjW4��:kܵ����av�K�0�,u��b��y�6&��J@ƚ�Um��j���V$�:^�N�IMwgƾ>�#�m9b���s�)C��C��]6�|�2;jwu�����Vi�:J 2s
�)�>k]ϳ�F-a+ǖ��ܣ*��"��1����:�HƜ8*j��*P���m�i��ly�|�Ҳ�vY�� �PZ��Z�*HF	�c,�N��bA�][�%y	#֙d�2.��P���櫊��6�c�{�-���JcN|����!�]�@{�[����@��*Ъ����vi3Y$6��;��`��a�Q�=�{����_��̳��F|3�.���/�$45<	�Ny
H�V0���:�M��qɎ)E��k�I\2I��8O&��g�JqT����E�:�Q�m?�ν5sPO��Ԯ�U���k�VB+�M���\�ԯ�$���+��%+4��U�"2.)Ǟ���˗�G}G7�z<�) ��Ě9�#{��<B�s�kySKԉ�?��m���?�H�� dE�.�O�i\P��{�G��#rd#W:<ȹ��{��mer������@�PQ����4��A�Tv�>�cm*'���[Jν��|�ĂG��N췦�bZr�C�}n4����s��&]Sx���e���Vh����.�)%ʚ�$���v��xr�)��8	w���Z�4HHaΕ!��(�	K�|�>����t}�Ԥ�^Hg���>i4�5�<���Z��;��Jc�g��?+���n-߲S��b'�F�bͯ�1P����L�\�˧?;�W	���K���g~���S�G�^ѱ����,��P�\My�����׬[Wm��gp�bP'�ǡA?�RoB�z�}��_t{���S��s��J��W;�+q���Yc{Zu��*V��Jsȓ��.��]���a�E�~�|��8Š=�߳��m>��a��5�l$%�0Q[#P[b�oг)�\�>,߄`�ڗl�b�SA�{r�$LQ�q+I.������t���rP�z>t_�jB���%ٍܦ^�]�87?,P��zy������`v��z����b����S�2�}LIWLc� D���p^~&�!56,h���O2��t�F��u��Ơ2TV5���(��Ժv�f�����D%���	�s )y/X3>6��Y�m��>Cv�0��#�Db Tݥ��Г`����b�ѠN=y����ʁ7f#��l)�\�!��ܗ\x)Fi��PD��#�i�3o�����w���I��A�c)���`R����"����+>s ��g{ձ
7����?��gN�-!�<�U���q��@��C���F�q`p�'��o���ɋ��a�Q/x�!����A��м�߯���v�JF�B���n��(���� ��II2�3�<�5fU&}�y����h��÷?�mO�2�o��v�P���e�����e�9-].M�ZԽ��oϜQB{Mu�lT�V6L^Q�8���R����ԁ�S��h�Ṇ���ب����J�l�&�t��Sg�5�]�2y]������	���L+�ƒd�q�%�n�ov��|v�i)X2�{���jq��N�����
���U�z>�u�%]���6H�p�!!v%�Ɵ	���0��#E���O��x@��|Ѓ���-q\�o7��� ;!o8.��ۨQ+��<:�n���⒴�l{�^���Ͼ�5_�~�g��'���2����ێ	��P�7u��{�n�Y~13%�>��pU�����U��|�VqLL�J���K�/j)�%a�$�d|!��'n����|t��uvT���^���Lv�����9�s�-t�q+,��\,�rX5g�S�&T�/s�.�o��s���T(�ŀf�pKN�����X��]���'|e�Aß��1�1�C**�sR��Ez)E<���T5o{_���}��e~�M�m.e_X�uB ��l��D�R��g�=��m�͊_��"^mC/� �<��ӛ"!,�1�b�T�A��ޟ�2ߠ��x��J
��_�$��O��Gm��J�sʮa*)�1	�!Po��-�Z�+uQ�I��B	�,)t-Ʌ�6Z�F�|bP�`my��Ӡt�-�_GJ�Ņ:�Gyw�٨�.��,o�!�A2A���bg��gGT����X�]�=������ԔY��eٗ�w�Q�v�e����7�qۇ����7\E��c䩳^N�,3�|Z���\����VȤV��L�vx��j� ��I��҈���-Ԗ���2�_�W�7�������@�z%��~tv��&��m.���.��`��2�2�����@:u/�� ����j�$:�j�/����Ҫ.9��-�E"�}�y�s.uճj����N�d�˿��t�`�X��Jm�ж���f"�$K������%�T�V]������PI�N��������V�\��}��=�/��Zs�������sr��0r��^�XF��%Vw�ZI��p׫� 2]�S��)�.��I�\�?�=���\�
�Ո�ڑxͺe�mY���j\č����c�u�]Tչ�=��?�=}D.7� �[�F�����6����Uӂ ��:�]x�א!���i�]����{��OF[)�*�R�"�I$:�!A�FQ �#"�2���ߒW����?$�4��C:j�k�|xh+�Y1-lH�`t�����\���G�cvg�;;�֖MG7��ֺ�S@�=��w��J9��Op�����'Jm(��[j٩YZ�jӭ(�C��� �$"^o�~J`^p'�`4�4E��yr�`���\�Зsj���b�B��v5����%���¨���[�^�5�!�fT�h��+�=l!�%E(�����U_Z����˄����go�����N"]��Ͱ`�"
��L���T�ᳬ�Lh���P3h��^�iX4�]&ß$� ��꫊��T�[T�X݇��zf< ��$� �}�e0�=Y��s%�]l����'J�X4�"�b��p���]��	�R}�� �u����5��L�^�U6��M�h���,�#_oPf)#I=o=��B��d��V��C≜��[u
דx�mъ�OeNL�{�˔+�@�pL�&��l�@��DΌn����5 FF��]���)���qX���8�=;�r���;!�s��^V/��������~�S�I��=-,<:h��d0,���9	�S�?f}���>�n�EiIG��>.���Tt�/<77i�L���H47D5�[�I}:��wQZC��	��Lm���_�}Z�,y�rW�@{ZW�b?0U�b���·�?����u�m���~����kk���޴6ND6U(W��SxbČZ����k��[�5X�>���]kH���d��������}l��aȄ� ��z�֣���P�f�5`'�����B/LE���-��9،0��8�O�@��ZvK�4]R�]�Ig�:*�\㴁Z$�q�=GP6Lu�2��(�o��y���S�[�eJ5�(Hv��^^y��V�&����oڤEׇ�R�b��VVH,�-Ă�/~�K�×@�t��1��
*�ئ�8�RE��K̇b�"���%�3�jD���W��[ e?�%�K��.}sD���M%|#��t�ꑉ�L��_��o��b����8�p���Vt{"�-K��5Ș	�w�pz�òҳd4|�m�{��e�F��{E��]5�}y����jZ�D���𸷬W��x}�Fi�������U+v\O�lF)��S[��qF���D�!l�4(�h5#�����_�D��v2B7V�]t~�8S��f'��^>0J���p������h�J�5|Xn�ƹ���|$'��c�p?�h=��gO���j�� �[�0�"ы1r2ƕ�M�j�wu�C�q���wimy:Tn��7����ܰ�u��/  �^�����v�u��;�O�����k�(��5�ܖ�Q�x�s܃(����4kGs�=�q��PK^�+���d�χ���Ĕ�4(� Ɍh�\t��5?��YP�E�#{�`�>6Sp&[gDJ����U���S��+N���Ӕ��6څʺ'�!}��L`r��m�����g~am�R�r]y����[H�	y l�k2T�B�J!�Q�8�[���s�WA,��[W���jU�J~����j���Ԑ
(��)���$$-�>�����6�?0�@k��x(�za�[�j)��4��&�X�L&�� �c*�涮`���
�NY9E|X��B9�����L~���T��Q :J�8i�6��6q�w]Kl}�Ea>P$FK�q�Ҳ�Z�Gc�:�{����'C����ӗ��q�8!PM�]d�|��#�$f�����������p�y�;y���I����(�³%
eBt�&2m+9m��vޞ�6S����0�-�Y��H_Ԩ`�Br6��!�vu��H
�功��n�hy8a��0�������84x:�W-�� �w�"�i��F�۹LE�5Ħ�מV�x�y�,X�&�u��r�*ҊU�_?�ϧX�
�P�8��C��T����A0n��84��u����X�>�3�?�m�O����R(aFnk-HU�O�~�^(pN���/�x�h�G�*q]س2|d�!�H/�fk��S7�+f��Aޝ��ZW�/��O@1��������n2�z��ӽm🴻8�3��WM�C�/f�O�ڂ:����8���H�4�?!�j���Ӑ��i3u�}%GF��1i��k��Zz��4�����#J`��Q��,��~q��u
�k��s�>t��s�Ǌ�Z�H�r��/}�/5����S�[�X�Tv�A�W���KS/����i){��q�]q8�|��ե��7�mP}�n� �0�œ��
vD�4Ł?���*N��z� k���Ĝ?D��h�Қ~�Uv�5�~Y�Tʓ���8(��.v��W1�2�
�Z*d�к'����Ou_�a��P���m׉�H/C*YO.d��V>r�:����;�b��DV��^�_�}�w�ƻe)`r��q�XUl4�aG�<�gky��ְtl/�mW�y��{B�3k���!Ԣ���Ӿ�1�q����p���}ճ4uM�"�����`l.*m�[� +�'�W96���9u,X���Y��1] �����I��?�)�C0&��e��}�����f��-�����;~��_��l�m��y��]�=���qO��'�eT͞v�]���UAA?z��:�}�z�54ڨ�|R�
6�"I��{֭e���d�&,2h���h5�Z�h�	�|%J�Y�TJ"�R�����J�H��\f@,\Fqe����G��A�c�Dnp���[���pVʄb3���QZ�A�P�n�%Ii���Z���2Esn��^�;q���*Z�QP��S��q���KЇ�}xzj���͚������KsZ�W ��dbGkD���ޘA�R;@�|���vl�G�g}`���|��5��@R��D�S^�A���W�|(�gl�jP�w�*>�s	-u��H�}���{���s��D��Y;���J�ޑ`g
"Jռ��r�#h�E� �8׍�|>}��4�;j,���EGaF�[��eC>S "����w�-����SSs"b<�u�V��.�ee�)F�cq�fq�Bl�MhL+���&�'��3�<'uR�NQ�
��[l'��300�u�� �p�Is�^�K M���BM�����i��L̩{�W��ɣ�pq�9_��$.���\>F��C/'��o�a���Ԗ$��'�P�Y�2F�8g�g��J
|j�-sa&���8�GO��ݐn;$��V��q(�S"�8͹7�@�mf���d��E[5 ee3w}�����|�Y�F��������ԃ�fV�p��~�>�R\ߥiv�1�����o�ƾ�}��QH��y�ˑl��+iQ�C���g�<78�4���^	�-iczؗb�%\�5�9�Xr����rT^Q��v�H9��1�����=��h
v�o(����+$���O����#�U�hMwv�#%�W�}��,y��wI�	��mP�����3��[=،Sb�����q�:q�<Q�w���ff-��OA�Cy��9�|+�؊���$D7o�����_�%h�ץ�K�I���+#^��<�s��/j�������l��ۦ��}ۙ��J��C�3'8Ev֩�B֘@0�$G�86f�>�v�����3(��|���)�E�pmX#�T�=��ˤ҄A�H�S��i��ϩ���X�hi�ê����1��X�ǉ��W�)��� �]��z�}UL�m���O�C
����fJQ^�/M_��2������'%������~�b ��Z���X����`�(m�������"�C1���P��@�D2���������
�[ f�g��1�׍�f�G
�{R�����':�G5l��������S(`��4țJ�;�J���x�JP�e�Hɢ�'unT`6Q��I��O�f$�9�eV�7�8Eh�}�qV��q��C��.��Փ��R�xu\�;Q��NZ�����$نT�_]�y�&�f���Uz����TU�9+��aa���աa7U�Lb7ZBKl,ML]�(K���@��������/��u��K������;&���]��No�������?��{��8r=o�}�R��7k.Dx=+��ڥ ��U�D�B��$������_+хq���]����`M�E��A3~p�O復��t�"�ڮ�<�<��m ���́a�.�xț�����^w��J��Á߱vBn� U�����غY`���4��,*<Y���R��������wh�ܸ�t7��mT�O����K����$]D/qz �6�M�|bT=�T( ��I�T�F:H�M�
�BE�򙆢-^d��6���i535��C��JH��U��S(~���� �mKw��o������t���h��,��g�	�+�G(^��j�����uBߦϝ*W���o��6�ϫ�CZ�F?���@�Ǧ��mF�#fy����v�����,���:�np�	i���W�8A�>8$�:儃�8������#�y��(Mj�[��0��;����Xx]N�<YRO�|��4� �_%����*���<d�bN�^������H�#c������j�¡lѼ��!$�`D6�N#�RYVY�����GX>�Z�K��?a����u�O�w�ˍ��Փ^�8�b��=J�yݍ�S�O��n�y/w2�guK$��Wf
�^ZpI�cy����@�w���m����9�g��&�iJU:��)g4�eK]���D�=�D),l���i0��(nӤ[eQWi����ݷ*�&���Q�c�|���P�j���]�����΀Mwo�S9���ZoSi�l��3�qb����hb	Mqί��:�:�j���h���0_rI�%F��*�k�O+�9�h�/�f&3�*�0��m����Y���)���v����x}���s���A+c-\CbE_��̐��.V�k�E�F�+ih�(}.T�;k2��!�&[�Viإ�2�p�R��%���j����Ւ%>�S�܅�BnmC.���0a&���}�m�7srЩ��gz��V�\Ĩ_�}[4�Z�>nDZ8�ww	to�؍І���ԛ��gUCm���"}��`2��4��Art�g��y@�ꂇu���&k������b-t������Ke���@�c���e�1wa���-.V�i̘o��M%ٵ�����g}ߟ���
��ç�G���үD�x�.D'��/g�l�9Z��{qF�O����<U���8q�[o��u���ȜVC�1���ɚ&���e^E:o�۶����{��H�C�5���\]A��fi���#���
cASm�#��v�Dƛ?"D[�#ȩ�;񧶢��mVɆ�:	��wV�$ƓV ��ȋ_{��>X�[���V&ڷf=J�S�l�?IXqR�暩��b/��eif���	e��r�_х�%�:�,�7xe�\'�"\�x3m/�k�]��P^ +{a�f> �G���U�$��ƥ2g-�1��ނ�"5x��8�f���GP"�K6�;B��Mi�5Lc�H��tvԌH���M��}K��V�;s �pW���^#b+�����GV�V�}�<e�����}�H�>�CN8�w�I���"����D���v2�ʣ* ����_ԙ���Ч��82������Q���L,T�jü(Y����a~��9�msV��"-ðHC����1f�;��t�sP�O�2cyiS�pCj���~�s�:8Yh��Y�ȅY�"/���ke�"�6I;��i�����E!�a�ʃ'����	�>G?�5Ñ(iV �i����M���1�^D�ٳ�x���}�H�~ULNJ�b�wv#Fʯ>�d��pA�i+��m���i,���"�f-���5y�AՑ9<���&��E�p�sC��p�p���ʑ�����Xm���I���e��+�2��T���ݾ�o�.^�$�7wy�8M�'�6s� ����8v�,�����Y.��(� łٖU����z��怍Պu��������8q%�sMJ��﫚jW^�bquBeR�M<Q��!@�^Y�aݍ�������(���(�����?�BMZ���n�����"�e�I(��k�������{�<�q���g�Tk�ܦ���Ob?����G���Ү�c�K����	#����l����͝��vE��\귟<m�?֯��b*�?J���)ý<J{6�yX���E۞o{��afH��z��^��k�-��Ǌ>S�d���	Ʌ����y�İ���ßkq{��m���Or)N���L����8�E��wFن�V+{�sQ;��m?��*��'~��.>Z˅
Zq�b
1�$�<�bOF�F���>��[U�0t����߫q�9p/U��>�\�S�t���Kp�  %V7s�#�����R�G6~XH�Dv�I�������>0�����'0������o��Z�4$��7ӳ��Mn��z����+d[n�5��:�bJ