��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|ḱ	I*�y��&��U���RvV��>O�lP[��/�=&9$'Hj�2R���_n���l�2���2��s�+C�J�9?;�}�hBXW�z1�$��Z����V,��F�ݨ��"�5�H�p�Ŷ9�^�@�%����I{��"�I
R�R����� �ov��ҭd&�U���{�y�s���;$���0�k�Ϛ��P&^�u|�� <�g�Ԃ��i�v�K�9�#�������_PO�LK%�䦟}�(B��+7K�sWT�B5�67@�(�G�O�%�U�K��˲]5I�ؕ
�Cu��t��Y>z<�%��v�%���)��>�_HY�@
��~��0O� �ޏb��$���eQ�W�s�|��f|J�%��0�*�7�W���+�d7&%G�Ʒ���<v]ܽ�h���X�{��iFy��Լ�e��M���h�;��n*Y3�����
�I�ǜ�_�!w�(Rje����yn4���a�mNf�������iSE5ep87;����6��"���|>'�#��/��3��\���`��_3���x�����;�'[���Hv��Jt��y��;�D�/���A�daT��*=�d�E��"�Q˺,C�$N����m�q&Va`tW��	�DFcҌ aG��8�)�5�����u�v���D#��0��ܵ��Twçzj��T�2��$ш%˄� �N@�p&�2ԪZ�V�Կ�6'���FLI%���1��z�#j�Lrר�\}3O'9+d,VqS�ݘ�a}h���Wd?�<qخ�A�X�e��P �^lO1ױC�t����R����fo��\k��i5"�L���������Ad�~�$g]�yDʕ�&	������EC�;�6�&7������S��$X�4�Ľ��?��qt��Gf�9J�}�o)/2~��5�V�_�2ef'�
������=@<ع�K��^ CTe+(����l��4(ـK/�����o.��'����	i�i�������d��6[�|���e�h)v��\�s��9SZ�b��]rr�.}��ʃE��Ir���R�y����boR|����G˗A��ށ���!h=���Ad�>��6��̻�p{}�Ӎ���j��[R�)w3-&�"��8��vCQ��FA��p��~t��1<����)'\��:�n8�o��D�NV̈́L:p�&��&���_�� R2��̯�~Ȣ"iқY�eI�}���j:�0��l19�q�AN/(��A�D�-p�B3�p�i��,�/�O�������@9$�=O����e����b�����Ç�uU5�U�^Յ�L��E�י��z���	l��}�[R������H��񢌋��Q+��g؈$�����2�����r���W6d�eɏ�~�p����$}�B{ٱ��d���^�p#Ǫ���v���4BBR��+�5�!��.P\���A<=�1)���R2� 5����*w>~lt�Y�>��vv"C��k<��<��=�f�)u܈��q�/܆�(V�g�`���]��x�b�5�x)����}eR�������]�N#�M��r�h�
��Э%΄H�rm����̭|s�sj��΃���~]'�PW'���q]/�,�ܛy�Ƨ´� /��b�H'
�2�#,sИ
kãcԿ:�Z���%���5/&��q��`�He��h�j~_h�{��jg�I�}��H�qUK�ݾ4;�ߦ��KY�f����D��T��2�X��8�;H~!�&�эn�/�{P�dbZ�C�QL����^UzZ�yZ�(�u��߰�s�>k���La�MK���ꪐ�XK,В����i��U�`d%p ��}0k<�9,��ʎ$F\�N�����o��'��� �L�����̀��&]�Q�;�n���َ��7(��� �:#���z~*8vд�@ۖ�J����#o�yuq���
�l�4�j������%�b&w/�'���0�������@���'e��P�& �X��u�g��d0p0�y�`oL���rZ�j���<<g\�<3����>��m��Y�EN�Q�g4��/��LK�ަ_u]9�;����g�'�P�AK�[~��T��h�/Mb�x�T�);=�� U�A��RS �zBo��ǡٞ�PR�j$ُ2�{���<	�n:_-��0|k{��D��Aj��WD����d�W����M�EP�P稜��<�[�u8�0��|��o��=��b|��X[��ϔ���AG2�.\UG��XMD�\ �L��8�n�w���"��9�C�S��]�cr�W��v�5��]1�U�1;|�;�԰��h�|e��V�u����n �q��h�\Ĺ%�oo�U���0��R�g7���k�����@�{���V ��vV:8�}����ҝ]Ӿ�1Xb- �/y��BzQ�d���:k]t]w_ˑ��T���V>z��:��*4�ؔP_��94N2Xa���\!d~�䆐5�P�9��|�������V����+�!.��!����Ѡ���<	`V�VC�\\(7�|��Q��FԂ��+ �
�eY��C����6�nH��?Cz��g��U��p+2{x(|�3>~�$�N� � ;GQee'�q�<��BQ?J"�Z�0�:5�H��+Ŗ��p�ʞ?���%��۠T��w��$�J̻�6~I8�����=��M��;E�ƨ�x#A�2�_�R��'��9���� H=ꛧ�Ԥ�aϙ��V6��!x4�h��Z��h��=7�xU������sqp���M�9���PF'�{ ��J�P��"�4WF|)^���ض�0���t)$%��i��K���pS�4����ߙx�:o���s�Tģ�4��r]z�F����"b���j��I^o^�W�,�f��PU�_D��{�`�,�9��3��]�.�HYv{�`a|?A�ץ��
`�~ً�Dv��7�Hj2Lh$��F�,����?/r��`��$�l�Ʊ�w�-�;/�}|	<�Hh���<����{�o���sb7?]옵1�2�L'�N���]����=���k��Ճ�	%�6�'
�)У3A|#�"9���@p���q�i�2�Y+�Cg�;|/7�e<ec�I.�v�IP��=��Q��a��c8�< w���#��" p.�bD)�A#�v4Y�����Z:� ��	��M�
�ɞ�� ����6co�sc�rZ��H>}*I��<�(f^�j0�\,R��X7�(�ԡ��� i�eK�7�9���jE�#�04�c �D�%,�#�u�ӭ2C�j
�z�,�hݘ.�NnS��]��r�5�kM�6�
�@�lh�]��m��Q$�+v�T����s�܈��r��=`6��F3����!j��pX8oE��|���\���^Z����<�:�0�4U
����|��(6��UC�v�,߻���[��1+�떝1)��45��󽼤ꗳU�U��ŭ[�S�؂: nLi0�֭}<����h<Ó;S,�݀����Я��Ҟ�����8s'�$�yRw�Z�Qx�K;.{�Z
4������s��%ή`���DrOup�,�P)W�SL@`�FT��t1��G��j�7�۪��������i����$۫�p�c���-�c{�E�Ob�Km�Nu����fh�����e�6pGg0K)�v�`0vQ^1<����K����H�=≥z��t��m�ö���j�5/�p���,|����t�����X^����V
�:�B���y<N��c�T���z�m��ő[�	�-�!�	�������u��D�R��5^#�F�k\��ڜ�6�׹���D�J�-��-��㋏n��f9��� ���4�<Օ1R�m�����N����&�����b�d�}����A���Δh���przR ��� g�4vB�څVc�=�?�Y������2v����Q�4�+wpϝ�����bz�Eވ�~Y�~"	J~�T���$�~����6�:�v��h(/�ܲA<���@�~��.yg�騡 ��:��!IAݚ^���*�k�Q����oq��t�A07"�Y	���|��9���s�p�ni�kϘK�L����QZ��^��Cg�,�d�����m���SR��1�>=�q0��"78����j�c#rWg����H�I�>����p�={[E�!�U�������������+�����`v+�Ȝ+�45�J!�Cv�:�7����RW$�F�#�� ����R���Pb5��cE�(���ƴ?�ط��a�(�tl`!緯ŵn������*��5,ҋ���CGĜ��lfV��e*�S�tq3�����\�c�є�B&�y.1P��\Q;S��o՜�r�[ɲ�pU�!(�YZ��Z��x���X���������yL����@��l��ьoα	�X�'h/?�+r(�G�q.�|��'���LQ�<^2K5'�Ai�
�SP�&��<��.䴖��®�[Rl�faAW&���Dw��$��C�c|C�5�O�G�W(��B��
�Ĕ���Q�Ӛ���|�ɣ�Q�B�C����Y�5ς��,�OU�PQ�:���:/��c4���_�m�T��0���u}zǕL�^	��-- 3S6���������+q�Ci�V5���nm6c&j��@���^�+oj���{�zz#����κ��$���`�W!�Έ�~�u�P��u�7�w��7��5���W��s�y9�giLC�V��)���Aq�)Nx��K�g��|0�Miwm������� (��a��D4Ծ{n\v���r�8$tR���Zu������'��[���2�3��ȐE�ȉ���]m7��2s�P����1�����V6��W+L�K���.�ҟ����a��g�1��*J"��۽=������}�fc��8-��� �ߗ�,�R�.�t:��:���.�O�~�ؙ��q����C��҉�g���q���udE�!�h͆Q�6�<�����_���2�I����5��M�i+0И;�r� ^D��υJ���,��~x�_���bTڌ���r���A��;�s7� D�����5�eN�fC/��3`�r�~�ʡ0�F���| rO���;����t��8k]e>��%�����α���d�8K'y�tb�T���<L��d��}-���[�t�/�!E�lF���5�ʈ��ܰ�:���w1mh��Qs�Ux�rp5�q&|�Jl����z��*���@�قOBm0>K��D�/z�H45�H��A��↨iC��<�2���iҘ����;�Y�Z���j�$�}kr�0��:(f��%�<ÆU��ѹ!�gTLS ��}�ϸ��= �����>�
!m�^W��)Ě��C�`(�?��u}֣����ߖ��<�L��<��
��7Ikkh��V�А����e����1����n �t�C�����;.�W=��d8. w����n�-T<K����qF��k�.�Ga݄�Z����#�iސ�?�(CK��rR+�%�
;�G��w�`�Hm��kre?m�LVX�7t��|�Pwl��&a#�
4���g���g1�d�D�3�����1�I,j�+4�/`�^o#�F(V���K�	����*d�`]l9nsO6�HC`�� �R׎#m2��"��S����dԈ|<^!-�05����[b��C���U�l�)��R�6ޥ����Dz�� �׆@� �4��Cۊ�>��g��})�զ�)�� ���c����ǣVlml�_���g�=R��"�'�:���8t�v��HW;��_�*1�l���+Y�ũ�6]�����-�CY�; �s�s8b��b�����  �0��i>qxJ��&W��6����2g�|�z}?v�)1�m��FE�|W"mBg�(�SԳ�4�����Y��w�jнPݰՎ>p���1F[ƶ؇��������,'�kTx��2W]�16ң�\�k�WFѻ�zn=p�m���\�pllyF�mxn�"B��w����o��`/�c�಄	��������?�$DЎk��!�_�]��C�K��P.�|x�$�c�7�к��J���#�vk�Z�w3P5������ J-ڴC|qv�q?Y䅝o���(�ׄ�	7ͯh�~��=�K��y�̂����}I�_����!Aҫ��^} ��=B�p�-�D;#�C+���{�ϧQ8� vUH�4�N\B�$�����s�+�k::[��|׿*���ȃ��H��_��a:�B�6��9���$7��ܟ�`wS���rB8�KҸ��
ϥ�>�E3?Zu�������p��u�#�"L�I�g�7kI�D��G�@��
�����޲Ew!��Mۡ�劍�O��&F��#p�`dWcpj�]�0��w���zj���>��ج9`���3(�D�}��9'�������o/A�����])�%��ML����.�mQ�`k)"�(c����L�z�:]��]�
�Y�Cʹ�����d�%���FF��d*�w$��poX�V��)��~��A��v�*;|Uo~c�)9'&���u�]�0%|ʁ��d���1Ũڑ���V������0/�P}�x��3\�!���� ����N��q��G��v_�����k�g�$�`a��iY�ג��I����(C�7:�1 ��z,������Aq�(~�[؍
�ҪDH��M�H�����;McC�!���E��:��\��0L;ӃI?���H�N�9q�VuY���j��r^�J��]��#% ^ƻ��;�Ù\�
Ĥ�k�5�-�L� ߤ�#!~�WeLDW��z���� �p4��=��h���ü��F24M����M��6�'��Ӓ�iC3�N����b��8gp�!��{�_<�AJ��!l��Y�fМ'�K�-ɓ��Q��:Vlj��a�d�챩�yޣ�=�.|�F����O�����b����3�]���!	��<�X��k�B�k&�pёY%#�z�š��0~�O����B�XQ���IՎ�؎2M8����:�4;c����3:�|��y~�F���5���|�u�ix8ծn�7����g6��S0��Iq��21E,�v��4�躩dl�Y�'9Q��T*��Z޺��_��I5;Sr�;;t;$$�!�/�N?��(OܴU��G=�53R>:�p�(�T�/�M��x�Ŀ�s/u;{y?��F:I/r�u�W9�H�D��t����@�-�0�{-;tt�Z�������P��ضK.Lʒ@�4�
"��V+�Ѩ�,�*��ȁ6�˸���>�� �����w�l~�1����~�����^�nb�	/"���=ޒ �\i<�1/t_���OX7�p��A�~�.�+Z;Nhl�I��戝oy�͗�~ѢQ醨6;������RL�b����e ���ު��6��|��_�9/eޞ�Ԝ�y��f%�2�T�J_�қ��H����ޥ�~+�Y�,�K�F��!���bϹu�~Q�E����u"��U�I��[w�E�Y쭔�
{|`�.��[�db�]w���S����9<�<�p��ʷ����z?��@8�@[�O�y#���y�+9�3e�+�ur<��� ����bm��Zfc
���uܰ��iڣ�� {w�e�o{���8���,Rx{�?���C���I���{��Jn��\��i��e0�E�h�tUJ�E��V�g��n�X�Qȑ8�@��<��G�,����=!'�k�1la/2}�NOpYKԄ�z�Z��n�˅�X���[y>��C��Y�:��$��:)%_NF1-y�m�4=�z�M�l�i\V�@)V�Y�h�DT���p��Z�پ�T?��������y���!�יg��]�2����=�	h���5e�����R�(_�؛�U6��J6w$��|�03�_@�#@;*XFN.U"2vK2�S�WE�������T���Oja����u�ljQB$rǉ���#z~����s_�P��1_說���������A�:�R㉝��Uy.*��ͅ[k��&� e�z=1w#�O�	�>�鳃����#S�@?m���ԉWspH�����kK��nc��[ƯU��r>z����
�~�j�]jx���`��uG �9�6�BpuՕ{�0��G�	M�8��x|,U2��]y36���	B��QzRhPB��[�gY��K��c/j������g�Vx>�v�M������4�� �Xܼ��P�t"Ep�G��p'�����'V��z%�����/��6��N���ZC2�P��p�3y��H7�{���������sV5���Y����ϲ�� ��K!F"oX�+`)�*{g9���<��ZW�fֱ��]m�.��PV����?�
r
�
pU�f���˔�\�G�~ZJ��#�l�z��eg�����9n�j2ɒ&W[�i�!r) ҹ��n�rO����⹄�ݜ@$���*��h�ɮpX���K�?!8[f�Cy*�J��=g�+:1i������Ҹ���u�1d"��y�%�ѫ�ٜ�AK������~�ԀY���~��ί��臦k�I�O@9�� ��wڼy�P�"=}^��,_dM�"�版mc{f?�����Gp�F('���_�q���h�Q��%|�-�v��jTG?���F��.4C��z�S�(}E_�����S=4i��
	(�Q��a��W�I+�$����G���h�/>��"���b���SI�J���.۷'J-6�K�J�@T���i2�)Kr>4-��1p����]B}@�.��Y�B���!"K�v�]��5aSI���ɴ���	+��d�o,�n�@�/��Z��f�~.{Ҡlb�sm/�j�������r�.��ɇ|'7�|�XW�FA�t�,����M�c����T�����
z�e9�1��N�p3�.Pkt��m���76R���?+�j
v��iV)L�m��M9b�7�-��3���G�Me�0_
�܅�3���D>��l��a�5�"���pl�a�[��'���a�@
EW�c���R�S;,��ADX���j���$�3�<�V]E��ʺ��4����L+΁��D��>d�M4ৃ�Cu��^���9�>(�zYʯ8PԂ�Զ���X� �Y���~/3�s=�4���Mw�'>�[��#��@�l�ĉ�1�^�κ��vΟ����r�������G��b��Qx-zy1�etx����1F
G�f�L�EO�/:�'AW�xm�#��9�$9��_���֙��,c���6����û#"�N�Q��]d�	�[�H/k�4�~R;g
��\����S�g<����p�
�+IEY���[W�$kW�T\e#͓�O���rqD���-�r�@��C�D��hW�b<�{�X��S ����>ф������a�uţ��6������Q�*��ݦ��(�̛���6:��?ץ6nΝ[��%��}38�;�s���f%a�h�T?�8����}H�*}0��u<$�z:p�3��?�bo����Έ(F�8⿴�^c֓��K���� �7����*��]�!���[�y ���&����*6i*-uTI��?����A��o%c,���cP]C;S #,�7��M9��q#��3��?tr>��f_Em��)Iќe�X^'_�*���N�I�v�-Jdr̴����X���0Z[nz���Z䱵��'LcJ���7py>���s��[�1;L�;s����#��[��M�3 =���8x���}͓}�� 	q����rNS���BM�vE��E�S�`;��ԫ��Ю� ���7y��B��X�ѷ6���1�7���,�1;~Vj*���/�����v�E��cf���A�c~�h���ul���Az,V�ߺ���Egt�����e!z!�ld����g��m1&(�9l\�B�`��Dd�Cry�Gt���·!�N��|_�-H�3�Mz��d�xd=]���}�9���i�|s�Y�{^ۙ�8�,��4y�h��E�Ww�u���L����K^��킪�_�����f(��)y�KH.)�E�{6,-����L�9�aɅfs|�)�M(1�R�^�=��F�k,'HM�5�~]cݷQr�s
�On&C�Zm0.�X�YFF��L�����p�s�Dp�o��l�a�.no��T�����Bc敜|�Y���8�$���b�v_]��3Q>�Yx�,Xz�8�X��"}j8�Bm �Ki>�;�$wB�Ū����I�D��UŰ�n<�,�I��4w-`tQ82��|X?L6�]�i.�0��z�t�3���OM�GA'�Dw��b��Qe0֕T'NI�B��H`ɞ����%4!��!4l��Z1wp����Q�Ch:�\�F��E�-#Jw�{N��%s�o��Q�j���ϤG��&�c���F wn��1���WNqtDsm#��,_��=ˮ�8(��YUh(?<k�l�����jǝL|oC���3��2�֦x�������y��Ҟ�P��	��P�vP���9y�@(TK�.��� �ʢ�p�� V��r�V����0'��Q����;_;{T��栵�Dn��ּ���oّ1?��15v��<&.�]�b���|�_��NO�n�g2<�F���zY&�lH�]�(�/ӻS��A�(]k�q5�-:Dw�	�l��9e���~�bB��ꢠ��7�s��w��+�|]�J	V42�,uh��a���D~ޑ� �8�ټ���hK�|�Q��/o#���od[��#��M��yR��6"PG%���Eb�b�e!_A�b� �H`�Ch x~s�؋��\���Edl�b��0�$�d��������U�wY�3�/��0"�"O��c�=)}n�dH:�����Wqv쎇����`�n��xQPt?p���kH���T��̋����*y�:ݤ�ވI�eosY���K�En�s����ΣHk��bыOBL�h�+
̛-�s�E>��ݳ�c|���ō-�A�� ����D�dB5յ��V�z��]By`�ҿ�̓�}�$N�F#@��n��x-�5��A-���6�Ƃ����_�s�wD�FOݟ`��_+E�I�<6i8���9����6?���Zu�F�-�{O|�ӹ�|)EJϯ����<~���Lm�mj.�ܜ2�o��~��!Et!8���\X�ҵ��GX|�PqlM�k�w�_=oQ�x-G�(�Gh,�d�K��˥Xb͓vL�ﰠ�f��P��+��WT��m��	�(���/n��Ɯٚ��#<�w���ms�����`2�!4T5��,��mf ]��˂؁�U���6�O�z!�
{���.D�A'�B�Mq]|���i�:�|7['���;�`׆�aJ��s� �1�<0�^+�����2Egp+\6>���i�c�=*�!ߵw���ih��M��S�\�+�r\9�_�p�$e�n��<��������L��'ylG*��:zpB�V�v��\u�<]�[�0&�ϗ��7t}�o�u->�#a8JE������n�1���=�����t?��z�s�Ź������^�2MS�&�8��n�ts���4^iԫ��.�fe�C��Fa斘��&Lm -O�K�������E�^b�ݬ�IZc,�x��x�>Ŭ��C�o4&��f^8�rnE'|!�G�4�6��QP)ݶ�����=uE#B�kEߏ=5X�>��ϗ"�%we�z'�>�0S뀱;�@	�a��l���0_��y��_8�7��5�2S�\Q ����KYƫ�!��l��?Vq�2v�K\���Q(�Uȝ�z��}D�6k�p����,�@�ֺ��U�B(7&(l�KAP�7�#"�4G�TX��4� ���G�l�_�m����A�V�����r���s/~G=�$De��B4��aΧ�Θ�~?��D[�Å~�<Yz��� \��b�	�Pup	~g��;�SZqbɠ���;NL.0�h�C�Vi�sZn���O��uRB܄��'�gϤ=��ճ�T���9،������5B	�R�(�j$�U3�p�_j��C�,�k��͢�+�C{[�e{��v�����*�`���5J�c�f���b+���s����m��D:3�k�4m������~#@��2Qh�xJ��0;��Nʯ�i����+�o�i8�/�-�z���_�&�3_Ff�v/���'����aA>Um<�
}Q���4���*"�3K܂�=;�
��Լ�Q/�,����T��S=�/ī���r���U��e%�5�4�rV���S��z�ި1�*<ۘ��j���D���+��<=��Wt6D�%��ҸoS�,Fx�����'U�sqg��Ѝ��O��)�`o������A������n-G_��w-L��T1�ID�_*�����������
�.�F�Sh�L1R|�.�.�
��$�����e��:^���y�T��=�����xh���)~J�UG���m{9=�p��p�6� �v�ǅ*��/
s�y<�P�N����V<�hT	T��n�7���z`���o���$�_Vvk3YL�X!DJ��$WQը�������\w<����^��^�{��dG��^��RҒ�)=T
k9��y1&"M�~ c��*R�;���!����m�4\}�v���һ�����6℘Z�X����)u�@({CIXE�l�S��c{�	K3fds��E����u�ǳDa��i��5^������2AM"&���>2�����y�N��s4>���3GR��/S}��ȱ�LG^Ig��i�v�zO�WK_�5)�kW}�kZ��Y]/2���8[���C/�6�m�t�fm�����A�1T*sݐ �����Ȍ��$S\�~W;!2F�6��IJ�\����Ӗ��^�p�ac�Z~�Ŷ�M^KE2�wս�L&�#�rz������I�����_1.��&���7�f9�ף������.�Yg���c��v�$*�u*�do�F�LNzTA��U����E� Zz���9����Q��}�H�)ɏ�Q��7��Q�`��&(�mI�T^uƣm`?�������}���H>3���6��"Z����_5��_�D�-(*���B�zU��b	�4]w���a�"zLX8k?Ns���$�V��sD�X'�Λ�@�F��[���O'"�qj�B�.K�JW��<�"4��X��Kg��2�ɤ�J����mR�z�U�Û�������u�Y(�zo���1(���j���Wr8�s�����\'%Z��
�s`�1���V�� S�Mk���lU��LS���є ���果|��%��tbڱ�B�K��A��&�k V]��3�Z�ʳ�J��Z��W >@BԘ�a�YD��-��v|e1�pV508��`���7}����;G�r��~{E2���ȼ��cMB�z�؟�5Q���������!߈�u���W5��Z�O�ϋ��V��/Pү��|�ҫ:��t+$��B�y:z<C���|�ˏ�ŝ���6v�%��0#��?���9���<Ă�y1��Z�ǀײݣ��U�LHИ\�v�h�� ���������,h�K
U'_ۗC�0E�zWÍ�Z^��1�5Q6t�-��-�2bά�Ԝ�N�K���z���>5B��qH�ՃR ��´���d>ʲ��K�E�%3E8�zdA��F�C����V��T�-�nC�s�� ܐKqE�u����nz�dt��������L:lky���q���b��^�m��f��gnA)o/y�(�}��hЛ��8��e��8��9x���aF��Y��&B����9�h�UwG�������J?��}H�q�/��K����!s׶BТ����>n���%	�,��=�JT2[�R�ζ���9��Ь�x��G�=���Cuo�������g닛��O܉���L�`�@/
��Шb%�~(���5��O��"��0��K���5�4ܿӮ�U$	�>�Pv~X�٣�F���=y�(_ݒg�qx��=��-��R�W�5V�G��UN䪧>�
^��䊨 V�����;��G�A�=@��X�]������~۴4��N4H5����d����l�G�p�1Az�`S���!���/M>��OJLz����w��J���^Rlh��,�?�x��PmiO���W>b�3e��a��+\�EP�����P֢3A��呀`�rTp���}Ǐg'��${M�~lj��W}��� )O�W�O��ָW���v�}�K�)�MHy�~B1�d �gAV|���'���@5hX^(2��/R)n���vᷩ=�J���n:�OEq3~�_��+I�����n0"¢�.�XH��-��w��u�.wӝ�^��4PnڅO#�!�ZmC1�Oę�&�|�Ġ�f7b�;-C�	�<����ʢ�T0yW�ɨ���N>~���N�Yj(=���zܥ�u,]�`�/��k�)���Nn��l�pu�(L$n�:i�si�q\��S`{�\>5K���^ 9����E�r#,_��=�4`�fr�`���/��0����ż��*z��;�����P�Y)��NMVK����lXJ���?ݔXq����(KJo�����,�K�i��K�!x#L���b����yϸˈ��
^zLĊ���O`�y���s+�@�L���������5�cx5�����Ę��_��C�45���N;,
Q�8�5�RE�[T�!��Z4�N�#�t�#�g������*/R+D�M�F-0x�j5�!�`C|f��a{2�!�cw�-��d A�6^��X�-22O���(�����q c��
v���k�EN��hH�A���/�e��ȕ�=��t�'x=q�9���oěI�v'gࡘ	����w�$(t?�H�7I=X�ypVr��Y_�����_f��L��%���4Ώ�����ķ�� `�T�g��|��dG���Ho�L��u!MC�hko��6���� RrC�;u�z�I�S.C٥��>S@��(5�"��u�4GE(�vC���Y�4J�3��3m��yU��\)3?+����p�����[0���+q\0���h�)���*�;�4L-�[S��q��h'q�D��0����1i�<|I($��ڶI����g��z�ʈ�Ճ�s�K��,;�:I��Ŝ��%�U!�<�����h/�0�6huDLP�gP��\�}*<�oak��ߍ�=HR�y��5���_t���I��'���~�_���p��h#{_�챒��Z�"[�g_���T� ���4Xu|!r�~�>�mo�Jh�^B��¡M�U�E���Y�KYnB�j�J-j--��^�K�;��w����&��ȜMp�4J�j�ʜb+hN��5XA�۩�	B�˅�I�@#φ�h������C"�G~�ٺ��K��@����\{_5o���.ȍ�;@)��,>c{����"�� ٣����#�-M\�B�n��(%���%���,k��?��XE4�\�[J�A��VyQ��^7c���բ����Z�.����c_kU� J�8F�Ѳc�\Pͭ��j��J�r:oIe���M����Kp����on$�qC���yn���u���m`��&����Ǵ=����X���Y����6�ܰS����`%��[��A�w$�g��5GDFË��L��'�f]��έ�U�]'�J��j��W8F�� �w�T�9;�q3��E./��6X��݂�wc�g���Nu�E\"&洞�����M���7�'C�����ҫ}�gR���mY��Γ�G��A�W���.�B��Z`�0�c;��ߢO�Q������:��2�9�|Z�@-6IA�Wdc��a�5>E��t[H�]t�=Gǵ{-�P
4��*�/}H U�8�?����,[�od�U�@>3"񵟵#��JOҔ�SH4�8x��r�IM��0�������Ҩ��ZP5Fa���^U�$�&�����jX��jȎ�ˑب�:Y���$-ѱ�Ԑ����-:��"!7�_=*$��HO��|�X�RTUˣR留�����V�p1Q�k詬V�� v�|4��O��0_��g��5�hT�(���R��	�g��H�;�4n/�(d�SJj�4�W,W���(�z�����q�yz����)v�r����04�in�|��`9*���#pU�z&��
*}�����H�N�0��dk���)�*�o��؀���*T ��|tf!ȶS����K���vȌ����u~+~��ɠS�`.�Y�=��:_I��H]��x��Ǯ���go~!�����vC�
��+5�Șc�F3uy���(JV�&"=�D��(��0�>A���>��"�t}��g�|�5[N����T*�fx}k���+k�V�x5ϥ���3#��A5��+0*�`��",I��-K�c�ک2cl���t
�=���=Q�#/]���Ep�\	�D�;T4�ݽy������̇/��^�1;���>���?&x��]�d5H/:���^0M�$6����Q�P�3���;�M)�pG�D��/|C
_���|%��ܚ���gHt(iK�6�%IY���gH�Q��ە"QI QB�,tm� 
ONi�8�`Y���ؑSY����,o+��11E�ǎ����sy��\��+�AR&��9��(Hf�6���lO5�*���[u�����i���C�'��������2�`�K ,��ǐ2M�Nsߗ�K��PN��Q�}�Y��O�,��+5�'��_&/9��x���#�C�,�-q�R��@���<��W�\���Q}n/�=灙ըojO��6��p�7}�r��a�qٽM�g��� �[b+��¢E�	�Kt�"��� ��I�����0�/�6��ʇ7�tv)�x*��9�����_U�	�]��4?u
.je�p�������CT�ͭ�E�_v	�i����CVBn
F�
?�/Z��Ǚ��T�\ �,+ π;F	�E!ֹ��)0Z������_gru�H�'�`�l���;�"�X�	�+%`}_C���7~����:�r �/#���,y���;��x@;��6���	�-�Y7 �=�1s\�
�I�C�S�E!�[�~�.=/ߧ�@����]R{��½�t�)�[�������2(�/p� :�b��������̈�k����UKٗ��O�`�0���4w��龷$.dM����^7��0�W[:(ew/�0��u�0�J�+�Q�Ma9�Ǯ�RYt��/��n�5C��"�lF���H2�c����J�G��M=YE�uڽ	&Ӭ����<�\�ǳ��{z�l���FO����]A��TF���I��Y�T��`�Ǧl*O��6ʲρ�]%��E�6ҼL7[����g�7W�܍s�y󾋫�+E��	�1�FYiT��)p���Y ��P��`7�S�����-q�G����eFs��?E��\��#>�R�?I����T�A3)#�-9�U	��sC,qiuZ�}��ݽ�g �V�A],.$�Δ�N�$�� ����V��0)Sj�S�X����a#�-ֱ�ax��7��	I:���Z�.�y%s6|C�ʴ�[��46l�W�x��Ż FQY��w���;q�=�I+�m�����c���z�6��R���������(�k�$��.�!Ӹ�Jk���0���W@�;��B�Z�C�������r��{��u��R	�g��/�����'�g���;�:��g��{�l�ӯ<��V�	�[�Gn�����xU3����d:��U 31��dFrw���OP r?�l/���K���t�w7�9�t3x}H�A����X�?�r����ZQ�����~p[2z�K�v�U�J��^"�ݏǶ�2��anz,�s�_Q=;]@�2;��rv٘t�ۧ� ���JT��bdD*du������ZY]�v J���S�0��x�[�x�k�"ByK�im8��+:Ӎ�!�_����3�瑜���r����dkY�p�p)QB���f����wQJQZ�5�vȄc�oܫif�­����'� }�C�K�os��8����lk��?��y�@<Bj��&�W9�X�f��D��U���� �~�iK4<�ە��-�2�o'-���~l���d�47X_�Q8m���R 7�&�1+��`�j��7x�T��@�J�s�ȿ*U��=���h#( c� :,C$�m(�޳ڸ��f�	�_�v�^8FۓG\!''��脄+��n؎B#��Q��B�Nѯ���L\<Q9V�n���؛�$�,S�n��Zx܋��LC�8�9h�g�)��))��r1r��
b(N�#LĀZU��{+�T�����#��r��� P��
����4a��5�7e�������l��%��8K���ŁAZ�ۿ���EE�g���57Ѹ#��0�T�Oqa��゘J$s_MOr�$u3��aH)XH��r ,�	{tT�}�.��!ds��m�jh���{� �E��%nw����ۀ�&Nx�A�5A�緇xLt��y�#�����44�%��/�Mk�]O.:�݂�����ԝ��mB4e.	`Vw�+D�N��aڼ�I*��/d�4a�0w��TlV��U7K?�g�A�W��^pJ�{��r��:�T�Bs6_�wkBa�ȳ�o�P(ï���lw745sc�8Ǽ�Ys�-�ђs�^�v��!��.:��^hqc��P�S�E����WAS4���^��a�5t�2�(	���s�@�y��$lv����7G��i2�ǌy�k!y:�ѧ�B�Q��B��Ülډ��I6�8�Y,��耔��6��v�o�du鏛���Z��^R�-�˙����X�c�_�;h-�:�x'��V��BA�>̳ޅ���vi�BC�XE�W~���K����d9f��!�bR?5
��x�?�r\R�P�IMp/� ��A4�+��%��!M�|إ녙�J���g��3�r�CX@87��	�_��`��40�Ԅ��эmk-e���b��� �NN $��r˂b��݀[m]��M�.�n
ʘ�p4��a�����.��5H�7����Mw|��ײ��QP>����Y]��m��Io�{�������8�8-q<�nW�X3v���¾�{7���߾���H����ƨϓ�]���ͥ0Rit3�+V���V���3j a�n�Mϙ9֎�$Y�5_��|�3/�J6�t�V���zZV���s�;ַt@�����;��h��B4�����)~���S=fp"f~w/+i(׹;��^7������ly=)e,�Y�RBiI���p-��0������]LF���G��R����L�K_��ӡ&�e;HY9�;�_4Z���W��(�qQ>B񐋃6{��+������_LӍ�-[Y��I�v�!��@���J��9�[>X�f%E]�x97�d��Y�\*���a?Tr�L���G�=���C[�lh�pQ���������Qs�Tjs>��4�O�2�M4g �l�j1���p)�}3�����f�&X�
�3�A�K����}�(8��!+�aC���R{>�%�����,F'�P����_;�ݹv*d��<2����H�&ٹL�\�.�A��3U����b�1~jaX]�`g�G+k�0T86��5J��L&3{���[UZ"�=�&AAֱР�*%���%�~��ϵ���5�RD�RI�ܹN�mJ(aV���|�u���ry"Z�f�${��C�I���|��1ن���U�9o��J<�V�	N�׆1��6��''�����aЂ��kU}�9�R�����K��Km ޫ��|�Uo�/���:��]�VHQrI&$F�ڟ���ߘe0L�_��>M�1��nU����}߉�iO��1�Ro1mޢ�<cL���y��H;n�;�[�_�c��e�-�A�̢�Jq�F�bj7�|ſE�CF1M�,�%��>c-��a��S���Xq0)2���\���~L�a]*��Ө�l������q
Cɵ��ӭZ�������������:��o^�r��s�?!�+n_L_?5�(�k��ޛ�ڛ9���
��0����	��y�o�_�Ȳ4PA�%@��?���o�F� >2���ßD�d��P�t�o�����'���k|)���P��s���ƥ�Q���]`F9	%H����H�;x<W���T��iΛ�_:䃸�)��M�:/��G�����m� D[�8�������*n��}��R�`=�s�Zr��_W-�ǽ��qS�����'�?�"���BVR�Β�[���b���^y�����<n���?�'�j�p`	}�i�Ya �3���Gx`�-����M�rj~���-$zf�����SV��Z6�ao�,Ύ}�O��G�P5B,�g����lF�������q�JЧ�&pN]�E����r[%�f:G�Նb�EXcW�j�:����ط��fh4���t����Rmy[���4��8�_�a�ܷ�.G���Q"mD�qʽ���v�FϫFG��V>5�B'��Fwm��������l���!y�5#E�ڐg��ix�lA`c���-��^r�#+\��}6Fʻ�Ր3���X��Gi�j#VS�WRk��~��\�-�5��{��*�\��|t,����˯�zP��dU�D�Xg8��i�L�:2����8hpj ]
�i.��K�{�MPoLڊ��PyX��N�Lo�G�#��K�3�.(�'�ԳTΗ5pM�)����:��|<�(f�s�� �j�B,TLbo!�����"&*g�,#�J��}�W�ԗ�5��VШ.e��u��yN�T:��z�����إ�w����E�=Yw��jX�W����K�>�Sň�(�I��H�H��y��wݑ{��;:�IG/QJ:'&n�R���W���p|~@Rm�mk����F��Z�e3��,u�"Wo�G��;�3v���y7 ��8�Df1�m�����u�i�S�a�B}R�$��:���S�ޞ���?�ܮ\-W`%�?����7`��'#}G@OKj��$V5�}���X#�4� =vj��V��hMy.82'���*�"L���YL���v���#��C��Ξu�C!9��N3���g���M��H]�@ �[�U��_��sf8���C����"w]��`�cw�.&�g�:���Q����g�[�6�o�g�1B;���ᱲ>2���mb��2�v��s�B�:���?Ќd2���ҡ}R��jPS,��͆�􂯈�K�'�-Iy�J]�i���|����j�j;KV�p+"��&�W|o��L^V���/�k��zqܙK���G0M�@����� h���`���R������-QiY$�����}� ��e��vԘ���խs(sy��g��@�&Y��6OH�C�{�8�5�~� ��^�'=�ڸ����p.|����Z�1�md
�=㭅?'��}M�|X��g5.�g��ȁ,iWD{��Ó�Y..@kp�ۡ�0�W�U!�B���&{^��hV��%���$7HiW���=j�o�cD�����B/����p�b9�j�&F�h,%�B�}�/���_-Z����1l"�4�f�z��=ӷd^�M胞�SO��\ٚ>l>É�{5���b��YS�ml&M>|��r���%�]"S����0�0 �����������J��ɭh7�8$*���M>�4��XxY�v�"���t}��\ۻ.���Wht�}�W���A�d0�� 3��a�h�<�z~!���aûT�ƯVix@�d�KJ��F�\7�Ȉ%��1=��&/-�4^�3JJ���0�Rm�VV�C�{�����&kl��ۢ.B�!����SZ�J���h|��,9����O@����|���/����p��r�}(�X�^<�Z�5R���}s���U�f�@��ɥ�;$v"�eq`�;�{��f�X.���q;x��c��>M��Y��-�n{���d<���(ED�	��w�uM��B��=1Y)�;����9�]�|C�V��c�㊇h_~���ȗe\[���M�%���ں���t^8x%Q��f�y>ϮN�|��qSz�vu�A�y+5~EW���`�l l�\&$�˃pȀY#��4��!u�Ș
�C"�g�s�2��\��{x��� ��f�!{���ͽvǊĳo�a�G�}� @N\����J�1�|��p#�#b��x:�H1����wql�MJ� �$�p��?�c��!�Y�	YcP�pOdB,"�(���S�5��(��]j�\--��A�E:��nsi�OJ�Ή$���~��3�<��B���*�@1�3t�'��w�