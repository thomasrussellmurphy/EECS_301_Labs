��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\���V�fnvx��ÍG_;�ȅe�~�>���9�>��Y;�0GW�=��_����lL��*��b=yE�uy�^ĝ�r������}�����;��� &>E��Sz\7b(t���pB�5�xm��|���I��{�qr��ó�s���U$��|�܂/68+bl��,��1-@��/X��G����'~Z��{m5��y�5	xz��ݚ{�0
G���:{��7�]�.!4���[OLx���P�~��=j�I�렿���*`}z�	a�]����U�x�]��d�D�\�Ou�n�|̦f]�����S���4Q�N�':�/H�g���FH�l�e��'@�v��9%�2���ͿwΕXD�o��%���x0�Y˯��Yv[<�Z�@��P�Y�2r0r$�WE�����)�Nv���Y��X��=1`wl>6���CyW�����8D�e��gR�c+�����|\���ЮV�H��ͧ��:t�{�_�� &f�ls��l����#�� a�k+X���x�_)G��*�ŗ;���}�i��wx��2}����`�ƳE:I�x<����dħ�د���T�d��x����^ɂ����u�E���H=��k���t�h�c��qhф*��sN�D�8j�봍+czd��ꮙU��	"���jD,-�\���瀎��^�����g����j��n�F�(o�XF&�G�|y��\��}Z��u��8��u�T�b�}���%a�g�po/�a|��#�]�=�
t��� =��� ����g���[Q� >A�A�/89o�0S��}{�˅F`Z]ٺ�d뢻�ɗ��Ўn0� ��PB���Q��P]I�6�V)�C�(������hE9���S�[�U�%����
��D�!ִz�� �T�|T��a���7�>�i�óXk����wl��xp��� �a FG& ��g'ng9Y�QKR�v����a�w��(��k�T��h�uO:��VI�}���(x���5l?�G�s�۪F��ػ����B���l|$����(+><�͂m������0We��;�\�y`�D�m��ݎ�"%��)���jgD%tQ�+X-����Lw<�ź��,�eJ{{�#��|�+^���GܯжI�xq�6�BC�_�Hؽ�����z5��늗����d�<�����N�j:F��dt����H\����#��u��Wn.���Q�NZ�9��ja||�}�b���`r���`p��	68|Wǐ���+�'�w۾n���S��15����
��O@�#���[��8r3E������E�5j�O�)�£�1h���r�jV51�6��	�:�瑙?b��F3T�� _v���	�d��tHk���7w�#����)!�\~�%�oX�ۤ�4vס�4�Rڥ:0�r��(}	��V����ĩ�����RcY�jS�� b����&�#�Cj�Gn����'�S-��m��]d�3G�f^��Z~WE˘Q�߸�
������������q� ���Kw�Ǯ=�8u��h����Bl�W�a����6 x#]Ōw O��,j�ݧ7�  �",e�b9N���Z|+I$�"��rK �n�%D�^؉pj��8���+��xP9�U2Έ����,���4��G�#���	�7�o�����^�wq�/�؍T�.�),S0�v��ax> ���")��ᛑ"$.}�k�='������AR��=>��Xhd�Y% ������+�Մ�����VV��ߞ"K���д.}v`V�Z��KB���.̃c��֥��nl:�ܠ���Л����ě�3n:�.u�c?�����q��X��;��{�-�HM�H>邽<{���h�^zL2&'�����7vz
�ۍ��)�|�Lq��b��\1~�[��R������[?��+�iZU��,�t8C��}��rg��&ip?�����z�:x$��'�{x,����_���zr|����h�ܶ�ܜ�ƛ���z.�Qg����!M㼸nV!�X����Ӊo.); ��b\�����Y�9��@o�3�H��<���JVf���,�<~B��z�*�Ń�
X�S��\G�|� �� lv_�)\���DNi����6�/\�G_�����%a}��k���,~��5�I�Sb�ܴ�H�@�s��� ~�Ax��M�F�oJ�1��/�zPY��㰓u�K>�{�#O�Y\�a"��Jf�~�'�Ug��|1G���|���D-�੖����tP���-�YđWv����j��7��O�\`6R��;�a��e�;��ߠ8Zy�8�@�؈wN�0��7�[�*���C\_��>*�����>�~z�R���}>�^Q�I�� 7K�SsiM�V�%�i����z��(�م���|��6��i�J]��?
T�
���h�H��;��ΐ,ࣵ0h"�n8������y��(S�H�Z��lͥͩ��t퇳�(��z�u�#u��������:R���; �Y��/x&��Y����(���Lr��5-w[��j-��x��K�TC (A1\&�%�Әr���2��u�Z@��fKD-�ep�,��Pn�W��S���~�#$�gvu��mbݪ�hIؕ.l@X�2�T2I�y5�0���2K���#}(8m����ȉ�j�=�e���5�(6��b�ݵP��oݿ�
+p��ŴKMQV7"R%d~`  ��.�gR2��[}��:��X뎃(.��C^Y-��Y���w�C*G�}�	�z.{O��J�Q^���x� ��Y���c0�n}�Q;v�M��5�#9)�Be:�����h?.б��X������g���2��_�G�s���B�d]����V``�������@͸�\��w%!Ar߸�/ ���Q�&*S�1�럓�ta�,�W=���?0��m�O�>Z]���p�A��ٸ�A��A񳇼{���ng=���|u�NaR��"�v��m�~;t�I��5ߠ�̘��m��{Fy�q�Fe��w���4@8 EIJY��Z,�����vU��&� C�T�TzG巨�	g��
D�WU��E���:���9~R��|S�J?�r��z�*����ك$.��	� ��n���Ͳ�ClL@1�����8ۀ�/���`����,=ze�L
�Z�o��H
V;��y�%�3p�-��m�ɵ������YE�c�3BH�<��(�}�,��.�8�>�����Ρ�����\J��~GP��@'�����S���oy�ɗ����#yU����z.���6�<uV�����kQ�#V���v�S0-A�.�>JB�u�v�y)�C���3J	 t�w����F��Sb��p�����}�5�J2rz�,�C���T��'*6���+�S�'�����SMe��o�_|��b����r?_����@� @��]O��ɶ�R��	��}��"iZ�A�M��|��nN��S�=Q���X��a�ڏ"�D���"k�x���3R �MLs@����S�z�xݗ�����W�j9��U��Hj�XOQ�����#mO�I��<�[eXRw�����sYb>�'�H�S��8zi/�Jy�m�%6���������1AJ�Ŭ_	�+_�2��P�IB�����&῍��Wl����)�%"��W0�R�.Ȑvr��Q�m��͂��H�;��O��<�s�L��X�o!�yE�[�J�6m�ﺡ�;S�
q��-Rl!���������K!�U�pK� b{��K�آ7�"����P�O[^?8�s�Gsh|WmC��١�����.$]sZ��6Yؙ'SF�S�9���O�z� ���=`�Gקa{�,���q=q,+��\��DJ��n�CD��d�(���H&r)�7��0`lw��ь�F�}Vv->�+v1��ձ˚hJx��ѕ��kF�H�Φ��dr[_���Ύ��d�N�J�7�n^r���_Ī|�OIMT� u�M#@���ג�>^`��G���29Ƥ��Ɨr�X�o�8��ҁ ����Cv�:�ȁ!��=0���My����o��bx�Б,�rC�m1Ed]�L#��f����ȴ��n�+���I{u%k��I'"��F����9Y�t'��)��SfɅ�1Ρua�BP�1����"�%��=P�;�%�5��C��" �_�u��=p]��HGS�b;,�J2Yb�C:ZoL	|�9�������^��M"���1lv%]ĳ��s�B�9��b��l7c�Z�g����r͎�3���/��"�!�bKn���L�x�Z����S3۫��p&��x������C㋝6����5�u�'PL���{
��ͩ����3�����g�IE�����Pʪ~�;_43��>oD�ж662� v*9?� N��}��ۢ�~0��g�j}6�$�KB��f��'�6��e$.���XA����Լ����P1���B�̣�����3
p=�q�K���������ゼ#�3�����B��]�%�N��=�&'�'���&�|�Z����O��qo�30�ZB���:8:S�9�J�)ykff9ˌ�Π��$�j��}�7;�T(�O����*�t�?��%�Τr�x�Mn%)/���K`Axд��ñ[��H���BIHri�t�4g�-�����5�<Ԙu�c6�\�ZF���32����I�V[�!(��b2�	 ��Ҧ9s���l��ꗢt�(�?u�x��*�r!
��8l��jI�}�D7�j�$��޺�aV�0��M��֘�q-L���tZ�H9�}�ꔌ��x�hS]*��l�8g��U�(����/��}dg��"�����_jw�Xv�13�8 ��!L���T���q���A�᩿�*��ʛ&f��G���y��u�1	]�+�t��[Z���A��u�f�WGQL�Px0x�io�mF�n���)�j���;�@�ꕐΟή��,'�ǽ��t�l���w�k��w��F��ɯ��l3�C�⎱�ϑ
u�f3m�ڎ��$KPB��_�H�?~�v3RӲO��pp���Y���M�`���{/ե~)'��~�O��,d��*�9�����v 0�ŔM���*���c@`��,� ���B��L�=�HJ�j�2�5�!��dYN���[2�]��1���4�s�ZǗ�&፻h��2�E��� B���$�J�V �8r���$����5������ `8i_���u��7@-��s���T�7#�f�;�P�������3�/%�����-}nS��]�%��!����d�k��w�2s������8�>�w�t����E�Y�����QoKG��!�	8L7�`|XT%#,8i�pZ���W/kmu�+pr.�]��Wi�:�j����oJr	o�Jf�h�݊��a�n<����A�Nӿ�EA1H�_��fč5U-Y`�˞���������9����� ��wEMd��[d�zt2��{(��@��qAq|�J�H����ь�V���`c�_���r���Ǽ
�X��E�?��B�V�C3�p.v�j�kVB���'d��|��I���Um�t�=#0�ץhM���O��II5�{�TQ�L��؏v�<��=�;���Ǫ/�y�u����_��\$<�Hڦ�N���J��ȇD�' ��X���Ϣd<)�Ƀ����U�%ުj2߹���q$8�h�O����Vű� _�p	~�0T�s�?p� ��!b�c� 5�mR `PzP��f�/�y����K���`���S��	�]�O[cB��m��M-b�Ş��kI�����1r�|+�ћ�Nl���W`��o�쫁�z &JQ�k�t�a��k�$7�
�;Dp��7��)�l��s�d�N�������	`9��(�)��gLK�I�u�ߚ�uN�n��X��5S'˟�]����`QI�֘%<��D�"j&�+4��U��.�#%��47A��N��N	�X��`�!E'N7h:m� '���;���x_�;�Q�}�^j�d�,�x���������?�O��V����B�p�b=���~��|Q�`O_��y�ᖑA��}��;� *?G�l�8���?��T|�R�:�LM�/�ņd����CO6�m�R`�\�����]$�gx��a�p��ح�8�y�!l���e�F��(-@:��Gl�`�hQ���Z��	�q��<�:M@,U�{]���i�H�n2�3��tBu,\��E�
����P���ެ>r�+�޽e�m�������4��2a�hB׻]"�����E��"�����X���}P��*.;�PW𴃣�ŐM ���������J�2{�9�chg�@&+��h�j]��ۋDy�@ji��H�k�Q���w5wm���	<!����P`�,������<,�SE�ނ'��Ď9Ąy>��^�Ww�>��pnFiON����_#�|'S��%���A�bu'�O�ۘ$%S?�~�N���,s��l�I i�@�j	��r��π/�#'�c��v��������C$ �ئ(z��@=?��Q��meaug�KqńqtC�*�O��=��/��Z�~���ߠpv_	{�ɚ�u/M�uz��P|�o��~�\�:j��
��1j�(u��< ���B%_�|0M� ��qaV������w�=��c؅�}��,ٍ	�=#A�n��='wh�F�Lٵ!�-�xK��j��� .�ܚ&�F9��)p)�q��c䖿38�U�k�h�n�kt���-(qA3e��oS9�,�gG�W���[6��?���S.�b�G�"*U	O��zt;��j��7�!Z�M��¢�Z�~Z�3\�&����M��1~l���ґL�P����5��.!m�0�ꔧ�s�ik�U!���<U;���ӵ�=��u�R6��̹��½g�$�bjF"�`N�-�m���!�7AŘF$�6,�����N�x,��tb�K��O��2����{�Y jͿ��;���-7&Ӑ��l"h7�y�9T�F�dcٵP��3.3�QR�ƌ�Xj�AG�1J��r2 T�R�ռ�q��`�����q�K�] ��,w.I�1��R;y)�obr
B}St�i���7H ��D��R���Y5o�/�}�އ�yBk�׌�j0k���`죀m��@)�Ӕ�a�0cV���㌢J���x��E]�!��z���tZv+����my�}+��`�5��X
�\�f:^jB[��'.xP�J��� ��#��a�$��zl�N�įT��[)�mt���K�I�Z�?��G�f,��gRI�%��,����:�'pt�C��,!%J�-�7��L�����p�;�~�KC��|j/��ErW�h������9�'�k��GU�a��1�1�.�������u��zج4P
I���R;`���lM��M�z��4f����T��0�T�c՗�����7�g�an��A�����į_��R�㴯���70o8�%��F� ǎ�M\u��Y�8�RjV��o��FU���:
}��ƋىL�2�H��tU�]2�k�;v9�Lܥ ��y�X���0.BU��&�ဒ��),J-��Ou~g~�����������L�t,Pq5��M͞��?�����8�ԃB�V+H��Ԁ�G��:�37�_��\�Q(�C٣���Xv��V������<773��e]q��ﱖ�t#��x{M�5�|n�1���'K[���a���\�� ���,����r��ûlז�;�W��~���V�2[o'v��Xǣ��2d��c���� '*���9'�����E���T�2��×��*��5�F�'+z��4gB�f�H�G��p-���G��3#Q�T�D\N�J?���-��73{z�~���#?�iJ�"-�e�[LtpD�𦈨�J���O5|kJӃn�*QV0z�qA�M��e�v�o�*3����S�"�.0�2��
���t�F��)�O�^;��)�:����w�vs~�Y����4#qe�L�����]3��2�HU=J��Ä��4������*n1</��9�$��/V�Yi��:*�:�HeG�+C�eL������EE����W�wR���u�e�l�TB�=m���@$�	Tm-@TOg��n���
��h��|	�Uɺ7�AUd���<|=��Y�P�f@!,�������R�6�c�v��ٛ��w�U=��k�;�?��qͬh����(��H�,�6Mצ�U�y�C!�[h��mO�t���&b/>����I��Ɵ4?��D$�	������>7 �A)�6˒�s[���`t�5�b�\-��+�E��xD���|#vH�	waF-۵�yY�nI�^�rɚ<\�狽�;�g
K,��7���&s3�{�R2.�i���{!*4����itG+Hl]�ɕC�k! 
�ݱ# ��̸SrB&ْ��+N7'g����_��@�,��+r�,���.�zpb�,��D%r����/�����iO�8�W�>̎yX?�<�n�A����0@�!ڐ ��L��&�\����C�+���ݢn�W��D6Y�"���RLAy�����[N~б3fo�{.�
b<�Ȅ�1LOR�qx���0x�4�I�:<�yGHa���"h,w~���R�.ŦΊ��&3�+M�I�^pXt�,>�� ��VY�q���h�'��zu��.î��k4Â@_������ D�OXn�X�9��!J����Wy��K5#4֯�lPG9�,�����4��W�D�1
��[V���j9ydaVHF�} i�����Ysx�E�'(����:H�X-����\c��j��
��~BPX�g|7X�~���Tݔ:�H;{ۏ�( q۶4&z����"��Gi}uYG�W���fZ��t�`��2:���[�&�>�R�Iͼ>��iߡt�aCXޱ��Y
Fܕ-<�3�7�,��W�2ݤx"�$�6�]O1E����W�0L��S�Z	����q��/Ų��.������Ů�JX^�!�T���&����u_�_���B��+�GPbYn��A�r����G�(��