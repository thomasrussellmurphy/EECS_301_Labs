��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_����m�e"kxu�Uٲ"#oB2�-g�j��h�p� M T�(�P�+M��&�[���+"�:%V_��	�Ξ�܉�����_̯��֛%�����A�Y��Y]b������ju��e�c"VoH��7��ۆ9O�5�ҋهO;�������w}7:��yFP~�%ti�_����q`�$H�,,��Y���^�h����?U�=��56VG{-�O��D��y
a�=���B2�w�@�Ad\՝al�O�P{��|���//.qtq�cI���{���q}��՜�A�)r{s��!9���2=��pSO&.V=�f��R��_�(^,Ak�MF t;-�ó��]�s��s�8I5�L��1
W͋P���m|ߝ�@0Nu��ӎ�CJ���L�v�9���>x4/=�7/�TZ��5���ra�q���1P��%׶Gmz�'����k��&����ȏ���ޏ㐉�#%ea�u��m(	B~�1�o�ku����#��z��L����_���aT�b��g��"�#$���j$C������$��r��ը��X�K�q��8}1�銘���q�i�z�����-jk߇�0k�$W�]Q���K"7/�V�ώ�׳�VT��\P�����v�����Z�N��$�Oyyt�*B��W����#*v@5�ƙ����s��v[⿽K��^c�8�}d�l��55xҍn����X��PW��m��[�ǵ�t�ҥ�]�(�e�A����K���Hg��B���9Yd�AD�`��5���z�+�E�ښ8�����.�������>����$��Jg:%����6��X���,p�E��sZf�965l�]f9A`\�����3��{%<6��Ʒ.�G�o��"��H�>, �L�-=�EW4� <2E��� l�{�γʿ���Aݧ�e��%��EC��,����]v��`ٟׅ�T��^���4W̷�<[�`Th�����1���8�a~�����
�/R�<O�r����J���e����C�V�/m��E5�<�i
�Zf."�T����}�|M)���hB�L�Ho&�>Al]��l����/�*{$X�b7���[�p�h��0��.�6%��l���H��$�U��z�W�ީ��ǭ�,QlXP���!fo���-p� |N��\kh�#�_�L����;�9�6䋑�с}�BdcA�D��E~�#s4߹�I��L�8�K�>�_� �YJMe�ֹ!"�̡W���u2Oΰ�]~�'�5�sݻd�7�7�P9�p~�����[f��q��#J�:�=��
\��K���gA��/>�T�s�ŭ�4G�'�D���c#��#e&�L��ҷ<T=~���,Md��nCѯ|�XD{�=�����v��C�RǑ#Ma�,95,�-�wLLg0�mF_~��%)ϝU^�u�ɵ��6��D��Wc)�@��:��9�i, ��F��L[C5���@Aޖpq-ዘט�� �.��a �I�{orƬ��7mi�rG�$����k���|-��K}h���{��`l� 
Tl�� s5�0��g��I�����ƥ��ab�47����^)]JC��D�Bv(��� �]v�B��v76�/X�ϙ/�B���Q���`/$�S�Ϫ���� �q�5N��%�����p�,H۹�H뺊�,2�CtM�Q���b+��'O|{=(��T��XPՍו�S�-J./�]Nb��A�'"k�@ ��]��:�Ȋ�'�\�H���P���lM���Y.ܦ|b�#���zg%N� �!۹�e�rB�=ʌ�@ߞ���r6gw�L� �^�e;�w@�R�ν33����ϽZ +#b6�`���}�����}v���J��?bv��j���zɷ�e���g|:`�����$�"������5�(2����?M�&�r+;s�?�<Q27�s=nF�����F5
p����o��������g�l�2���v�����)o�g�=��"N�>��������g;n+]p�g�1� ħ�-_�=q����SXb�2���M��ݟTr���!����,x��VQъ^>|�j'�4��qY|H�~a�F� �Y=�2{�;�&�G�D=����&�&j����m{q�bً&<�w�.�����Q�U��Q	�i�� b���d��¥�4҇. 4p�e�0V7H��!P��"4X��i��%�$�AS��sG|�	�|����j��O��5+�+���̮��M�0l�Lh�H=�"���M.߶��_0����1� ��x���X�}�XqBxB��>RU���	C����*ՃGv�s��W!��O��~�I�s{��s�N�D�Г�4y�أ!�p��o���.�M"z^��/�
/��������L�nj��B���v�Z�A?w\y2���<wF9
Ux�h�X5���=o�j{�bO��Hd�B�M�Oڳ�UV/3� XU�"��k8F\Z]r~P��9'.0��25���`��0&�ȧbϪ�n�� �TI���:n}��><��%|r���j�k^ݼ�@{,�0s�5�0S���~�\���"��l @��m^
|�7h�S/���w�_��RUt�h�A�z�.T�kO��}��ςŤvx,dN��7�4n��A��(�$J׃�d����+�csn��u����b�=�gI9߃ӭ����U�����7ǝ�dq�֏������3ze��H�։���P?�(�����ϒia��kZ4����Xol�#�a�&�!w|V�����|`/D�g-_	��eĭy��t��lBYD�bW �E����� ���;�YKv�����a��N