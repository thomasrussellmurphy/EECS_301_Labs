��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|����z=+���v����Tn{������&��o���R_6��F!k��j{.H��y$�n`�)n�Y�Gbbd���-�*��������͝�8Q:|[��@����K�L]��W�*+#��l4|���~3�r\��kB�s"�(Ӏ(}@�Q�~ZJ~�*d���@:��[6��V�!g1���F?���Tcf&OH�g�9��
�I��.,�R$LC�ng�ǉ;i�a}��V�G�첿B�����~��xsz��(�R6j��wk&P'A;It���/DK�h��߼��6�9�kS���*��\��e��u ������'#hl딀�Tj�������N[Pvn�������X�|rꝢsW���n���n��l$��l���б�ݻLтRe�Fn=���"��T�{���F~���	?�G��_s���$�[�"²:L�	p1r�nj�6��!����P�|�.�F�2��{�����T:_%@���Z���*��׋�2����6��k�:�ٺJ��"J&IQ&��"�C���u�H�b�ɴZV��*�褀�6��([�;I=L���]�?�A�ś���lm��7�w�#�����%��J��J|�ԁnw�00E���aO2��@ėU[!�T���̊�U`���zy ؈,	���s�r�����_����^��kq����4c<�G�!9Ɛ��\(�BP���$�h@.���>��:w|�����I7aІ'�.�
�������t�%s����*�C|X����U�hç;��|
L�`�*r�=�K����eG���DZ "��E�I�{%��jg�˫ZG���>�zo��A]��R.��@S⹝�z�*uKx����W� ��$D>�2�أ:���|�;����l�
o��\�����-�'%&��������K}�5��~v��Ո�H7����y��9��c�\R�r�ܔ��!I5���/�z���2C�7�;u�/���b�*@�T��m���-�J��A�/V�`��*vr�|�Tz� *�4lЀ"�������p�Ph�[O�r̪�v��nE.��@�Al3���^X���Y����LaE���ض|�F�*��Y�&�I[�x��&��1�V`��U�=BT0h .^k4��xz<U�{ɈV��{b��M�f�d1xv���*���Cpk=F�U�$L;,a#?C��d~r��I|�u�]X�FbT�)�c57~>���yz{�m���dh.8���q�4����>ol�E:�8�������I*�{M7����]=�ܘT3]���H�2���3S�~7CC�m�m�bӡ?d=^�Tk���(h%�y�붵7~\���88sW:���=����
�Ҡ)���
6��M�`�p���F��T�m{d�u��4�`�#�C��~�5�M|�G�+/�
$�6�昗��S���v7UV�<��W�c���ߔ�wj 0�ߏ��=�*�Z����8�7��M�$�x���°'R���ͷ<��GO!R %]�
���7������Yr���/�2�3�P�Hf�g�8����oq4Z�$yQ)��}�ES���H'��ف�r$�^$������a0=Zm ~�G��Ji��8JQ0P����
��s�Kn/+m�vG���B��#*�הoNK%����~.T�x5~�%5�ux0k�VW��A��2C���\�̵�wSng��k2>�,g�o���MJF��Šw��u����2���|Q�(]�{ �)9���C���!�0A�,M	�0H���ɹD�H�0�m�����_X��f����z�o͖��~a�B@#x�Qt9/zIn�	^�Ӗ�
�-�Xu	J;��-���89<q;�
��鵮T�L��2b�$NEwV͹	�a4��<�*�k4-�(Zhс� �JZ�V�gȴwl��b�����k���H❍�k!�H1�R�4-�Ix�Y>�gOע�n�\%����fv�#(oI\Gc��$sR�*��ʌ�_,��g#$!gl�z�
y�@F�Wab�0�Y����?���Y �C�:�BPm؉�Q�5n��bc��U�����k7��X	x�q|���C?���]}w��:WA�w�x�D�̏R�u����˯�y������*�7醧��ѽ��!��M6
��P�m(�$�|�ŭ�zA:�N�nr�Y��X0a��/5�A��TO@��dC��e|�����B�Uk�&�>v���0)eh݊}�v�ͱh�G��L�N���kH^@��:j�q�#"*�R�50���;�y���g\�\èz���Z����,H+�L�yf����¢ʎe�՛Z��F���XFn����riT!1"�Z�TM�!����M
��P^Av��ҍ��D���d��]�wu=_���O��"���*>i��a(�y�ɐJ��;ü�i�Jy���/m=-`�XaB�ʀ�ǖ��}��o�q2��#[��=�$�����Zd�J2'-^�j\�"�d��*�2/V��m�z~լ���0\&�Ҏ�o���[J�R�T�(�?[S��{?MH_��r�D�cv�Yj�3x�D�Fr;���EQ�+:��A��Y�9R�sۣQez�?�����H܉�[��΍�N���@jA�%6Q{�ۆJFw� ?=o�`�;���5�����y����*#2
�O	 ��m�ՉI&��=xt��z��	q��
��L1�x(�&i�:�9�=���9c�/��l��U�Z�@CM)���S=��-�A���&�L|�d�ڃ��N,5d`����{���RÉ�,�% �ܳ"=ςif����3Y�]Ȉ�]�<��{�<b/��c�ˍA�6�Ǩ��_�� [�q� H3�����Q��N.��)	�0S���I���`��Ae��x��ҩޕ4�]&dK.!�v�aE�;K�n&�=$i$(�r}?��(ѱ�6����".�MS�*l%Kt~� ��0[O?����0̒�3��sɨ5��D�� �CX?g!�GZ_��v��#1�eV�l7�v�$�2�
g�&�
a�ڒ$e��-Ư�q�H���7rq���UX��b���Ek��Nl�U�b�--7���n�j�(V�g:N5��Rz7�/0y�&�̞=ˠ0�D�-6̥����q���p���7�oN@TaȋvZR|��/��>_��XZ�P�5��{��J��߇A��	=x�qn0<��F	}6���/f�r�GyO�}of���ܤ��3��� 0S�{�~W��Q|0�w|Hܭ|G�V��D')-���5��䷾e~��`3�"�1��3�o��:��|�-�끔ٺ!��(CT�O����s܃�@�������y�b�T
hNQ1�3�ˤƩ}�=����mwŵzHq O8��`���6	w�H��V�)$�c�*��f�pE�u� 4�e��_��l�&a�?*���"Aj�g�Ȃ{栫���	k�*�@�@�_�1��9,�=���Ky��3��o��E���D�a��;W��Y
��Ri�e��<��b$�{�ӕ(�2F����E\P-���m��Î8�zB؄,�An������ճ����;e�P �f@ψk� �����"��/��p��x��-�e���Ѥf�!���