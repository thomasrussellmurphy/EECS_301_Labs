��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\���V�fnvx��ÍG_;�ȅe�~�>���9�>��Y;�0Ga�%m郵��DTZ�!��}TU�M�4V�f{��A����m�dڔ��ċR����Ďa���"����/ �V��Y7��k���=&-�k���H��5�;�3��������ԇ}�$���MG L�<)8��b��SR7Z���fG��ER`�rE���D�ORl�%Ġ��P�˕���n7��%�i1�`�[21Me��Ҭ9	[='���\��-��p���U�r4d�{������d��H�	M�����S�k��i;��W�/�-skcFbLv�k��N@�8����eޫ*X���L�^�o$���$ �N�#��-j.f6�+_�^��4G�2�� ��P��7n�]��=`������U�[Cd���o�}�֝K��`x����߷��%�dz���(^hpf2�v�OWI���}]��,�4�-�cb�TE��,��G)ޡ�$��[1�miK;wW�"��x�e��sˎIY��m�&��y#6",���*�<�9D����Z��.�#X���\��Ȟ��VoD��{�Q���<o�?ZD�D�	�ҹ+���������S��XFuZ;���0������.���E0
\`�X�ε耨9�Ê�9��i���ŕ�v3R+2�,��	�R�ʲ�A�j����5��q�x(��9TD<f[d�*	��ā�$_|s�he��	ғ懬�֗���i\,��:��w���p�E��;�1���F����Ͻ��
�/A����rYZ6��2�T�߭喝��a���-z�1T�$sY/����R6IۤG�6���(�y��q�q�P��{���(O9���@[JA��W����2.(� ߣ��'I��Ĥ��Oh��+��|�2��K�2fSC�!8)��X�+h�<���cmWZ��j0��é�(�m�	[s���	ܐ;2�)8�tD3\ZaD��99諨,*��cq
�2tƥ��Utt8�W�3'��v�K���̣��XZpM���NQ+ݎF��J'�c���Z�`����oI�6i|(=5%��=�������-!vP�ĭG}� 6��_&B�����*O���\<��iA4^��jk��1N���tF�+`�4	�˂r��O����d��4�&'�����)��Vr+���$�*=MaQ?X�Gi����d���'��b��q���	xI/�ߓU�y�����8�u�E��BpZ��燬�R���ͬ$�5AO��a��O���ik�"�ٚ�#��>"7�y��U�B�r$-�����B��7����W�3�K]�ى�[����!oN'ΐxF.x�5B���^�v�@_����N��`o ��iz�^���=?���d1d7�=�����lM� ,j���-.�������J�y;�ϰ���|���M��@$��Tt�h)`8��
_��e4Qa�	��V�G�Z�p�l��fV,�ޜ�މ}��z��׼�V��}�6 �^�W�Y썫S�)�4��4��o��+��a.��!>=�o�i��R%'�CĒ�x�T"A�AT���T�uց���L4�Jʥ�����h:%)�M���� ë*W���FS�̓{���?�~��Fe�F�Kw�=<t"� L�`�H�6О�#y�H|c�Ǳ["�������0�O~n�j�$�p&�ﺬSL
�ӣ�Zp�iT!-�H~Q���&�;c������-8��P�ⰵ: �m���͝��w!��m��Q��ch�y��oR��)FĦ���p�ޮ�!*�et�`;/��<Y�}�򉁏�����V��!B��������߱���(?���Jdџ��v@�K JD>���]��yf]H�z�  p�;�t���F!��O�'�V�!8��q��f8_�:1�W�����Y����e�%�O<��4�6��;$eD >s���g��0X�c���5e�S����5R�� �t@��hmT���q"Y�+O�,�qFZol����{�Wq��[���.S��q=���fhk�;��/����ب�������jщL�;�uHO�W�����k��=�eDd�<�pкA2�d3�����tȁ��=M�fZ���om).�Q&�T��
�)��[$�㛻)��`�Jn?p��۟Y�O�IvBlqg,�.B*������x2���ww�;i^^Rd�3�?I`�E��w�y��{Y�6����o��B݇��v�	1�%A$M/�K]�P��켶�|�.�w�n�#p�ĭ�����O�[g9��|�S �ڛC�8���hy��R)�=�Ԅ��b�����O�G��_ge��AtF�Ŏ��΀����PZ#�����䞋�w�(��������6��:�"���Z�m�������:�*J?���MƷ�Y���:�$9�[���R�u��9R�ǳoD���1�-q>���(P�镸q�,O�x��'{��gz��E����@�x����Z�x:_�]@��3px����(�Q�咎�m��/�'�2
�?�@�H|�24��$����S����� 'l�|?:���^�I�W
�k{����u���plH���p;�A��N�����ݙ�,�����{�< ��Q��Ȝ:l������ɉG��a���3�W��S�8�:�
�R����{a���s��=U�~�[��¤e���F��5��a���W��1�h���
��P�p4��Z6�P#�P���j���!���	�{�s�W�+�#�O��H��@H�\��]��8��є��p�ōv�sP֤"˘.X�fQ2��Cؐ�_��)����(x*%��X��Ԑ��.�W���Ҷ/�Lo�`�Q~H�+�T�cgk��O�0�m�Ju��1���|�����J�\0����Ryo��\���e��H��B���;j0/g����ʃ�nD
y�}��K|��e0vaO&��WA��s��}��W�T\���n�w�0�c�>�*^�iHɳ  �G@�H��t�1��&�p�R^z&Z��D
<^n��w���_�p��������*�X�L~y*����δG�^�N �'��\��M� �+ۍ�C)pfQOZ�	���U���!U#yP��E������{i7�F�ʳa��^�ʱ�D�_����d�lKH�c�Z���ῥ)�O�^ރ�Ĕ1v��ؒ�y��!� �g�q�`��w���_4f2=xk�#�m8��!�+����T��}����k�Sҝ�2!�nAҷ�Y��0���0��;���"k��Oq1�����a�����5:m��	�vB��ע�b�ɿ,�q4�DS����xX�7�V-{�ǎ�x^{��W3�ΎY�7���+HOCaO@�.K ���+���^�E�]�Y�y������$�-[�	g,[@6�R�uv���4ƓW�?qL/K��,4���qٕ^�3ΈsV�� >*���~%o y��׈��|�d|�C�,Xl(�%G�<_�J��Y�'�=��[���''3i+&_�LbX�^���F��O�YZ�#���"���۱%1��'��/_�R��T<��8!|��a4�+@�|̓\�3�m)�c����J�8S�fA�<�O��H�E���Ň�Q�흅�^wX�w���ǪR���G�[��!΁S�'�x�Au{�z�Dd�]*_2���!ܔ ��HN�-���0�[-�N��h�8�d�;���:��������˺.i[�Y�k�
�Θ˷�7��0g�C�DqMG���=F�1�
�ƒ)����/�/H� i�6H���#as
��	ۂVs�p;w�8Ŧ�6�/����^E�G��]7vw��{&�ưj/�7�:�Z'79>B�@�U��#g:w7��6g/p���@Y4B�{7�#�Ήm^��E�Cb��x�v����T�fl����ޯn���u� �V��X����\c[�U%:�����R��2���4��}�x:B,�����t����J��}gߨ(N�I6+�8F���w>O&�ڀt+�#��<�QТ��|X�i��0��L�lZW����4��`�<���I�[?4Y|oT�t�K��e�怱D�u`*"u�����/=�<`�v��a����B8\9Ϥ�`Ȓ>�R�Ѿ�����(1����1=�� �mDaNѾͪ� 
Y���Hv��[������K�+U��]q��G%_ux�::��U[�Gus�d`EL��fpP��N�S{�7"i��k憐$��ii�Kv���$[9�q.Z�����/�E� MK�uV���5�(��؎ث�f���j��Ɓ�|/�*fvi�5o{��$���Sl�*M�X��ҟ����PG���k���R��v�l�O���D��VU$`�4k��"e�o,�X�_�;��U��K����q����?t���.��F�&9��{ �l���S65Xu��>/ړ�Q��<��@���r�:�����1[y�K�t|�c�@,��~j�K �}ߕz������LN���Fz�����έ�*�d;��~c�*��=b�����m���j�|�L�K��p3Z�'^�^
QD�s��)�U���6z�Σ����;��>9ͤd0HR��*�@G���?��`�U&4��II�PS�G�gQ��غ�<�B���<q���"��ԉ��%���K�*�7�˸�6&w�%Fޓܾ�,Vp87��&yb�bp���3�Y��k��]�|�@���s���X�a�Q>�27�H�kZ��yb�a{�)<�g�>�A��hC*���8��U�S���T�i0�zj�8ű��D
؍�'(e�%W7��VuēU��yVI�f������*\L�H	�(�s����_����i߉l�8͹u����s$��c75
��1p#BR���ɱ{|���f�!*�`��A5Vgd��KH���S�� X�^̩�I�5��#��#"�f��(�7�ͨ�N��8�x�zc�Hq�@��k%�ނ�@��cR��d��/�5dnկ�5� ��5��U��	��ϗóD������r�s�q�t�u�Ku"|���[*>��uP��)��زc��Ќ:�)��0	b��5�/�9>�~ �.��X��{$?���;��?!�AgН���Y�Y���i�y@��������ʆ{���;�ֶ���ΰ�Tlk��Q�e$���P�n��m�{c���J20�������=��}��5�{�Zՠ��6Tܰ*���N�B;EY!Y���&�z)ػݗ��~P�[p��7���w`;)��Nu�Ba�z;nFg�|(�}��O�p��2�<������GB
�W���ol�/8a]D,�* Cu.��R�/��(�����Ò��3���o8����x�$N�����c����j����5Ff����F7�F����e��e��������+0�# mT�)��u���'� ���~"9��0\���w���4��dGA�N��J���S�F�0�_	��"��T���w��>��/q>h����%U�ƍ$�Ӎ4�Ϫ�0��Q���6�X$&��/���Y�\�[�9�&���x�)DdNG������lcM9��n �$B�SY��?�Ov��#rs�Q�������ԝ�Y����aR�;�H4�(E!^��d= |�5��<��v���x��P;�}����C\
qٲ���ȧ��ƙ-j;�rom~w��{��_��?���L����i��biF�e����.�������M0�����1��5�g���.�c)2�n7N(W��PoM��,~+����4_ɸIlO�x�_�EA�I*� �d#���$لO��9+��?�0��'�򼦾�z@y9��Դe$Rxa�����J+k՛}�ri�$j���{��Εk f7s?_��l8m­�E�Ǽ�L���f?`#�\ )��J.�5+�d����ܞ� b,N��yf�]8Eu.�kQ��)�wn�4S���_v����;�B�嗜)�����d�A����Z3���U uR%n�V�wJ
m1,�x��5�{#f�	�8�_��>OLm�<wS��X�ak���MV�8�.��n,�� e�j������]W Fu	�� ��* �-�!e�0�
�h_�0-�щn#Ȁp/M�	�I�@Os��R�1n&�8��5H�ҡ�#A�5�2����e�L�8>�4�n�=�S���/�__�.+v����3_��+��\ӽ����Q�/��}�ֺT����1H�E��+�8UA�;Y-a��ǃƶ�]V��7�����s f��ϒs*'�#�}dV�YÑ��&;���Q0h�?�f�D
����������w�"�!�*oT�_[���j�兔8$��J����H����=�?���Č�F�P������mQ
+�Om��l����H��2���u�=]�=ke��3:C��rs('Te�r�(���(��Y"R�尚'�*����{|��Z������������Ta������X�@��I��уS�nE��h�#�+������!e~,O$��a�,����1�2E&���`Xݔ���
'9N��h.��L����R�Z�0�+70���U!W�I|�����,u��`k|Q �h&�[��1l��rE�8���U��ۍQH
+�݀�dA�β=T�&	X�!�5U	N��N���K}�֗"1� Oΐ��S��'��}*�x:hJlG��8�'�+_��n�G���:�߶���
����7m�4#g�{H��%)�1�_e1��QG��L�5�n�ou@��_�.̼����ϓS����h�$��b
�K�4��?	[ya1(�����f7 �W��"��S�{B*MٹR�	�W(����_�s�K@xx�W�2��7y�*$��� {^���xY.�J�p�1�#�F����8��j$�P���P�	����o�k}��:$uYg1�~�������2��qE��*�L+��NR�c��go; �N�@��kd��"��^p^�a�v|h}��$1Bn���L\�D�7��KUp��O��Ѝ��������4d����A�� ����
q��/�(
�O�5�9��ꍁ?`�v�!�/���|w�O<E<�����.�D�U'O9�B�c�]8���7���Eރ�N�(��}B�s�}��W����,Q������eӷ��F�zV1Y7�~��������R��ih[l
�{�@�O/b����H�y֎LyhxFk�1�w���'34R�EV`6T����)"KvIڐ�9m�{�A�͉*�
+��j��(���-,���\��
�֣t�HcJD��25��i1�##ì��#r#ܔ+��"�y�{�K�7��s�9���nT�ޙ��X��˴�g�qE�i\�̏$�g8+/��
���B~�������cj���K����V��'j��]�~	��P�tJMNj����k�z�o3+�,81�O�����@n��:������rI͚�D~���_.�."ep�<Q���փj�]`��"c;Y�`�c�Nf��w\<,�r7�i���)�g/@��-@s�Pd,��}9Z�B]�6{&���_۰j�[!��w<J��`L�����eP�5�TU� R����d�}`��`� �Gj��v�v�C`�wvKޡF	����7d��B���"`Ilx�HQ&fS��'�6xF��ٙ@M�-˰/e�QK�[�!��އm���%��(�e�R�T�P��$bm�m��>N��l�5}3��1a�T,>�_ G���[ʙ��C�4�gS�G��r�Ĝ��F��B�-�fH$��>��q��\����K��ߢ�k�q)�-)�̩�?��?%>����-?��!��H�fa�I|tp���/��P���{��̕ ^��.`u��fV��%��Ť��/t5;�\���G��72���r��-�yh����	����\�,�����æV�+V��i���q$�0�|��5�c���Un��`h���bleDk�=�Z���V��3QΜ�S&�l�q 	���.V���5�W��T���+&1��[�˱Y�3�w��

b!����#a����!&��3֥�v�\��G�q&����U�>���w�|��+���U���~ƞ�  �q�n�^A��rw��#�U����y����S�F��]Z!e+���������A�ͲG]�d��'�tPY���$'��T���(�4���'z�I2q��{%�2���ii��+�D�E�F�f�}_g�!'���p�*3��h^��YS�p[~{��ҏ��������<d�h�>T�B�)m����W
CZ0CSJq�QE9��Ր�ɫ�a�S�VA�v��0����i�Z<��3d����@����{t�2�����&�fЬn����ǥ���jQ�<�#lkƈ}��0�uNj���QK>�nU.��)5=1���xI6������^�������#���{U���&�o4%��Ua1����,��ؤ�-�,�B�J�u��:E'������W�mDɘ�ش�A���X'�?h�i &5����B^5�U����ԟ�ONA�0ʏ��t�cp�#��s� I�PfD�i�+X`�S*�PwL����c ��GY��3���Ln:�?CvF���צ��Q��DΧ!|������*����dxX����o��k2X��Θ��{�^��c�L�\W��:�Ru�������Eo$�	G�~K% ��Փ�[��g���;/:Ӟ����T�u�ꆐ�'N�\��n��w3E"�M�6�s�b|˗:�79������<��ۍW��u�5����"�a�S�Xe�W��G�3��m�Y�o!���.h(UY��{�T��K��Õ-q�7�N`���7�Z����cSEq�9zAfzr���)�\��%�5���P�a���4�˥s^���H��t1��{�UV��oy���;��[�G�{T^���e-;�d��a��p��,l���Hc�{%2{�c9G�
X�􊥄g�)C@.v§=�lDG0(�'����}1A��.�30�H�6��$�I��V	ܧ����<���e��l2��S�����z^�hj�x͝N�<�:1�1�6���L�YB0���������2n�i�M��m������3^�J;�Xqؿ��������-]r�LRoz1��j�#��-�]��_|!T�`��ѷ_��T7�~�w@�'a�Z4��~�m�S�}����eT7�3�,ؗs�R�>�����vI���9U}6��F���:1��޻�$�Ȍ�����-�S����z�dˈ�k������=�<�3v�F�i��(D�`���kh;d��|.}]�t���3���Yh9��7�A7����I��a�t!L$�pBĵ

W��÷���D%�JBy~�&�e��&�x9l��p���n�L�TP�X�U5!a�9�c�U��ib�S��hw
��3$�Ԑ�%S��=���Ո�m3.5��0����ܵ�*Kd���֏Bۅ��mka>M@�#��qþ�`����-n�p�\���LZ!��1<�O\��8C���j�]�]���5��h�Ž{D�6�����uz�״�[b����ySJA��)Y��,�R �����B��d�v��?�9��}���� &k4��!1Z��������x3�ځj,�%��t}TJj)1GZ�y�+!���G�N�w!�߹5�H���O�eC��d>��(������f�o�]���6Q��%d,!���;�&{P)�y�pV�&R2g
��{�۠T�HE���dw\ �:	��
y�?��i�.� �(ݩ
���Oh"�)qvW�_�mQ~E�Z�����D�Y��B&��ajy�Ѣ�S�~��7mmj����(�������n~��k�ŁKc`�la���2���
И`շ��UPg��V�p�g��Veg �*�@n��N>  j�ޙ��B�*�Qb�W�������z!�!Nda�G�TF��M�Կ��� 8)�r�ޏ�]��F�����p�?�����N>�B �<���y�Ùa�k��6�-���OLrr�a��$	���o.���r�ڼq�^��Х�5�A�ח���$�����-�����.%����J�i(��Ǿ�u��&kw�BH����Bq��^)簐����>����ߎ'h�����c�N���",��x�7�?=�Y��B�V��A��y(؞ #"�|�����������.`�	1�ק��_Z�Z'6i��A���&V2�� ���sb���I�e-s�Y���ǅ}nXv�V�сHj�g&.w�*��6�MR�L��Q�d3��E|j@�Pz��=��"(DS8��l�檝\�,|�!_��#�3�D{��ގ�/���U&��qS�}[}���2�)�Y��!��*v�3��Q�#v��֗��*�-�=ww�I(��ޘi�Ӳ����/<�����]+��̉�#�O�wT�r:�x�Ȃ�v�|�\q�h��H�Nix�T�ƙ��G{�yN,1�7��������NC�O2��H��B���Y�K���(M&�N3�8*�癏�ŎH��p2���L�L�4b��\Z��Kzw����E���>cX�]'"Y5���?uA�"�u�X�B�>�Ҷ�D0(c������]0��u1�T4N:-��8Zd�|����BV����ަ �.~�w_v֡��u�]�ϓߊ�����,��{�wsoU���'1P*�w��k9�鴫.-SW� ��&�i�
��[��?�`Qh\-x����1u��V�tړ�����������Ŵ�8;f*:ߤAo;�xm��'�z�i�P�1
Bb��N�/$	��bj*X/t���d~��3Q$�9�<��&�cR�4�����>�4R6I!�]�8k�.��8Mo�)V)K�f0��#�J*^>}Cs[i�b��y����B��Z�/���A �	��F=F
��)q�H(�&�k5�_.zrT�׏��轾�\���h��z���O]yt�/K�;Q���EJ1.�!-�	톟&�\iG��'#3kx�7��Ãz#L��~z��{� ����������g|s4�;�z�@����v�?Py��c��g9(r�O:wE���	kL~*a![2Z6�B��d֝�bL>���VW����us2�Qɻ����߱
���v�΂���;�Ұ�~�K����i��vɍuw5���������V�)g��^'��|��]꿝S��v��o�7�]��uj�8i�1US rq��{ ��\��
��,�5t8�u?wFx|�g�D�<ę�s����Ɏ�6~7�1����8gh���WP�*s�ٷ��M�.	�k�Mc�*�ִA�<w-ҳ���[cb�q�GN�w��*r�R���CH�<���~�t0�O��!Y�S��JWх��E�AQu�c/6�J�ŏ�W�
:3F��5p�+vG��U�Y@��ξ(�?�
n���`s��NR� (�E�W~��a �\0��+�]�׍���Fa�:�z��� i��9�4,=]�7dm^�ɭ�M���X��� �@��	��s[9x����v[f@�τ/_�g�
���=:�m��B�d�?*��\K��#)���j��'p�fX� ��!Ul��5�,�V!��h��U>�����0�u�?�����|��FI��S�'wQ�����"���t:�h����s � �K��^\mӶ[k"ʷ�m@��I1�	��:wj_�#�M)��	&�dF�Ym����Pv���� G��`#�N���C�}îNu�%����0�ޣv�N�@�K��a�����v���T!x��ܹD����oJ0�WWMK@bX={d�y��F�g�\��z�=�%��HZe���|*�3�1w������r���C�W��~�eŠ�$����܁ճ�{�֣}u��[\��'V�x����z�S��	�c��h+���̺Z�ص�3PeS�nIm>����0&�C��S"]
N���SJuxʹ��	9�w�K�K}���w�w�Mq-/i/��z�O$R�<?c/�d��l!�<q*D�K27`�)�d"|�{��gz�}�fg�v����BG1�<���jף�nߚ�ƍ�]��&�"V�6�[t��i.�U(�H�$��ҳ����W�h ��f��>WW[��w�iޒ�[��nAB'�'��ˣ�DHK�Vz
���M�M�a>(�]�{�?1W-���+7��Lg�q3���,&&�5��2�B[���2���{ s������&�D�;i	�C��z��:���������b2u ɡ0��I�����T�z^���0������7�hCd?�J��Q~�N3X���껶ċv�@��z�V�$k>=ha\5�3w�<m�X.�o��b(R��>$$Tщ�Ut��i[��g��ŵ�8���[�.pFJ��lϦ',u*4�h���Rb.����`��b?��=��R�l��>8W����疇ս��V�u�on���d��Al[��w�Ѫxϟ��+@ .Zbg|�\�0�$̥sU�����R�B� I���@�����fI3�)"Go���:e�I>��<����y]��׬��Y1����7���x|�ԣc�&�E,�Mг���Z��yZgюe��L�n�$9����w�r��f1�@�\̀�
&�4gV�wI��	2S�0[�4FB���҄�C���㧃'"���[�z�����wu�k���72����dA"��r������R>)v��-F��'�F�
W�3x.Խ��]��ŵS����U�}��Q�	#3�6�3S���LO�K ��ei���73l�+ȏ{����ao�#�ܶIx{7A�  W<ݿ}	E�S�����0��S� ��r�<3�,^^ui�\V�D�� ~�� ��!��c���d�{�A���;��������,sYx���*�$����q�����+(ja^�����ޡ�D�o�C���a}���- *�|�7�r��#}�����G��� ����'�L��<�b��E�=#ꡎ��.1].����Z����`ᬾx�W�����U�|�~���s]y��s`{l,D���Kf��4��B�A����n��f4H��U�̊�(��,��F�C{ۭgv	x�'�8
'����2qv�s����~�ǂț�΂Ͽ�����o'Z8��O�9������evLbMM�u���������ϡ�/�5�*c3�"� a0�K��w�{�ф#�0B ����I��
ړ?u#����{�/lM'b�fp�0�{^�6�H��}�����]��(���^8��y�%��7�k��M׭|���1��w����L�C���χ:D��U�G�O���N/Wq���1��V���3��_�,�\۶�����e�^�G9��?_`l�E���-k�@�BȱVs�CB�c���y0��wmo�&��~����ó�۸ը%�&�Q]�o�M�0��*ۄ(M��:$��������3uE�F��|e����mӌ����ev�GٚC�ʧi���|4�uߺ��^�� ��6 v��d^���чS��%p�p�g���߄Dg�5�N�yU쾆s38�0��K@qeˋ�Q�pK8W���+�EnF��Fv�	�L�+�e�*���Cf4�m�Ԙ:˻)�l3��mB�v�P	������r��}2
Aɐ��hF�}�����?N8h@��q�>����sg�)U*q�r�C nyw� �p�.�U��|dؓ���:Fߠ��YK�U���F��5��O�ch
��dҟ���2p=UX���}�aOJ�n+��9�D�il�����)E�����|D���ƚ� �E͎�;^$�A@��eK��{���<eUg�S��7�T��u�Wл�ݳt���%����o�f<a���9	����~�����$;a,��
���ya6<��&0e����Hu'cXDD�<��� c����S�d��GJ��#���-J�nň�N�e����{.-���[l��p���)��/*�r�.�{���u���g�����i͕-��_G�N~�R�׹Ww��w�4��
�JӃ���U"���*��<��qx���t���~ ��6^�޾ZEW�2�R��1_�%�x���EF�ؐ��m8�B���t���l'{U�j��	X��l&��qpھD�Q�n��!p�WUq��r�D�6x�%<Pk�^��Z1�hs������K�>����Y�mh�aŞWD��9`%j�<l��;�qeY`��کM;)�H�p���~�����rF��(�f��rB�>y^ە�퉏p` 5�@8~_ͮM��guϊ�aZ��$װ�Z��Y��Ho�;:`�q��Q��_���M��u�,��ZI�c1,&��,��57b��7P��V"f��г��p�s"�n �Oq]��t�.��	V�G�5�~�4Q�M����׈XIS��:ˎ��mEX kv�<����@�W��X�r�D�[3��A��u����MW���(��=8�o��'�c����i�eQ��qHH2-�GtNge��[!O[���%a
�W}I��}�<�1�;#}��0�m!4,$�H�:�X��G��4���ۚ�E�֋��P�|1	5�(HX�6���^ъ�K�k���;qw��L��:��x�Ol"�DT_�=w(ʅ���nbN9�BcI(�yU+[��HZ9p��
Φ�[��~�]���z�z{ ١!��Tv�4��_� Ƶk���c�͎���y+��0ɂ�_;d�Z�xv�DV"E�-���n�$�_.��G-I-�|��/��q1|͟�pmd?�Jo� @�(��zb��Q�dD�4kD:���������J�~1��rW��Y�}����R��ԓpV$�=%����"�^7b�cZĠ��2(��8���D�FAs T\�����"�"r�dZ��S�����H�.�Tk3��9�p��u�>���3��G�^�1�;��ɤ�
_q7��r58� L� J�2H�`�Ĺz1��fZ�{ww=��Ժ

�{4(�j��Z�����?}gk��!'}�d��/1�T;(ΊC���kx7N>���:6Pz���aN�4290p�4���~~��U*�
��D��p)�BIyѻ�Et�mʽ�x�"yЈ���Ǥ�NT�ء����O�����3Ul��?ܑV�c��ہK]��Ţq��j�.N!;1�/b�IrO�Dlǹ����I0j 
L؜�Q؈�[�=�l�l@��l�ж۲J�qw�]��>/��CT�T#B.�=�G��E2d�D�5!mg�E�{���_zc���#_��FĀ�i�ژ��s2���<J���_��x�1%�� d���Y��^m����*��_ǽ^��/q�m��y0	vq��7J$�~e	��!�:����|�M/���Q��@�	k��u��;���l�lȇ^|T����3�� �\�=��"�WP��V�$�_��}:��V��}h���a�} g�Q�Ъ��Ф��6*S��V�!��+�B��[���ҨM���
g�Nu-������/�����R�\Z� �ꓙ.�2��!��hf[��cA�2�����ȉ�r��Q��w�����Պmt{MA�)������ .��
-�mt����nK][��iy�7q�p�.��ۆ\P���qNA2ޭeʧu�����I���	�&���J^���0l��Tj���v��]��f3f�r�?��Aۘ��:bQ�e�� ���A���ғ=������Fs7O�UT$�~#UszitdWM�w\!�ˎ��ʣJ��QR��wx{�!���g��\���K�ד��K����㾌��5�c�:�|����N���]��,�I(�h,�=��.�é4�����"��Le�
�' ��s���e
b�%y���B�5@&��R�%�ݭu�B%ᛁ�=��Ԁ'��[�ҋ[�	Y��v\4�k��y�N!����~��BZ�����ϼ�fHo��[�L����N��%�6��XvJ"���YrG;q��_�R
�S��cŦs֢pCk����|�d5=��#�	H������L��X�����uJ�������G�d�'��bY������[�)/zL�����F��)&"?�f��9qQ2�)��)tW�����uP��Z�����3trKm#u
�q��Z��9��q��Q5?�/&g`E�Ru��[m�j��?�Sq�Q~�(��������#��}��O�OM�6�)ΐro�~mw�m��}(&�YZ��a+P������$y�m�a�
S�E�;K&��1������5g��S�[~H�[2��Ñ$��E�#���;�4�Oˑ:�%]z���N��Q�i&��g$n9��=�u�M��̒)�ܰ#���[���Qt ���l��ǀ��7P�g�.�/�`����vQY����ug�F�^����L�˧�;�6�򥪀�3��w��r�C#ܿS�"��	�����Y�"q�5�����I<"�
:+��u��հ�9�����AO%t���ne�ef�	�[b�㖥x����ϭ%��@ea+_n�(�θ{�$��
ޟ��#^+���Zڈ}T�?�^��O����_�w�s}/�K�$����A�Fd���uD%��7 5�����q�"�L��3���e��]�|d�6�'پfK���g��.T�ƍ�a��&x�l]� �,�£W�(�������* ��@A�*�����h;�V���dT��EVE"X�N��W��<�b�.����B��26�*{<�;�bWy�&�az�Q�cB��(c��f�h��7,�?j�F�˧9��ئ���t��\q��}�H�HU�I,@E��Y�G�'���s�"
(a���ۯ�D��j�MPaXA����w��O�H̄",���/x���_��PA��s�^-��f��Һ>x�5TBr���+u�gV&:���7�p4�-�<�J��Ј�}��r}U�'�Fd����9�4���o2���o��tM��ws<[z�8���S+��:ײV�-������1CUA�ފ��[󃝟縬�[M�&0��8��N/���ɧ��Ja��
�Ζ?�We1��*y�bLkK�l���l��i���#�'Z�u�L�̼��&�lڌӳe���0,(�U5	,�@$�RM(�̊��P�����C�e"�����$ŗ�n��=�;����mHrZ;V�I^�{��el�IQK��u���|AMp]i4I��w�l-Wɰ����=�����]�R�f^;E������`���v�D%}�˽w�<�d�vmsff�3'o��XqO�ސ���j&��y���9]ѓ�rvj� C`2�5�airXPu�wV�ؠCn��rhn�PlG)-�`i�#N�K; E2՝5{��#� �� �V���	8tnW�J�m��
y�%����Ga9���ܬA���/J��kS��o�!#)3*��_��r�IIXUq�v����x�du6�����w{I�����2��������$P]���ѿϘbt��r:��3O�/�,4���{7ꋻDN�E�e�㹡��8����� Z��kk-�D��+�d��:>�>h'q�� �QO��|������k�._"��4%��[�*���T;�G��d����=�(��<�0#��*�.N��I�����n܊���F:�2j�R�*�g�ܺ5Dv"26��Fp����3���bj��pY]�0x�F�ܷe��42��1$jQϿ���)�\�Uj9��|h0���i���(��"!sqpݢP9o�?�=�"i}%컭�������/3���]T�Fu�������(�Y�"c���x�2�z�JBr��A"�b]\�9��!�U�5 ��^P�o��Ԗ�?����9ef8�9�7J�,�
�i��k ��X��u{�Gm��)z����hB�Aڔ�TXxuDM�k�.|�Fs3m�32`}����Wj[��km��mѧf,[��>	��qb���09?a�摦�ˆqP�-�0��)[�7Cd�ي��q �&���]������`5S�K$k���s�ŝ`�S�^�</Pt��=m&�]v9�)����@yuyO%��6&ޭ� ��҉�H��A5:����=�D��2���3!�����x�4-2�t��˛�����8��qR��V�+z��;��[�U+�0z�#hs�h�O�⧉�P,t�}!f���٪�H-��x�'NY7�"(�mF�,|-�ٖo\�ә�Ώ���a��Z��w�GG2yi���=2�l>��ͪr��B_�`=�B;���-/��m��"�/�I��ɗ��G��I��K�z�S_z��G�_s ��C����@e��3|�Zj3�୷>�k�~��A�����'(�R���u�t��Kv� ����*.0$X #�&M����=����z�=[���0��ѯ�A+�N���j��ǥ�N� "��I�-14�ϳ��/�gU` %n�5r�~M���rj��Gh��I��i��/��/� �b��R�,M]����{.b�-:���$�u�^�����R!XY]=5R�r`Ηoy|��%I0����C��X#������#P�sx9���M�v說x ��x�Ege��us˖;�Q������5Bz\V6M*�o��_�dA�,e��=��H���d����a�[<B�m�m{K����~�R�i `�-y�w8_�T+��xsއ�����R�\cÄ�/zG��_4X{�X�T8�C�A��O��zpJ�.�9f�ۙf���B����+�.B�<��i���f&*\M":ۅ��DPM�p:C!����_!KAa[����|c��TS���q��w�q�n`������١��g�NNsPC���#�6�F.����)ba�ԱV� \Ϧ���zZ�"ۚ��gi���L'h��1��e=��R����\䁑�SeH��T���ꉮ�j��#a�]U�4�߈Ӧ�@HQ����`f��	_^2֦w)T�}mMS26n���[�w[����^��ȋ��-�c I��^�<�b�p8h(�d����ژ۴Hz��~��7���r��`�W�ٸ�e����Cnj9Y�=��S�|B�'
���_�uF�Z��D��@�����4J�`cw� to�4z�t7��!��m��Z߃����	��keW�����lH��Ä�9� �d"X?5��"%��#�)MR�ϵ@���B�p��'_I�c\�ڊ�OL��'Sm��ҭt��8��4A���Fi�f�l��L�zN�帔Y��)����e�H>pw�\��~��y��k[��*�8=aN��[${rE��/R�)�B���3v���;y�V\%Wp��D-� ª	Ss� K��E�,����	�����Q۞u'�)�)t��YkZ�a	A�^R�/e����9�RB�^\�D�z�}1F�XC�RYw��Լp��9Ҩp���.��~�K�oٖ�0p:bj^W}���Yv%_5�t9��<̶�\]��6_P�3�b��5���'t���J8ҷ���ߛ�u�*\�������'�� Y4�4��mЧ��\g���ru 8s�4z��T9���KAC�/6$��~d_���Ǟ~Km��w�`!�yrm�uğ8�YG����vꟽ��]�1^$�G7���̓�a�J0�/@��`�`�]�ˊx<Is!���
e��U��U�{ ��e],J4��^m�r��_u_�:���Y�ΰ����#����Wb��;qr��礵֭a��J��睋y���z�x7��J�O �j�yʚH`ף�7┖Jx�g���Ƨy%��M��d��D*���g�%���N4i��~�Г�5��nS
bQ+�g�%��W��0\��u
����P	�I�FI.�����z&�Oϙ�"̗�{x},ٖJ�>M�� �t�~}�����>��u���nWH6�"��!]g=+_"\�6�O6z���CY��\�I%������Ձ |I��܊.=��>�pV��}<6 /���*��4b����tZ|Ǧ�<]x񠺜��1��y�oq�#|���ݷ+�c�qcHg�\O͂��Fv o(��%��.l��z���W�����8Z��v���}Z����)����,l���:�z���%9��Z��6��uj1��^~ԝᴻ�ٗ%c�\�xa����FP�a+�)����%��܄���W�/|�N�7_�R�RD�?ՅU�J�@�p;�v#b?6U�Y�e^�W���]6-4����� M4�HN��R.���]H����{��8�3ߘi��5s�|2��X���q�ox��=q[h>1nZ�`���5��d��M��bV�W�����Ƒ���p�sVD��-��Q��Mbz��1�^�����ga�:�ߴVRl�W�j��Rys7�ǖm�jUhA�s�k�С��v��pm:�I[9Ul ��>�!��7����
P����1�:���<���>�NMn_;��^�z�$qH'MÌ{�a�Չ�`�/�E��)�vZyO��/]I4ϒ��iS��s��O ��3fV�,=-?g�T��Mݒу<�ĥA����ߢ�g{��1}en�vr��R4ܸ>�c��{?����&����[c�^���j�ĊO��4ŉt���=�a�ܨ_O磋�$nu'�|'jU���fz?:"��_83���̀HW�z�W�z�T�x�b�����7Au�&?� ʄ	#uʪ�"�<���H�����L�M��=�yq�#Y���}��ٔ��p�`���v=����׸�5�=����:�e��c"ܰk*�"��U��
C�v�l���R7Y�������6+��^�� 9U�R��~�9�I�&�/ڽf(k�j�DC&�ȩ���>d���J���广'DvS�<�.[�F5z��~�, �^�'��cj�%0wS�ɚ�pz{�򭲽�wӜ0�?=��d����/�]�*��4ܪ���{����!��mB�/p2�#v�B
�)���@���Z�14���ny&\��\?�V�N\���냨���ՠ�}>�Dwpr��܃��6/����W��&ݪ�ǳ0#�*(wK����'�ƭ�>����4L�!��eC"Ub�F!��<�DN��r�#:oc�ny�+䜆,hMo�D]m,}��^D����b��v�+-�����gB�3�Mr�qh<��˼.�!,D��Y��W1�����q:-�'�C��&�c4�T��>��L��d1���~i@nb�Θ%˂؁�����LƎ��LU(�}��O�GK��m�����β���Ctd��)5`�����܈�YΪ�=/��g�Sd h����.�u�~c�pm,�<�UJ
8e�b�`�H�᲏Χ�/w�z���;g�E���z�i\��cGB�%�Q�#�u m��a}��%q������ƫ�ub��rٜ�ڥ��*�V1J��x�}�#��V�8�2?�'�*:�χ���Ij��b�|P-�<N*Q�/���-��`�=α�yě���0V�����k��k���d�\��[�W�U�f�	n2\��)�E�u#�z��<�WO�ͦ�d]�17D?�g�[���!m-�2�ҳ۬����L*�.g�$xL
3X\�^2���w��g��|J���?���x�O1ͯnrg����了Ts>��SZ4g �o��R����OQ���۫�����8\x(ۍ.���$�p��[�PCOOZ>� \d^4�*�P! Q�(Y�6�{SF�΍nڤ�V���q ^P�X���93�ke��
m
(��ݽ��4�[8.��DoXq�%b�V���bo�� �r�#�����`Ǝ��Ê��5R��S=��Ջ�ݮK��4�ڻ}p�r��Vd��@ԩ�4���fF�����ο�������}�zѨqܴ�B#3���_E(p���}}�p�B( ����i��?C�u��P��SS{���}��Sz0��cz�d���o"�Y��O"Mx�	������<�r�ɽA-���u[Sn"��v�U��R����M��x8|7�M;I��.fK�{C�sc_<�q��+'�J���v���j�>aG8��~OCޡYB<ό����ʻ�W�&�N���TT?��=���GK�X�R2O�d}�s.��n�z�)�Ʀ�WNr�����(卾U5ØrfLȊ�N�S�Qe�|�4��Q7:�^���`XkA�pC�{���w�7w�
�5�[s�*�7�l�&�����t���q#B����b��"G��T&�{
<I��8�᳎~ϗ�R�7�S����h/FC���xV�O���hR��5囖�����荅_�n��fl�1�&o���EO���ib':Vv���}\�P��S���O���(�q		}Þ`�M�Љ�r�H�3�:����ҳ=�ȩa�x�
��J"��*&Kۧ_���{��i3|N�H���;�Y�t��x1;���H����x����Q��Cc[(��3.�x�N|*�6���6���^D<M`�z���g>B�'n�h,���Ym#'AL["��fH���H0�Ƨu+��?�4��Nd�\&��� ��4w�0:�2u�/�*�9�7��FG')��_d'�h%�"�}�b��[�������3��R�Vĥ.����fM��>����w�I] CW�
����A�ώ�w����݈�-�)V4���T�'��I��e}� U_��0t��CPw)�Yb�
�|�;���B����i<��Ȕ�Ҵ[�F�C#�����-q��՗nLIz9�r�a���6��5��M]`�%��À�{��h+d��_����3�����)Z6\��\�}Xp�4"����9�tm
w�<u�ŜC��п�٣̃�N��Ǒ��	��b{���֟i,ʉ*�i���YoLZ �!W5܆`�r���?T\~��,r���BA�t���Ҽ=S>o$�Φ����R�S�)`}e�__�q�j�F��H�CW���˜�b�=^M�c��T1_k�r=�pӪa�@Ko��m��;sT�5���K+Ј�P�{@23����D������#4
�F��!��!|��ǒtbݹ�$p�r,��ϝ�c��ݼ��1���B2�O7;��4�e2`���t%)U��5`M�6'-2���4����}�Q��<H�RjV��8����:/����.�32j@��i�<	��H�mNVK�������H�SyB:0pA{,�Tԫg_Xy�x��^Wj�Z;�*�su𦮡u�c3y`�F����d��M_�F��c�F�?y&+�-�W
��0��,�6.�%��1z�m�˼wd��j'Q(f�_Z��{��:�<Ǒ�)u�h$
 �G8��b�`��n��^~��:�Q���[Ac>��(�v6!k����N?z^�ER����o�ǎ����Z5���`	�U��D`����~~��*���P��I�& $S6D���4��d�_�C��"�
A8Cj��;(�D����4�~��T:�+������C�������}{d�,=�lj��&�͟�۝W�`�8�EUZS��j
�[<N���z��Y��.�-���A�j�fo��*�{ ���Ƭ�i�3������F+�����5��#���C�-��6wwr��Z��!���^��VK`�0�Zp��ﴽ��1Q�5�@���2��-Y �QB2�D�ݣ\Z?:�	�*0�o3�#�ݡ�9�Ƃ'`��qq�seB�8�\И2�L4��� 3
�� �f��x����A�؇����͇x�@&I�H�ԏ�[�|M:i��}�)���y�=۶�:G�V��okޒ\�i��x��wb�1��,[���료��b��:�I�ơ҆(r/?�e�+���c`���\�#�8r�������$���D�v���R=.yω(g5ϸ��7��O�q����n!!�@���,��}A�ƞ�>�;lko~��;�#�)��^��;w�����V��k(\N��j�����.�5|HPpys��P�$G}�2},��D��w�̗��8�dX��Pչ��W |�0�Y&:f�.ڲF�ی��谯N��q��<CJ�fv�6�y����:���u�"6�c��d�K}���82Q�sfv�c� ��y� ���m���p&y/�9���+�q>���icuu�Ŏ��۳�-/�a}�����G!%N|P*9_Xb=�F}[��Q�5��?r$�ݜ��	�W��/\$|�3���N�:���z�f[��Dq{��ą͆0	G�m^�����]p�Vb���ˏ:�l���KĿe�_�ܹ@���K�E�1s ��Of�G%̩�)(do}�%�^�9�k��� K�E��[�]�_)�L�e<P�w�Fk���(�a?�.lyp7�>i3��+&3z���G8dÙ:��f�՛�kg!�tؾcr]$���Ð([~	�Bj���-���z?L�:��������h)�V�5���"3���ZV���e#�4�b5���)b����S6=����>���I\(G)����ޙ[B��!�Uh�]/�w)	�i�bt@�-�.c��Sv��u��e"�g�^@�(�˔�a��,��%�t y�V�n�sl�(,���ON���C#�d������BuI��p��ޚ�\l�*N���8sp��{�a{�Ӎ��|T[�pb8�̎'�tr��S����Y���'�����F����ɚ�u%� �]՚$�<3����a�{�̝Q�齂;�������.�~����NQ���įLy�-���>4о�����~���Ղ�b#������W���qJ�ۋ�Ծ��kne�����@E#�%�˝���Mڎ����MX����¨�Sy
<EMS�a"��S�$�4�EK��s���Z�ci?��ؗ�쥲��Uȕ41
�~P�f�Zi���>�����6h�����|Q�9����+P�x+(P�è~N��DOH�'�~��PcH9�F0���]��&�����]��5���������u$��7*t�RvY��=�=�<5L���R$5����h��c'N�n)c׳EjN���S�`[FC^���E(�OS��9�*;�!r��Y�`�a�Ŧ{���H�X��}�)�M"(b���x���y4�2t�E����+�#˰	y(�ɵ�u���?�F������\3(��Z���V�e�����d ,1R�wt�����X��O��Fѿ��)2F�&���([׀���b��_��R����R��y�P�VN�э..2��2��P7�-,jj hQ���ǲʏ���C~6�a�:eU��l|<C��[�+I.�����*_�@�K�XX.�b��lAΠ2�PJ"](�;�Ƭ2�H�	�OFj��RR���fd?�e��m�*C�Q�#@a���AYaz�ԓ�-�-՝��^�91.6��	��#(���8���/Ǆ���tZ&�q��)%k@zJz%�S������sQo�?�!]K��r?����a������wJ�����Ɛ�0g�;>wM���37$O��ي�ڊÝY,x�Tx�;B�n�0�Wĺ+=.8<8'������9r�^�<�o׵N�S6��k�a�R�~Ωd/6m�p�{ATe�ϬQ�T*����$I�$�t�VPR1�֕���a�.%@P�ŉ�~�KE9И΃�1�]��v����V~)<^z�~�OQ��טː6c��	�;ː?�a|@�Bfa�F��:(Z/�=�p��G:Ƞ�C��Wg��jia}�a��5�F:����x]h3aU{��Lu��� #@ջ�2z0�y��Cƨ���2�qA�r�����I�}$'�݌7����^ �C��.ZN>��[~��X[)-M���Rh!=0���=�v���@���4E��󢿪߳�v��HU��|�;7����K�ƨ�T�����8�ʅ^���WF��5!�W#Cb�������f��d�?�4�8Ѱf�;��#�
L��1s#0�v�:�,��v'q��n�m�H�T�^ˊ`?�o�g�l�9�qc�u�@�/��q���ALA����8���T��LuN��7��:���
��8G�<I��"k*�J�½� ޘ�r����~۾5��4�\�'a�,�t�Zs(=Z�Z��0w��q�fGgw��Jd I�V�T�gA���^��ž6�Y@,�"pu/�Q^;��ol]SF�j�������y�w5�zU�ؒ��!�i����\���s��h���N�~�XF`Mv!�[s�۲O��]m���ӖT�L2.G�P��`0a%#=ױ�ȋa��bˇ��ü�q�W��ܓڿd�m���u��~/(���͊�A�Bf���׍���=��!�w�b4��)h���1��Pa��/c�	ɐl���r��၄�L��'��>@��/���wZ�7Q�N�(�,�W�y�ͬ0�?�@l��^����@�ǵ'��a!�ڃt�|��	ī1���D�(��F
r~(|
|��S���R#��Lp�θ������\۟�A@
_u%�H�&�s�B�a�T�mit�I�E�E�^ʨU�Ӄu�D6Dbz:����Y+����|��@�L|�H��u�*��Vd��~�g���)I3s=1�b��:y�#�PG��<p���Q�W܁��p�^�ɛ/��ާ�rm��՗h����v���u9����!�^�y�k���$��5**W�f<_��:NW�B��}�x@�k
���y[�YO�^�\�F��b��$���F-��n��=w.KE�h����3�ݠ�QLX�E3,�Ӳ�TeL&쮜� b����c�ڙ����q���$�P>�+�f�7�u�Q�7�Dp������cf�I���t^��;�T�u���ً�E$�j$�����|��~tw~4 �m��x���m�QZ�S��M�L\>��������c{[��l��.���Vd��G;����W�~�%}J��j���\2���V�w*�j����Ê|����i�ֿm�r�H�}K}x�o�]�B�bI�CPa�f����S��ީ���Tm��r+��ƑԊ��"l��Q�F�b�c^�,0�4�;�M@_�Ë�*�4g�{�헤Q��Ѯ^�G!
1�y���ė�/�L��l�~��ϫ���r�����X�9����U/�,"�K��/-�@jQ��IV�<��.:VV)��Ǿ93��b�6v5�i��\��¸�HG׾���p�=L�Հq��4~�L�Y�Ov�q@�=.�,C6͂���~H��o��`��h���� �VM.qxRU�V)yG�Ry��
����d�k	GS�:G��q��,Qd�w�&�WF��bB�c�ڠ��JG�<n�� �ù/:$۝귦�"6�����|�/��b���	g;��g3��m��&`�䩯�0(T����a|�(�ըB��G>�f;�Qah�f�C�Xى�_�+1ڻI�א�����U�P�Tk`�;�L�x�B/N��="M��>�땾ߡ�<(�v���9sl�HF/:o�X!�/��#M���ٟ�P��x�aC�m��vLּR����`�y�bY��e�U�.��#͆�-5z�ҿ=#eBx����|�os�c-N6��L-�{�q�f�J9/��"�Z-(�B�~QBSܽ�l�<�&����s��* U��)"b͘Q)ug��0ME���C9N�`�C,՞i(�o��4@��{z%�^D�42x�	o�� t�,�87w�V�U���8n S,��q�{�FG�+@�\F�)��16�N�
���0q[�B�te����e�z��o��D�CB����%�v!��9ˏ^ ,�X��j�T-r� ��Ҳx�K'�
�n?B\?��R��ǹ�V��g�=�M{�d�����}��q_'��K�nK1��N�r�Iz�*^������t��%R�=�Y���mm-�K7���H#7�;X"�㋼.O��w�J��KAsΜ�w�^�n��Ɨ���(t�{d�v��T�X�k�o��|ny� �ڷU�j�kp~
o����FeV�4̂-ܰ�<�c<�a<;8�r��4�u��WB@�����*uA�n�/>�Z9N3,ogTV� �R���C�&E�4���90f�� 9NVA�[lFU<���w�2>�E^�$�^	��^�v��k,A��%�8�����Me#d����5.l7"�Ћ�yL͔`2�mP2 7:�<����C�%�p�<�H9p:��LXd���Aqpnh�p�4��D�n�s�>Iz����%���.�(��q^���d�����viGP���%�G:�z.�_�Q�`��횽�d��R�3ey���]H���4�3>�%���L	��xb���wc�ůn���?�sQ����YA<�*e;\�6����?
�~a�+��J�l=D~-	7pB��>���矑<z��%��V]�����xJ��}'
C�l9	�Sź�7W�{]ll�xZ���Y��:������$Y*L�	�M@]�Ki �P�2�����ҢЧQ	A��Z��>��[���!0�uF�?_�5e�S	�&g�5� 4��!���&��k��qu�<Y�qn�U�t�3�$t��u*up������W��*i��Oͼ5�W�1:@QԻ�3* ��x�� )�w�oK�nVj�^�#�r���-9F�N���`���W[˖h�[��u?�������;�C���6�lvB�-�N�UJj��B��ahP��Ұ�!����X���oi.�����_��w����K��B�0�������|����G���Y��bĝ��ź��(6p0�U	|k����z<w]MVf&6Μ�G�<���k�dy�z�+m)�Z�jW�hSr���}ρ�h���{���H�6�Z[�	9��wʶ�.r70�P�ISkh�z��i��t7f�ݽf
��^��س�i��g���������.�2��9Ei+����V�����)`�����Vs����\�d��.~�S�ѢIƍ2P�t{0DeK5,�y1�L� :V��=p�{��\����wK���,Qy J� f�uJӞ�3b)�|�.��T��^�t�͞��Ī�Y2P�5<��Ȇ� h
�FT���'bF����<b��+S�H{)h�����Z������Ǽ�����?���|��cE~~���ݖ���rQYK��t �1Ii���RG����I
ᇳ^�ʱ�9�`��)?I�y��q�C7�r���=>E��[-�,�o���0堔)8S�gV��,����r�l��qi	
6���ߪ��eY8�֗3�z����{���$�\�9k,	��*�:�C��J�wk�����(Hx�k�L�
<F�!��+q�\��[��ۡW�
�z�_��D�0?/�N�����c����%��Җ���
h��������aZ��,iU��N��E=�"��3(y`KgT[:�5sjY�<��N�<+�E�3f��b�g���"*�t�x�v�^Vs���gn,�F��xC���}�T��X�)���0ݏ	̢@�:���b�����V�����}�$rh�Ɓ���f��-)�-.HRe��>~v/l$O�\聽��!�Y��|�"�7�v�0B�Y��%H�m��6��N٢�_��%�~��fY��	onr4�w��:AIG���m���&�����iU�!ނ@�"�*��-N�(濓�}�xo&!;2��\08�K��jo���F�p��d�̞��K{�\Gr���w���F�k�F��2\p���̡E��!��N�^g���Ǚ� �I&8N�@zs���K�8@M�O��D�Kܢ�΢��3�M�:����6�.l9��{�\�<N~�O�ƒ��j���^�v]�JJ�R!Dg��%�����"�-�g�O$(����@���ʮ�8x9��"g(j�U������F�&�^��#0!L`a����2���VZ3l��8'��Ǟ>g+T�]�\$
�[p��BtnE��q�������ٔ_�H��2�*B �Fp��	(1��8����5�%����p8��&C��C&Lo�^�#��о��p/|V�u�*�&��'�қ�J�mwjp�m���C�)8+�.$��7�qx��8ON\m�����;�^Ojw;��<�[����Ղ����qfʱ�Ьa[Mk���^�t�sD�� j[�wb�]�� MG�bxX݆�x/�w��
o��S]ű���À������0J5�=u2Y�aEM���/�y�<�M`��G
�I�'!W�z�&]c �����bg\8��b�k�}��u&�{�	fy�i�H||���W�n��^�h���u�o��� y�U�B�d�"��ld��;�&i���9.��i�*�w�0��!Ș����0����s\�ke)C��-���+�w$X�g�	�
�,��1��o-�P���)�=	_w�F��;>�|)���<��y����.�;(�Y{��;�A�X�P=�	��z��5��KA�Ų��o`
-\�Zjpa�-E�.�d��[K�V+�7oQ�@��.{�BA�3�b¶/P˲��L�J~P�,vS:�<�=�g4�V�Ȣ�Ll�M ���_\�â���0е�G�_5*,�^5��ږq�zz�؟M�I4��yݵ�K>,��Iw39��{�A�<*��u��yS��{ �e�]s�+����B-q���k����.���ה#ga�1��[��s�}���m���$�b_��j�+	"����T w`f�.lj�<y��'^��`H퇾9�
��6D�JؘZƁ2���F�34�&1��u�T|-L�)K]�Z�n�ȆU��
��W�j���%�jD�T�$Ho|p�ŭ��B��c_*�@��$
.y.4GK&ڣk�m��c�?]Ɓ������ֲ���y�g����3�$#`ơ��2��]�5s_TN�����i��,Ȳ�M?�\U�&�C�����e����jI�>���y8�W�����*�>�h�h��Ԗ��c�I "��g��v�n�5
���_~��H��]<]%�7��{���z<6��]���P��С,�Y�ܝ��0�2-A�r�~\�f��ƓYejeĴ�T���ⴿ98:����>N�NGd4,�	b��~7�A�P8Q�Lv�q�/�S�?��ʜ��@�b��:��'c
k.��(�b`�5ƞ���ơ�"\�J�3<b5v_-�[(�'���3tt6'��x�X~��Œ���Pr!.�&цO��CT�%R)it4mp|7�Hp	���~ �-ᅗ*����_r�h��W���|Ύ��zP�AN<�|���=6h0+iDW��=�y�i�[GMc��<����Ih������KsZ)ztC�O<�Վ����^��N2M�u]�`�|FM�K���i��u�«C®��2	}@��k,^��l���hUf�1������+�	�\鋍�}�b=$<�`V*;�^�9Ca����3����$�@�\�.�j)��O(�.<�{�N�$1�r���#��������?��M���?��f���ߠ?	JP^��W�C!�J�\ꫮl{��������\w�*�n�-p�����5B�}x�A .k㧉��O�6�R$�,���x�uU�3�B'\��LS!=z��k��gb��H�h��$�g~^�?,�Pg�A���N��V붵鲓]I#��O|��rr����������ձ��؃ `�}��`^(��&?��b?XL��_DvF�.�~�\��矫B�(TR��p��2�.*1Q������w���j��*������ �M���)�.,�Kũ1�h��FZ�&8~AW!9�%M�l��{��I��|%s��z�y�|�1O�@ c_�m�8Q5���0������oR �t���	���`���d� ���Z�W�����?���-�����6����(bIqH؉���Ԗ�(��~�)z�41���'��B�HW�CFN�
�1��8�7���t,����%C��]�������D��E6�%
4J[�1fr��[0�*�;�s�+���U�N4ei�ډ����ޟ��R�D�y�I����s�X�ۃ+M��ZB��s]��ps���Q~��a+d؍����)�s7z̭_�)^욛6e�\`yqJ��f;!��Z��͋n�FcP9�C�;׆���g^aƖh];Q��Ya�R���:{�#�qg�g�~�eA`�A�Fv�,,����7��AfP䒻�(����������Xm�㺮��~��������j���֪Z��3cT�N�Ƙ�����|���_?
<��H���]����^�d�֧��+�a$^�#ˤ��q�	y{�H�j���v[�KgK�dq��{!�|^I@���Ծ|�����EŲ�Ga�<]�Mw��UvN?�� �V�D}ɲ��f��?�q�7	lU�x���:�GD�!� ��h�������&�>���� �.�>������}TC��ß�l���n�)uG���dO��+����C�EBހ ����d������Z���d��- =���/��j����X��FPƨL��Vo!��0�W�ՄR��[���!/�5�x"#	���Ъ�Z�䜧_չ��^'aZ�5Z�4\(!mԱC����(:Ε��g���tj	���V,��%���"T��e�w�:]F�ܚj,ƪ՜�rY���!�(e��D�1�A��W��\��j�L�NZ���$0P�