��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|۶��-�E�����^�L>Ԗ�Tk@��ȼx[�ͧ���wa�d�y�~F����C�[M�P�r����s��*� T������/���ma����Gp$@�ћ��Il/&�f0#޼�����p���X1b/��]r�F�>`�Ʈ����/���Z׻�pc7�8�`��N	�����]�sO��'V[��jF֕2R�� �������>�7�S�w�9��O vr�� #2�)�
�~��K��b}Z~���}���[���*�{�I��'e�4O��?�w�A�����m^`;ڗ!#Jk:��1j%U�à�ZDׄ).G��R��`���ЋC��'5������5��(�y�צӅ��]cd��(�I��5����l��c.�� �Y������'��c�ç��-ѭ��W�}DzOJ^�����w��E���:���qX?�*��{�Q�4�#ٗ�Fa�jj�2���7��:|q��P���)��B�=���g{�8��%/
&�(%���H�C���v��21�vFqv�A� ��AE�o�A���ƈp�i�	���<%e~�L���?⧯�ˑqy��"��~�2�d�Baƛ[9�`_`��\K�SD  �,�5�AC��do�+�}Y�F+ccm�6��mEFV�DB2��C�e/h���%����X���g�%pI��1_-8�I��7����]�kұ�6F|�\�i����z�7�<=�+��yr��>��@>0�A�4
�!� h�M���;`k'�Ԑ���?<�&0������T4"�[x$��	���E9��y~�x﹜��^m�pT��5L�8��=���XzCaҳ�[Q� 6�U�������jK��^ͯ��GE��̜&�_� ���=k�mFj����7����(
�����3�[�m�3�0�L7�q]��H�ɠ�&W�ʎ�9�>��'�T�F�+��`_��=K�+0SP�8Tua~�[�H�8���Wn���1,7ZUH�խz0r��N3L��
\�v���DT����] �%�;�ff���P�>{/���j��w�$�P-�	���*��:����J8�m�!����뼍t�DU���?�T���N�c���(�DKX閷4�j*�	�����kb�"8>	�=�D���D�)��A�S�"���[}6��ބ�XY�Ź�Hj�#J-=���X���fn��OŭrqV@&�j�]Vn��}����/sK�'��bn�B��y�JQc��;�qm��Zʪ0��å�E�H�^ ����A�ܡ�2���5g	A��=��yFٕ��R�z�z �A�� 0��\9#�>{_�Ӕ)�"�p\������N�D�N����z�Wi������R��n�ؕk���
8�G8��SȻiz�pt\Oњ�A�9c����~���a�5�-l�%��I��M��}��ZSS[v�q n3Q1;�r`�[T. ͉�a�q`�It�VW�<��u�_�U�Y�}���g�9�qS7����� 4��!�?u�_��@�=5�ﹿ�&�&�wv�S��Qp>��d��MԽc����0��Q��8�Y(�r�~#���n��8��G9���?Y��vPX4:��׃�=m��B���_h��(sc����[g��n��x�*qVU�3YD-ч���u���(�zX�!Q�^AyO���FP�W���su�.Y��T9�)��yh�gΏ��i����|�A���e~y����^.���%i�C��3�?.Ӵ���0�R���	aˮ�-Y>��#x�\��-f�N�`�,�T4������f�3�6���^{���;��c�����	d��'�VQ�O:�G���De��|��Gȕ@te#?���h��^�xS�8Mc�"�v~�
�9W5�����j��Z_2L���p�KlK�q�����}^{=��� z�Av'	�%A����-9�A����|F���"�g+��4y���婵ԀN+�ܹ���I#��� 75&�=ac3���%�w���xF�<{oR�������*����L)�5|��d_�5A.��ȟ}��u� �?���j��4�
zI�h��I���3l�� �tV� rW����Q9y ��ܣ�^�,�`[alo��:e��M�=�`_W���E���?����}���ΊY�/!� W	?ݯ|����
�9�so� ��E���':|L>pZ�^�I�r��A���H.�g9	���ګ�HP����f�n���8~^m���@*�Q��<K}C�Q B`�Ƶ�Ȥ��M<�Қp	|��d��K���E��|rq�2�~̲���T5���Bd�R2f������T���؈�`H�[[-�sJ��YPŬ:n�%;1��m%��ɪi���ŵF�E�_Wy3'��M���ꏝR�D,��Qb��E��Ex8y.eS�j��_UT	�Ɇ��pv�D�s�QR��mY��ȣ�JF��ߎ�oԍ؟�&�Ċ����}t�)u�y�N�4��_�f��|��:k���u`Z�~��0K�~�4ɤ�c����[���Шl̔�Y���Cz^�`T	����;DP�uM�d���<~�	�}e��W�J��WS�?��ri��<G�D �ڪN� �X!��/��0�V�F�m��M*�����H�i.���@ރbM�R��_�;�����+��b^�[J��]}}�Q��!;����۪>�a2��������{�BSq=��~2:���*w�А*|d>}xڰ��U^ަ5�"Ta�!�o��y�����5�#�ǈ�ò�Q��F��l��}�"C��j�;wS Y�k�B�7����pg�`�ʼE���K-T����0�CMa\L&�[`R;��W�g,��n}�ҝ嚡*����NG2��T��+�C�3Z�+���T����Z�\8�R �Hqm�Qͧ4/��>gE��׏�d��>�@nd���.����7g�]f�J�aT���'�t�eL�ɧ:�H��+�τ��-4��I�=Q�E�^�ٓ�/ K�F�CN���cz������1�ck�	��q�h�X��lcT��d�R�ޒ$��RS`�����)7@�U�l]� :n�v���6!|}4㚇V�7wt�vYn��_�����VE����o���&Qw�Y!�ǻ���<�]����EȂzD�Utݏ�BT'��%Pa����0�-7���x������}��;
Ί	ǂbdy��W�.�� ���7S�����7�~���[������7o#��`F������N"_���Dl����̨�8v-��j���\d�S�w @JǊy�������]����8��%`��C�.X���	RT����@ ډY�	u��my�#�O���c��P���[�ûIL�[-,�*����W=S�2�5`m�c��e��ǡ���o�	���i3���#.�KdL�I��I����H��]�˛A�n튆rjo �cy�[�a7�9��N{�D	��0��x��*��K���.[�]�B��12���c��B	ؒN֯Mo�ى|�)?}e3u~C�L� ����`*��71�K�(L��J��G������*X��*W3��5
��B��,�_�8�p<���a���ðT/��H�����D��V��*G������B�(
q��AJHH��p�c����S�;�� ji|t��~�^��{ω���CIRX]�z��L�d�^ٳ	�-�����PD�p�qYAB|Tʵ���S�/PS��䐸鼾�;!�T�l6NfQ�vo?����I���S4���F���Æ��)��ǪW���w�Eu��R�E��������m=�!c1��?q���>\�/
��Y2��rEe6�NDa�����9��� "Jز�9�ԉ����q>xI���ѐ������
�$�GFt>�3
�����F�.|x�z�`���|SL6�W͛�{���OG�C���_[��w1z��\��(_�s�َ������ܚ�s{�Y�TE3������u�]~B�(b;����t����q^���n�Ԯ����G�4k�[=}#ίL��.�,�ŵl�-�\6<���{�yL��s��3Ŵ+E�,ķN&��W�~)D�I_i�"F�vJ� v��MԒ��h(�7��;(߹���a������]�+���?7O�eW���W�<T���V�@�nA���F�{��xy;
��@���1`��MHl -=���{��W�7����i�!����;fT�8� �8�����|�>�"$8d�8�}y�5�ˢ��$�1!C'��ч1�%�S���pYS��O��/&z+�Z��k%��ᘌ�R+��sZZQ� �N��xM�d�={��r"�]H�������|�ȃp5�����;���	�0��2h4ן�x5�d���J,ŝ�흋O��"�u���a��d`���՝��@ϝ)w	pԅZ��an����踶Ȗ��(	�D���k����A5Ԇ���������{_��B��W�:�;�O�E6_�(tM��O Oy�C�"s�âs2�g�����/#M�ۭe�I�r�/�g����#Y�7ʩ����;bI��{Y�ƿ|�y�{F�z��b}��Mn��cSQ���2�gb��u!B�wP��\ы�b@[[�ew�	�����f�]a����H�_d��Nf3܀��������t�þ�?�hY�ة�{�����nK�<�	������%*���A����c�*1�
�W�%_P��(�|�����[s
R̠x�b�YXd����D=�7%R�p�b�1Ӄ,��}
���vmY(T�=�c��Bk�j �욒7ueh3�h�L�m1B��<X�qi�g�>�L��D��k͹CUʮ7����������XA�t����0��^/�R_"J��NՌ��G|�'�����"�1]��}kf�d�Lpun�Q�q������bN%���Y�u�K���fj���a�̸�aQ�cm�#E��(t:w�FK��^�n����V���'Q���H�&�n�7e6�y&��f��'䀌l��h^R2�]�}���C�1�*N  ~ح�B
8;��L"b)��r?[��R��Go_��mY�t.���l�P��翛�J��!I����ƈ�ůW��r�7n5�!�<)��G��q��	�?a��U�5��X���/�t+(���!v	.@%]_���i�CiT�쵖����h�.Y�'�n��l3��sF>DpH�ܘ��3a�.|X������BܼN��u�gڎ�y�$�J�Z�HW<�kT]��; �]ƫ�w;?:{�T�k���/g;��q�̍/D},J1S�$ ��bd�Rb��if�}�{�	�7Վi����W���H�~�F�����PW����lصjQl��.��)�ЏLV�^��^���o�p!;P�E[p�j�1��K*�C"�	1Kgb)@`W����1aWkN?��!V~��k�V�	3�Wre��x��8)���U�!������v"�M"F�c�#���o�rF��
H�b�7���_6ܽ��J�rM}�t[��\�u*�����̌�*�A�Q��%v.a��z�;�x9�(d������v"I�q��׾\���]���PSx#.��Dz�zݳX�1[������2q�� ڥ�R��L� ~�,*�O����J��`1#*�"i$W����	T|��
aY �w
#��j�Ԑ�3 A|Kk���r(<z�i�=n��4I&Í����#�*,�zv^�
,�kI��'����P��T#)�-���wۖ����=VɊ����t�5��Ͱ��M��~��
#&y0*�2&�1�F:�#����4@�1R��~��Ѩ}�v殱 S�֡kR��厜v:��p��h�Mg���c�#[�N�����;�8�I+���2����B��d^�r8 ]Q��]�N���Ra�Vqϕ�)�"���T����������I�uL*=��*/`�ʈз���E�}Cn���ˉ�ܸ�g���J��E�����ߗ�e�O��{ͫ$��$����7{1ͬ����)��)���1J�4�u��7e-v��$�k��Z�v-D܁|?q��Vm�55�3�t>M��d_=$��g����J����/��V�K��:];pbZ��O5��\f��X��F��Bb�n{C	���YI�������4G#�De��m����4p1^���>�?���YM����@������h;��M��z>4��[I��^{'��u�7~�!o�TvUȩ�1.ɔ�<Cۉ�����HD�c��+�/��vAWA�C�݅ 6z�w�(�j74o�j<��XQ�6��!���-s�^�ǻB�KT��H���.f�x��M�`2Z��w�*��gBI��^ݻH�P�0D�y�����^)�/Ta��6(g8���K������1�]�����B	e�l��&���0vn]`�Ri��nƓ��H�Q�B ���%2��$9�g!g, E�y4Q}���.�]��ϒN`�f4�F�;tF�ɡUd��c��3ؗ~�������R�_�4�X�q�Z�|!�� ����JO8o3<7�?����|b�����xy/�B�6
ycfnM-��V�H��D;qm�P
��{^��ɥ�f$B>�c��U����ގڈ<Y�hw�V�Ī�H<��*v�t�2�!`�mTB�6�ϸv0[�����I�����8C�����UYHW��UB|�:_��t\���1dDJ�Z[�.3������R KV�D�<�3m?��t%%�>��<��$о�[��o�,|')nr�����F�#=��ѻ#,��ϔ.�V@#�!XK+�z��"�xGiN�5�Wm��>�O�!�I�
��VNGZ�'�|�c�7�(*Ǐ�uH����Ϙ�tH�� ���Н�1 �D�����]np����Ft7���Oo�6n��[�e�{�y7�t�G:��@�^��#����T�.�1Y��s���ׅl��V#�7���Z^2�,��b��~)O<���_m�&�d�h*�FM�S�O	�2�������NP�u�L�.�i�\����8P��[�2 ]R6����q�aNÚ���*O���a쥍�t��M���@��X]j�m��3u�0Ѐ3�{x�~��0������H�����7"��Y+F��Q�6��Ӛqo���%��$=w����gs��Q4$�ю�}�mW?M�|���Yj����4��U)�RU�|;�@0��f4�
̊預q�t�ie6|�?�0��yh�-�.mhV�:�)�OM��y��A��@�9SjV0��/�;����w�W�oϧF�Y��ʩ������;�ਨpr�����u[S'�@��t�i�=H�FK�f@>��J��CkL��՟既d��I��������P�>P�������Z~��[lS�Hk(�AH�����.��M��Ԍ�;r�>#�4<}u����@��]��C, DV��	Ȭ=��e+SsI&�I����ܾ�x��>=�A&��#�Ǒg�k߇��m�vf�CVi��N���b��������H�aBhA��4����WK�Y���/��c	�!O�x󨮣L��o1�2D��޽�%�MY�h�l1�?�α[�r��� MNy� Y�u���f喝?T��>Z��oH����3�
y
��`�,�j�S�2em�2�M`�O����leŻ�
�gx����W�RK���#��`��������<~y����pO�q���c�<6�7�w�LU0Z�j�f��u����m�I't�髷1���!G�}֛��W����wT<��"L�S���+��X#���'���:Mh��O�7�"�h��pýƃ׹���g�HW8A��XF���hc�\�C[S���$��\�疋���&�����h��R��3YS�8�L��nr�QF�U	xI�-�)\eS�oV�Ǔ�R=��V� �fZ���8�I|Ȼ�*5����Z�}�J���U�;$B̠�]�
��:n��X�M%Y�_���v�%/�u�����x��[$�E�%G4d\B�P��Sҹ��;�lYM;o��I`��h�Y�wAu�d�b��}'E�dIr<��_<q $I����ň)s���풳=���� ��*^1�!����� ����o����TW�z�둖`�w>���`�9a5�aC����+|�ټĖ�� �������J�Y��1䆶�ن����M�����`nc�{"K�sm�3�X�)��r#�� +IFӪ�(��D<���̉Y�RI���-�0bY��=hG'D�et8�~h��BCJ�n�/S�Y��&�t|,6�6%v{�݆����u��;%Q����7z[ۍ)�h�s~+m�<,�4��f�'�o���	U٭ 1b9������G��ذ��d�����ʿ���~`�A,��'.�E�v:�����*��f��/�|���rr��g:��)xN��t��ء`v��:�夏K�kL��������Y������kP�� FW�����4�dQ��1Q�yq~�Z�Y�F؅��}�[���� -o���g�"���ݙq�6�Ė���y�a�0�lI/`\m=����i���\\9��o���	Vf���s���pj��P�ʨp�� N�J/6�ćt�R���?U�p%� 8��v����޹�==H�l�\����R_���d�k$�R%h��P��������HVf��<��Np�.����V�O�?��&�{���j4Yt޿�d�bMwR���� �[�% /�F�K�Y#A�а8��E�3T�L9��;P�l#|�w��=و'f:�y� ���7y�C&��j���4уf�&��H�3XR�8.{�H"TLY���nxe�ǳa�:�J��~�`�|��uh���JH�2�9��.� {�N��,ɢ�pS6w�f�B�Zp1�84�TRQ4B���ʳf�������D�X>��uIK����T֠����O�s�n_*��k����q�����9XҒ	�/A��U+nƠ4!����3p�0����>�at������%��G: z�����@��v�G4�N�5�bB\�x|�/�5�aF1ȉ\�����`��
�30�ӄ��Q���<����t�$��K�P�+�s�)�Z������3"M9����|��<H��Ъ��Vo�E�-�x� ��� ���{�Y�b��	2�*O̑!l69h�_|���x9�vX�Rv2����i;��,*��|�)e�%���B�R�+�?1Dj�YF��^�
�Z�.z�-,Q��~���]�τ1�����/\���&=��$�G���fSm�|�M�h���]LJ�K��&vU��ޟ>`.�|��!KR�E����/�*���`��SU3��[�.%�~FA,@S�Akϯ�9�m\+mHdk�?Iϧ��n�:�P62v�&Ro�����\���1����1�uv��l���S�]^������۩���[�
I���K���Y?i�+xw�L=@�������Uf���3�3,m��U~u]*�4O]^��eL�R�a��B�l��A�w�Ř��?�X���`*G+0�%)��h��{w�����]���D�/cɂs�#� ��0k�,h5��0*a����s?P�D���`�~$o���A�cJ�فu�V��~�7$��t�;Ȭp>,�����uT�q�K��T���M̚��-?%�P�T
�!}�����~��DQ��nL3�/0��A�E���h�gH�D�̺��	�[¸��MM$�6��Coh���k��?Vn���g���YJ����(}I+/@���$��d�b�N�5��QT�^Q�J}GI��jw\�vMb[�Ö2��N�|&����4�V��@n̆I�?�9������N���(!j�("Y��Qj�5�vH�K�]��&�K4l6�I:Jn!u��-�^����O�p�&N1��%�d*�/.�3�]q��)=��u�s�I��8��M�_4 RL��Ea2΁8�
&��(o�MO�rf����Mm�>b�[(AY���l�'$��4�8�+����;3}���ɧ�w�
����/�3�M�̵ZJ�8~�ч���Q$�FH{?��C�}��*�`ddE�f�@}h��kH�S��g������CI�;y��[�.��$Ŋ���*�o���V@2[p�¯�s�d���5� ��Bob��~�tfv2���8�����u �#q^����kY�0� � �X%�_o��v�㙺�<������5I��zo��#�:X+�C��*:�#�B���n)�!z\qI�N��������Rҳ7h!���|RRp;<�3qF�`�;�Z/7����9�ipt�y{'���+�5h���=��EZO�2 3�&�ӵo�,�1�eY�|F�{�ߪ@�6����;�U�܂i}[�� ȍ:'���B��3H��mh|:�c�=�A�"20T���[���y��x`��"e�w#l9�����m=���9*�>�%�@���r[7`
0�e�ܷ}]-��Eŵ
XB�$>S���?`	^��?⸇�[姆#�\p=�Vz�V�j�	ț< �%���%����x,p��Zc� ��>mג���F)�M��y\��ߩ�x�+m��D���{f�U/����ȴ?�w�mټ�F,������+$L�dz�8�{QB�W�p6�� �qc*ut��H�0FC&���#�����9�?ێys��
en�J�C� 9��˿y'Ŏ�>��@1�N_�1]��c;��+� os��"	��K):��L�Pb]aR�w�����s��)�{��;J6��uzT��Z(���Z������2�=l� 
�C{�^F� �3�b[�B
�x�=�3����m�Nz�E3�	�a�EJ�A��cu_h��n���H5t��,��g��	������'����VES��LlL��d��G!��������	 ��C�>=Q��%,�)[�q� �p���6�t�4* ?��Q�i;nןR����P\k���
jw����ӗ�nS7ܹ��q��3	�������
e2��ծ��$�yj�p�'YsL���d6$��� �����,�)�yF/��:���"wmH��L���:@!�&�E��条�^KK�eҟgK�CLс󚟓��}�z����wb&�'ϴr0�Ŵ�
�f�sj�b�2�H��ﺟ��7��"��M��/�lj%ˢyU���qR�����m#R�O�S ��DRb]���Bd!KU}��D�5��HE�z���r��9IS��l�L�ċ��L�]X���4.ѵ�[��V�"dr���V�UO�E�5�� }�o�]�A�?�%-��&F�!���,O�g� y�:��)k�@<�)DB�Ճ��ɍb^3�jA57���54LYK߭�T2L�f;�4'���"�a/ЂD��@�س�����w:�MzqR��|��YE�xj��gEWFJq/�T1���X�k0��I����|&i..��sR���m�x�h��(���ǥ� �)�$����D$ �MWP�]H�ۡ��-�|@���-&�����R7AwޞK-a�p� �F��X7�X�!�s��WBbO��A��:ఢQ�6 �n#�J�+}
?����[�:�A�]�D�Lfv��-mor�����E����',�A��o(�T���U
�I����EyȠ(�d˶�̮�̘F[0h�g�g�^��d{j�b��ʻ�f^��V9�˯/W+�Ճ%`�Q����\_?K)�� ���{	��YG6�"�B-����8��v���%�u��g�0��k8�c<m|E�ι���Fw��S��t|���0$V����7z��_�>^���ɛ�?��돡9#4���1/�]�D�@V}w�{�m������c�d����i4���УF��ƌY�m�I�u`��I%7��pN����(BK����Fb���%��9Q�*Q24Fh��'�=`�0�����17�|W�Zs��v�U��F�P����"]������0������R[��J�T_ʹ�>��	��(� Hl6�C���Qh㌳C�U�|�:ƞk��;s{9� ��gQp���M0y~��ʣxQ���Z	ea�<��:".J>R~�C�q膅�x��y(=aeR�	�og�<_4��õ"�JGs�_c�ir�����o�(�yk���
�!5���IG�/U*D�ɢgO!ź$$(NɃFh�i|�@���G��𒱠���z�rZ;��XwB!�4χ�֭��d�M�>";|�����\FY�饔HY꽄�|/5 ��]�����b�i~��2��E
3��SW��d����W����j��r(bWW�{�U��:=�|���#%�yM_������sB��tr�R��az�;�uK*u�<X���bT�ѩ�$���H	��Sޫ�Iu>C�`��"��fHH�;�^1n�&�-)T�7�;���Y#EN�.�\�DQ�f�K�$D+�|��͝Q����,]�_�	�L���m�Q�Қ��:�Dc�iB����8@AH�Dƞ!nu v��Q)d�^H��ȭ��l>Hm�:!���i�O�Sf��ȹR�������k���adۃ� �}�I[��9�P\ǒ�c�} 2>�L5��ɹ�f�������Y75�x��>�5�+IfT�z�Y���'8+�ױr+9O)H�0~e�[��S���G�A`E���p��V�E�y�S�ϛ�`
o�,��`h�/�]�TE)
�1m4L��C���A�&��Z�]�eZ_&�B������#�2E���7��`�P�l�u^����7�r���,N]_m��7���	nw���U�Q&y�h�Vf�-��H���2���_�7�A�__�X�i�⺜0�Qy{zb6u1���9Μ;>".w����_����k$�n�)�H`��xa\P˶�J05 ���}&`��@2c��^��T� `�����L!���G5�r/��Y�J�?Wx怒1��0��؞H�=#'`�Y��ŧ��f}u��p�V��&h�M����kb3�}Qi��T?�;����H�Y���]'Ɗ����73�Z��3�J/���ҸB���;� h��eG���7R��ōqp�i�H}6֪��֋x��6�	�Y��{ַ���4�@�H�b����VӁl�N��VR�m�o����T/�fҴ�{�wJ���DkV�� �pm������^�b�f	}���&�N��r����__���C8..��6:��Ƕ��8���,�oF.�g6����mA-��P����6)���:�m���<;��(٨�8a2Z<�&���h��7��6a+��@�$@a�b$u��B+jT:�����Ғ�x�>�^ &[nvK	9���������� �z۞� ��C�>��Pak@y�"��p�I/���ji�?�*S�Yb?I��H
�B趘��\��V�a06�¥t6��qP\�(�1�9�7�5�����F��)��Qv���5���?H�;��/�؅�w��k�Ԣ��k����6�d~�7�X;����'�
���Wڏ�������?�q��!���A�x�D6��V��������%a��]�H��S�gԫs���Ǎ|$�j]���֮�}b%tV�c>.IJ�o$2\7�>z���Z���ٝ�E�b�k�$��<��w4nK�.?���P���NP�C����e�
�����A��Y>
��=|Ɗ�3i��`P�.ۊ�s�(d�`�V��
-�ty`�!�ۦKA������f�>�OPyQD`���p��^S���4vگ��7���S�ǘ�E���<<=ZJ�A���a�$=��G@@�ʿG�E�lKO���D.�:���Vo}3ԚiB�yZ��֧�#W����}V�^n�y�n6AD"Nʼ��*�Dg-�+\9q_�BJ'��ΘR���q2]����q��1y��b�����E\0��5�`b6�}�4�p�PN;:��)h���/O���%�gx�N�	+�o��b��R��u��&�4d�����
:Z�2Cj�Á�qˆ45��d#7�<�'"�����l7�|�7%��a�9�ګ\d���GJ�]�0������lآ�M%r��8��ӣ���V����Z�10�g���Q���w:S�*Ԏ%��:\���N�n���c�x�Y�K��F�����eC�_Yה$�,�OR��@�㘭��f����`�0�s���:��Nc��I��y�y�7�^��'Yh���b�c�nh����[���Wb��s����1���w�k�0_�b��ޭ�kkq"�Yñ��V�[$���Ew�cK�\|Ā�0�3ibW(���Fx��c���v��I��ܦ��2DH�k������<]�2�ͬ��q��N� ����'�7���+�kG���@*��D���ekƅ-����wU���|w�n�i:����B�&+���w�t��3�>Ō�zNc�L�[��	w�K�C� T�����i~T�,|�g��"�[F쒲�`��e��$�/����TK��C�����
ٯ2Z{� ��@�S�X�Q%�$�C���VL�K,_��㓍�AY�nyV7Ä���@y����f��a�k�;u\V.��#9�JW��X��tdEf� ���\�2���[) �Q����6<�����̝p��>?c��!�\�5�u���H+�ȳ)���p]��L3h'�	ϟ2�_�v�$w�zQ����li�F����yC�.BNۥz5��ףF-L�_6�,�o��'�
�#��o���=�İO{��N�J,`jq}�}�q2~��G��@�(���7\�9e%����Cj) ��VNKP�ad,�q�hcd�J�XW4�� ! ��
E�l̠�)�*�3ЫI/>KK	�"pa'p'�?���Z�:���Js^�
�%��#;��0�=���~�Rآo+l��_RPBJX@Q_8��z| �ǋ@߃�7�I A�R�y��t��a����@1@�?C9a��Wߠ�3�S�@�V�>�lχf_~��4o�]�#Ǵ$�e��ﭖ�����Į��Cy%�sC�	���t���_I4�
�ӂ.�mG���>LJT�+a]�����A2�/��zz���'���v��� >���A�9ǻ���6�#p��y�L;�[�Q>Z�Ï���~�:���#�%ͧjؐ���y��X u���y P<u�P֩�����}�&wvK����$�&�<�	�p���!\@����l�}��=��ZZ�u�S���'z�96A�	BlߋU�x�t�k�U�x[�$�É�����e�T�_�U3О�ʲ��!)��F�m�^�B�S����{��ω��>� �G �:��d�g��s�H���y���ݨ޶�G��m3�"��g�	�"���<+�2��9x^ȧ�<?�<Y��xq�����KS���(�,6V�o�fg����n�75�X�N$�5؇+xVj��-�P$U
���ԣ�o� ���N��w�4�p�����ř+���� �Ō�|u�%�vv�?�-�^kDKZ3?����~����+#�.��P�:�	��Q1k����)�#�~8&������!ϟytLkN��[N0�D55��05g�Z�
�Tq����[�7B�0@��r.���Wcn���L��%�*�u8�u�X�!�>K���;�)���q� ������م Л1��gF�X�74�10�"�4S�Ż��`������JSƤ��Έo�����IuJ�MWE>��;,��J�<_�'3F"Q\߶ʙc��Ƹz�Ul�_��үTK�i����v9˳k��E�:����i2��VGL��ݼQ`�1+0���[D�\��Aw�kvڪ�>T.~�(w1@��4�D`�y���	�gra9>�V3
���t��<�r�A7�������f������!����`��
�AC^߬5�Ȥ�X�z���~S1�)R����=���1ǲB�:��x���8ؖ=��2x�%��1,��B�+Z�XU@�Xj d5�f�ˢ뷹��Jk7�y�qDH��U�sΟ�:r���(�&D&����C������e��D��.q�sv�`]��Zk�'��G_/���7E!��J|)>3���"ʢ�|���ӯ�]����#Uk���}��\�h�6f�j��4MdHu��)ó���ӻ�W7ec����cfgS�/��e��"FC��a�%\�'g$����'}�`zyz"�>�NSW�2�kR~�GC�:�~Ы9�N�ojih.Q��ica��5���sC%q��Q�v���	!�<����"ɖ�������U�Q\Jj~�>��pWl[H��#���P��p�@���q�w�Mo��k��p�S��"�p�^lh��;��� $P�'E�<zPT�;�[1��g��ʮD�$}r���1��<r�|�5�޸ԉ]7-�Be>���[XI�턩䘡g���������0����v�0陭HҀ\o��&:�/��Dˡ]�"����N��|T�a�v��l<��!���������?��d4`���ڭ-��x�|{�S��5�
*�TɭB����V͆n@�LR����	:?��.?���4fV�%�n�Sx���$�OÑ����q߀��_�0w!S��9�=0�����iF;J�8˝Q� ��pW����g��]N'bB�HtW5F��S��
./�G|�R�W�[E��B!�� l.G�~WX��UHvw"���A���Y-���!�jBE��%R&��&��i���&WY�S�R�\F���������w��7	fT�YQn�X���N�'�	,�	O��,Ȃ����[(7
V��&�J�5W�zӐah�r�ݼ=l;D�N#��V�-p�t��.���L��K�Q$��\/<{�DI�l�Aɵa[�Q�N�u���0Ku���S�,�S�1�t���vę���J��A޾D@�|�ͬh��r�\�x	t���'wU��嫉���2YH�k�KH�^zC������$�A<��Xt�;�����k��g>�	hʝ��|O3���б�Fw���E5@>�<�7�E�/qߞ�� �~�7!~��̜����M�I�����)ٶ���bz���<��&}jlhB>�j<SK��{���lq���Ǧu�R�'˶�Y���0�(�S�V�zu{ȫ��N�_^4�)%��/U�>��ee���T�;l.�^L8>�P�*�L�5��ޚ�[5��(S�U��T����������Dq�� Ev.,+'R0��	;v1�~j6�EF�&`.�5��!�]���iB}��xأFN��r�JA�+����{A�����R���9�/"���R��J�o�m~37�~�[-��I��G��	фP���������̆�~T�K�6y(�SH����&�$(峟f���&�N�&S@��)��T��"�V��`�t=Rҭ��s5�A�b���o2G}�n�e��*Ǒ/r�qe���g@�o�Fq��g��S;�&$Y9����I��H���h���=�"�p� �3"\�i�޲B�Ӵ��
#�^�	� �l���-��|GT�Wkc��Ld�l���3e'\��Qz�|���7��K��Ν�<�]������!K=#ڽ���K�.��k���� ��z�L������� 7��ˡ�f혨֬J�>u8w��劯�����h�p;��Q�<�nN��z�����=p�q��.�,1���#�oH�G���s��E�s�Y�F%��}�!s�9�gM�.�H@�q���An�Z�z�p�C��;,�t����ѮhW"�obk��T�0��A��<��V�Εl�7�;>�)ַ6g�\n%���Y{x%��o��~�$��aa�K¨q����]�]�D��k���W�˕)�eJq�[}/K~�����jsJ���.�Ak� ���+��K��1�>��*y0�nD.A%��I=!ea0!�c��Q�
;H]NL�w�����6��!'�T��Գǿ�ʿ+�( ompυ}���k���J�*�;��/����e��t��E��q���@7���d�2�O��k� ��(d���p}}��bL����$<���ڽT��.ha�d/�sʋm��I�4��%a�i9(�N��5b�K��}5)W�o�oV5 �S��T�{"�|!�״�ug���ͻ!��vBl�B�=�ݢ�:D�/��-��<�k��*9�TzY�����M�2/� ����E�5nV��b�e�8 �k���%n�=�D�y�iɅ�M��s�Y1�ޔl���B�%�]������y�у"ֹ� �'���k`�ϻ1����-�M0�ٛ�Z� Uy��O�&;յ��ҵ���O1���k�i�y~O��*��E3ЧT�η��E���{!ڛ#@2�x:ΚZ�lTm����^26խ3T8>����������0�	La@��hA�(��1
�ߛA�v����"ג����3#gf��}��XS�-�Xe��>�镪6�}Q�2�Ϟ�-��h�CM��P&GO���������[j�)YWA�ʰ�r�d�(S��[yme���ź�{��`��U�N��ld?2@���it��s&G�M!�T�xF��ňo�Wxg�ŰMݰ�:i9��wNڙ�04$���nm�*Ta��%�[h�W*�'���~���{��'�f�����F�F��ح�D�)X
����V�@�c�o���g=��:C�
˅|��+��%��8=&����<�(�����J��[- 	�*Ev��eN]XLY�Ŋ��I��]]_����ߖ&"�1�.5���m�-�t��J����(�gz��w���5�E]U��,�u�t��A�ڏG[;�o�ʖ	;��� ԯ��:�=�����T��-��gE\���b�U�]S˿��^��W�q\��o�8Op_΅;�"OR 9.� s��g���?���C&9�I�������!��KDn3׸�DJ��s0)a��ebE�������#���E^�q9j3F�y_9/��hsj ]�92P)R�(����_O9`�$��H��������oO�����A��9��\[�Y��d���`s�H`��D����q���|���M\m�p��Y:S��A�v�EZ�3�GS���f�<��5�u�߼��uOځL�����	����S�q�N�4J���"�� v�
��?�Ω ��Hvz�f?���R7������Fh8>�+H�Y��]�ɩ�ŹY_��&��8�!��	ќ'Y��QD8_=�e7v��CԔC�_��H�e2�*��b�W�l]"/*
��]Ggca&�����㲭��`a�&	���9�С'������}
��&����/����G�s36����?��GR%db��*y������M��c=��)S�7Z֖�''?;�׮�z�	r�`����Q��L�C��{�%
��2`����\a���~��PP[%a�PV�fg���qW'
ږf���~�(��p#�i�E���gW5Tq��ܣ(��hġ��*f�4�s�hN����ۑ��jK�}��B��[�"d���ش1h�"��S��'�be╇��u>�Z��]޾�z�߆���*e*���D�@N���9����u�U��Aݖl�R"m��>�C��Dt~y�=�)��W�f�Q)�F>��/( ��3��g&�'&�8����=^yS���J	����7"���v���ۤ jK�P�B�y�s���x��#;k\���A`ǜ9�x�E�1��x*ePf�Ub���m�����T��<���	ݤ���ըq�D2�Y��(F�⼏��_F3m�\$���iR�3dxZm��s>��T 8����SHfgW;$�:?�Y�h$5�"������<mv�����詈Q[m��"M�U�KS��.�fT�LK�/���HH��v�	��J�w�����l��k���`����.ёz�碪=��3n-�F�QGT1�l��_��۾Nt�-X����j-#y���ï��Hq�6R�{'�e�M%5i���SQ$��''��ܿ�:a�� �\?V��:����W���V��Ʒ٪AԈ�D���.=[�SO/���EcV�M"�A{ƀņ���u�S<�芝IH�nWX~���w�5�}����D����E�e�Ǥ\w�;�!��>�K}�ܳ�N�k1�xT��]ׂ*�8;G�*"_�D��kD�Ӷ�|ꙿ� �n[\�9V���������)�Z��~���7F��1Ā�D�r������;���������eQ&��4�>����|WTn�=�����,c�%�H�ͯ ��{�Uٶ�f���X����:G��YJ���<]d"W?�D��z$Oa8i<4�?'�m��������M�#+��_�.�f��!z	5:B�����9�:���tG��o�0�,Ǜ��X���z�f����0���K�~�?՗�2�;�	>`�����9'@���N�m���t��Lb5���U>��m�{������.��i��i^���-2XA��o�ۘ�aœV��[�ԁY�`Su�W1��Ģu+ǋ\�TŪ��!���2�� 15ZP�/NO*A8{d��#���=�QpA�܌E�R��Tɯ9�̪=�ϕ߆&��`�E��Ǜ�#R|i�����G�F�ɡ�L:<},�+�0�<��v��c���'�����<�F�;2��}Jº�"g�V�}���'R�9�7��Ԟ �B-޴�9j>�0R��sYt`6C,ƚ��I&Aw���ͫ��t����n��\�)�"����7�i�%�wK�T�-z d�T��ۤ>~/D-L�ǐ�v��:t�_��Z4��3g$	د��m�J��H]G�����z��S�L�'���"�W�r��U�\�n�;KM���V���}#h������ow�7TVUl3��h��.-#'�>}!�-\@ʅ9~?�{��;U��F����ϏT���qqk�B_����e��6�\��C���f��c���3��]�����A�ㄬXw4{�nC����jX��+(�`�"�q�~r?�ΞK�ܫf���u��ь�v�u7�"�R�z��!;O����m�G$��B�V�4E�I����{�&JTF����7�[�e�Wm�#e�a6�-�g����j�$��#�os�۾���@����:�g�ݡ�2���A3�&�qp1�k���z]4�u�DO�.�{��B�N)�6��⯩�JB���x�1���5}ĹA`��X�01B��Ki:�����&>��JX.氬��[9�t���T�B�A�T��U �� ,�;��7֫=G'��Y&��Ux`��/�u�,z����Tl��q��E��P�j����|��T��>/M?����̃������@+��`]��Ap�7`�:�*��l�e�jY��Qu�Ll^��K+.c�w��wwMޢ	ڇ~dBd	�e�q���ۥ�B�oF��ɻua[��5��x-��z���f����<'RYh�e>}Ik'��٘#�@�a��XS�z!ǒ�\�\�Xz�F5�E����v�YJ�|��U_D��5�+��J�yK���,�4�>�dG��y,��M��;�͍+�
��������Iv����"b�6$ ��K����X����u���XOQ<�M<�q_���<�D5W���B"�g�L`V�sB�Șt��c�/��5�����K�Ədfi���h(����3Yh1�P4R���U��Q$��s맮�"�n��>�֚�&dd��9]ے�'��t���T��,�eTHg5٤�\E4DJUD%vW��0��R��%,,s�S.�(C&�,_V���յ
I���Q�e�jA��ѧ�-a������	�ʛ�O�*�,.pIN���J���,
�=�I������s��\N�VmW���������U�� j�]d������,���mڗ��\O-�J<n�%��O�I'����g�4�ˋH��h���q�z�ñ0&���AwJɨ0_���\�Ns�vi�D�Y��9B��x�5�v�H<��~2�3�o�1�o�z�3�U��N�f�e�W'��\ԙ�"�5a���}���B��(�j�_b�%��mgOo8,�ҁ[���pޯ�P�lT����{��n���
�Xd���ƈ?�Yo}���y�|o.�+e�9I��9黋����W�I�-<���(�Ņ	��a*�V1�q:�I_�`泛��>5n���A��vz==o������#��98k���w|�:p�	��[/h�����j7�xކ��Ԣm����H�E��g���vJ��p�7և0��S��bJ|NշP�I�2�Ƌ*�t��^��N4p�(^�czH��p�˫//���
�f�Noe�M#j#�H�D�݋#�M%�R���\�
�� A�q�0��2c�-f�3rѹ'�o����F��_�.[��>4���Qy�\����r\�3S`�W���23M6��-͖N>S�\��s�u����%vrl��0�fl�lʧTtEO�\q&�Jܧ�߫GQ}�_8�$":3MQ����<�l������F�������E�l�o`���E����Ete�n���a�����b*�C�:��x�q�Мe"�a�,�ؕ$ �3��}pF+J�W��wF�ˋ]��_�0*�B������CJ0�A�]��5��/�-x���O>����<n��e}�AG�B��9<C���]i��R��4fꫯ?Q[�O�Am�|�'�4i�?oClY��B0�O�ʥ[��`���f�A�ζ��	��
 d1y�?E��v�L����DV��M���Än��u��;:g����%H�V�-�X&��m��� e���L�7�54���z
i��h�|�v�ũ�&GB\��F����7���4�:[�n�H~F�E���� ���
֪INCD�R���śﱮ�E�n��fm�,wZ�]<9_�b��PO��CC+�N]�k�6tzbIZ�=P�qr��J��lm��[Q67%�;O$ �~]�UCX�6M�Xл��=
��(��zLR��Q &�'��{1ו��;bhV�,���+5v�]<�Ҁ+�R!��x�̫'O#����9��>Nȳ������$4SU?L���Q��"�i��Y��7F����=W�)F��^��E7����>�d���\]�g~"��\7�~��ѿ�����o[�f�M��d��k�����e�k*�Vb)�@X�
�|���T�6�ϯ-�{;���ct�T�
 �y9�`(�y�+�j���\Fbɪ,���b�Ӣ:Jd.t���!��N4r'Gy���V�|�:9K:ʜU����p�D�uԂ	�l�*��e�%G�(��� �s���2Q4'��c��k�������:@��*{WlGm�R�Hu�9U6O�RU'���<4�`�J+U���T͵�F���2�\IʻW!T:�������qw�E�2xf�o�cҽ�'�l�J��({46��Sܩ�J�-i�q�>��nZc�^�Y���W\�t��D*�qz�?���=Yzy�P��d��c9 N�U�zl����׼Ⳅ�b�QfCC��vw��,�kj6���;�M������!h@Z_�R�\��?5N�)��||? �2�W��2A]V�������ij�iʜ��bXY�֚J�i(�>�l���)`�,��kU�m�h�8��ˑ�Г�ٻ��RNu\����Ƞ�s�P���R%�'j�21�ni&R�0���M#����rLcg�K�lF�U���\���h��#_�V�o\����?���R�51D�Z��#��}b�u�ܣte�E�sՊ`��}Au��E��f{c���7A�	+����)д_FЙ���0�um��L�qA�j	H8L�0��k�3m}J\��3�=�$�0]���7\���7���0�?^\Ð��38R�5�ZC8?���y1�L�q�'M|鬿��M�H��$�ŧfs}\e&r�p9�64D�S� �gr�8����`D�^P٣�5}i�S�F�⥺:�_�V�oF`!���A�/�`J�{9a+��1�j�(��Y�AX����4�f�y��u9�vt���o���ٺ�jC"��{nYr҆�x�i�-��G�t�>���[y��>�� T���R�eT�L���`fG���A�r>'|�pZ�Q�����:�(�D��!���=q����{j-ㄫ��
FQ���)𤄭��uĵlW�.���1�=/�>�r�y�]g��5�5��ΩL����t�(ت�h8��'�d^+}�,{�i: ����Z���$/j(8��ͫ$<��R&��mK�Bo/Q�&����wt�=k������U�fl�H���B��֛�H�ƕ����sdVa����=��p4��w3E�������s�u-f��0�~\;ԛ��R�C���<]�- ��j��]٘vE�
�^��L$$rp!�P�}2�y�b�jx=��E��Y��a|e!�G+��gX�5�β��e ʦא�c�"���v���xl.f���K�5x�Ʊ�x�.QBM
�������OZ����s ?���a?DC�������.@Aj���:��7B�!��7�3dw��+*��wA��\�4�*0�,9�xj�{/ΩY����K%ڗl���.���+�������U[����W!�/�1�hEj�vTH�.��2Ki@[�����A������yu̘��&�:6\g�>��_���yj$ �MX��-9�g�5��x7I ���/�;W�&c���M�/�׭�� ��@�ֲ�8�\�h���#���:k�h�-1���E�!�B/���tgP�1ѡ���9m����,���obb�v��S[��M��g�A�ę�Q?�!;[�	f�+jgv"��+m��0�Ͳ�{{/�C����"_�dj�M�
�

�e8��[�nMc�>(>,�-n�x�%��#i�Ɍy���e2��@]pw�A�1�E�fړ�@Yz�~��GK|Q��8��� 3��?KJ��+�G:����R4�Mؠ^�<���g|N��ܩ_X�EĞ�Z7���������)�����2��2����w��� c��ƕ�Z5�i^��6h�BI��o8J�0�$�"�'Y+Vۧ`r��O��G��+@�A���������:�j[����Lvm����
U�����hw )�`HZ����0����|���53ҍ9�0�ĝ�\5@�ݶe��� *�q�e�kc�p���d��!�Aa��>ρ��w�2<-�u�e��0��������f�rF��ؤ�D�6��~e��:M�m���3�A�ar�Qn�$-	��I�ʘ����8��~Q2��	�M����n�L�̽��(���F�ٽ�v���^P_���ۆ��s�lN��w��e8(ZCB��i�F@���^,�0�@�Ն��ًxhB*�s���5<������c9p
���y�^{I�+G���$_������Uq���50@>�{Bz
�gı��BPmF�]���o7Ĳ.a�o#0q��u���^��}��f%���Sb�Y�W;;[e2&��)�C�8w&� )o�
�K�R�������j? Y�S��=P���-���2ߡ� PU� 9,Ť8��yNSj,���r�.I�m�<��Z��X�����.�m�fWjGy9����Lť{����b��/�F�Kk��HHq�J��b[�9x�Ѳ��W�!S���~|��8��v���aƐ<,�����Չ+Z酟=l+<����j�PA�1Z�x�J����0����_G��E�q��dg�15����)�t����#Wy���fS��Go*���g9�Q�(�\85����a����ȼfk���cn����?������A��&y:e��Vh��>~��;�*=�+�c_�v�γ��{ Iy���
r���J��ǝ�s�IF���M$W�7@�Y�=�*�w��Tc&SD�s<���mYj��"|NB��C��i�(�E�ѩ�RI�V����'�ן��3"5�Ēe�!�${�;j@[�F��C�C��t�3 z�����[6�:Ύա�=�ݻ�����]��eifpIi>W���w`7/��=���[�ܱ4�Q���X���tf��w�F��{�!$_o1��-B2m���X�=�׿0���ا!�-��P�C����ъ�ĳD**���y䘆�!3��y\RgiBi����^�b�-�\S�W���W�_u�q��j�yi��e�������0�sY���r0�U�f����ghmV�*��^R j�[�F�D�����
���T��ɖ����F���~VHQ�'����V�gݲ�`�m��\�|�
�n<AWR��ךHp��j�r��gC��{���b_���<������I��J'���>%�� <�(���lxz^ʔ�Tš	��	v���(�R���鶼���*b͑��;�C�/��d�l_ѵ�Ց��1�3�q
�@z�͝���	j`R���0ÏM>���O�KIʳ�@B;vhnO8��jʈŖ�层�&�R�6����t%�����M�������W�ǰ�}�
�<��e^f],�(UϭML�|뱶P̡�6�xm:*#�Tv��h�߱*�@�Kgḵ 9��?�aY,*)��vn��Ic�����x�RU��X���}���lB�J��:�KR=�t��y�UT���v�d���f���*�GT-�^���T(�@�5�J��L)2�ʮn����?�z8��j�vƍڨp�f ��T����I�M�;oT��{}���E�,c�vͳ�$-s�x���X1���xKf���O
�7?����/P��v��5+:�ـ�PY�g�1�s��H�
�t�d��Aw��X�E�q��O���E١B���Z�i󵋺�Lr�a'\��^��y*sTЄ2~���h^o,B][FG�CuL ɤ���Q{�E=C�z���ּ�;�!�O!��/��K��aydC�4�/�U17��eőN�;�6�3�.���p)�#2���cGJ��� �ٶTJ�^G�Ӣ�ι���,�)�5(���
m
D�J�
����1�C�cڵ���4f�좵P`��v�iu�i��삓ʹ�N �k��RM�7���8����F�I�lak�w�<A��BW�������2;�{\�p��ƲWp�Ah��>�KA7d'���0���v���a�ϣ�<�3�e���<R?TE�+�/��R�[h�#�g�ʾ�r_P#Y5.P� 6�L b�s�E���I|�ܭ!ռ��g���ST,k�/�ώ���l;EaR�h�S��8?�2Ӗǐ�BUrI�{��ǬZH1s��cW�c�"�F�|q=�� ���e�A��QV��^A|�N�X��J���ow��U<��L(zw�U}�g�qB�	��n�G��ꕓ�,$�"(:.9����\��:~�5O����r���#x�F��;�S �h�`r�{�@�?�]��,����=�`Di}�9K���lT���.zZ�̈B���S�������r
R6U2-��;��sf
a}��Q���6��΅�ƥ�n��q}w��6`��%P�*��_��Z몴˺j�^C8
X*�f��٠��a��W�!��گD��w#3����"Z�Yn���i��y+A�A�c���TT��K5613!g�Q���f'�gS�jS���Y��Egz�I6�����	Џ����1RS�5�.s,��QӠ�v�$ͣ[
W}m2�[6�eiq�E|������f�E>�u�~xbky[y�RZۉ9)��/��ι��+�wq�"��"��[������j�	8�:U�����$�1�-:���.�����D �Z����&=�%����j�|=>��z����e�p�Q�w>��D�~/0�:���Δ}��h�N���<L��>+)���Z�������^����CC�M�jo���њ"M�,H���~��|8hzz�����TA�ulb�M�n]�4g��/��
�с_���[�~���7�yd��x
<k����r.��}!lQ� d�5*ʄ�@�P���e�|h	jF�2~�����Tx�90��]Z0B�\��9��A�FV^�<��h��^��-d�@��E�,���qN CZQ�UU��:�O��pl��W�m� ��7�س��ඐ��/�:`�ü�!3�:�k ���GV�9�!i^M�F�3e�b�}������: ��|���JE9a&w�2����h&�0m\��h`�lș�rՍ�9���Q�����C/��+cE���/�2NX�$����2F���G.r�{!�E�Z�p�A?��H(�o�$r9N���K)�ɻ�]I߸�)�k���go~��_�*hx� Pd=E�3�Iaqv��K}Y-�&THW<��n܌2�eU����}�Q7H���w1q�<�q�3�*dNB.H��_�9lW5SERs�?���]�<�b��媁���a�+{ꗕ�W�P���j������Ǡm�A%��P�sa�h���4�q�Xg7�.����4��2���.�^Ts���	�u�{��F�.��a��F-e��[�������"lsw>؍��w��^2Y&���_���^�R�ڼ w�[������)�(N��3��l%�Qٸ��y�!�>��+U}��J��A� �n,H&��#�e�P�����`ֳQ���'�uW��~7��,
�o��%����V�m]���m�ُw��|[W�&0��!�~&�I	^
��[�H�JD#m�B�/d�$:	n*��Wra�"��r�&KV��p�i#�)6��X��.�!S�������j��̀V�x�Z.�H�'RM��F�N�n�b�'s�n��5��r�}��uB�q��yÞ^�n�*:���Kh+s�U&S��#p�:љ ������_��5:������ ��ty}��R��	?D�j��l��W͐NA4�������R��k��Jt�R���=u�r����}���O$���5�=��~�b�Gu4`�T&^�lπ�{X{����{u#���L��s���G\�j�9�#�<B[;�\�%.��Rm�UC-��ޖ<9�X�+�q ��rF��2Ä�$V�7���2�CU�ͽ�['2wS_F~R���F��3�yꀔ�'�1�MY�k����s	�zv��C�� $[�V�f�����g�G>a��/+i�P���#���P�n���?�[�ӡ咉D8���տ�A�2o�^�r�$�I�ɯ?h��w��G=g��6�L	��:6=Ze�Z�2+W� ����Ů�X,��6��h��͂��x)�u6�Y�j\ꎚ��}9����R�uׯ/e,?V��3����?t�{�1#qi�?k n$OH{Չ��O	���,>����1r�S�7��� E�4m���C[�S+�b,��0]s�J�_�3����/�}��4{�ހ��.���n3?�`�}�-7��M�A~�d@*��
g����.ގ�~-Dt��GSˇ����ˇ(mb[Z.��{�F��M�H�3�Ë���T��Pe�M�Ɖ�g�S��Ab}�A��_���"K6�w����"O�v��7U3�D�8�D��H���E|���y/ZW�{�}���ۢ/\�{P�bE/�|�:�2�Tl	íӮ�[� eM؇�ۄ�-r	�X*2ʯYK�|	����bV3��y�������E~���g��6w��$F����UXM:#Xv�9��GM8?���	��摰����:�O�>e�?����/�H�o���2٠���s����J)=T�Vv@�ꊿ��-�:M��v��D�V�H�ڥ�v����RwK�4�����
��zD6��wi�\�b��*�V8E�G��0"A�����4kRE�G��6���uv=�q��\5�5�*K�	��Q�2J�*p�tVE18ZM��z	{EϢp[&�-��4�\	��,�H�I��+��X�l0�y��כN�q.Z���D�	^���I�r�R�~ �Yr�:�����X�������:|�3�p�u~���g^Ac?�t>��eZ�߃V�+�	������M���	�a����p���(惡ۀ�0λ��:56��f:��/�4Ħ���m6^�,Y3�a|-�n���o_��uѰ�Q�.da��D8��7��v�E�q�W�҉E@�~�Ƹ
S�G�b�d�Yٕ뷠-�DF� ���/-��[u�s��!'��t�+5�*���D����u"w�aA���D�B7��碒/��rU���S0�t�k)���d����X��F4�-�}y�?R�v@"�(�Nr����cG�s��`�:�e�0,����&��k��~��<�E�Yn��|o��set��
j�y嚘z�0{7��/�E,m�G~)��ǈ���%F�\���}bY��H�(�v��fا!&T~�������!���o<4Fl?�:ޗ,���A$��q��i��]N|<��R	&�?��ϒkH��C�B=}m��`5��x��(�f�O�lzw�^�0Ĕ^�����2pf�	p*�v��-Ȉ|C/�F��pԳg,)�k�H��/H�؝N4w��C�% 5\k1p^C�vvͰU%���`*��=���E|\1!��#��e��?�fW8��Qo�
1�8������ĳ�9#�C��`�y��H�P��y�Ifb)�h�Q�MO�r�t��=Wt��9�I�#�LFogWee��y��������l��3QЏC�FY��b�Q�*b ��y��/�ьR�9��'��A g�j�k�<��w�e�!�?Da���~U���郊9Y���LC�&�W8K���
{�*V�����Q&q��}U��׻��AG��C(� ~�w�\���4�z�[o��/S�u�şFr���nD�!T���u��z�+��3�6� r�7�xhf�2d�\2D��o��F�?إ��n��8�R�S�|35�2��x�2�B�RDBn��������Bq>̚�- E}2�n��h�������kY�;�T��wx��S�@XkCX����Ǫ����gȼ)TC�Eޣ����n�?�i�|��6bÀ��lӁ,����Bs0�I^Tg���g`����3(��|��<R����ş�;��*u�N��k�+��^n��+��m�e�U���k32f�Bq�=�ֲEj�v�;>����	�vyt$AY��������th+�i��{1�j�4�7VT�����-�{n����
��ٓ��a�b�}`PE20_�bD��n�=�8o�7�Ra����F z�ADv����������K
����Cu
�XF�����o�z��6_� �����|��-	��혭P�� �Cz�!7N
�C-���l�_2ڛ$[0a��}��$aLS��^(��G�~{qd&k�k��U����f�&ƞ��!2dMz6�r�}y̮z$f��hT���Ӑ�6 �}���_��H�}a1�h*L4D�X�r�Bf��W�`��"�\ڽ�D�I�	\�5�B�|�3G��	�C<��9׃���Lbhh�|c��v��~}�L|�G��w�����݆O����]��a�B��i��(%�˦|�|���`S"�N�7�%�<�����Z;~gVs��g�jQ�Oa�����`T4'K�w:,�Z�¥��p$NY#Ő�ZV
����X�����n����f���)s���^�_<��s���������a����Tm&�.E!Ҕ���Fÿ�����)�S�U��:E{J.��.yc���P�t�+������El�!��@��[Zꋑ�ZfC����u��-rxas�O���Z���"i�����Y����J����<�U���aֆ4|X��u��,+�-�c��3NxR*�X�5e�$M��®(�j�����ն���M'#D�9��ul��g�7�
�g}bV����z<������P0��Zry�d���O��#�|�'de(Fhc�1_�u�M�f�F������m�Lw���y����@��������f'@\��ލ�u۔�$~�r=5��r�XG:�,}I
��m;C�䌨�$�å�E�[�h�yg��r�i3%���_q���d���f�pR"�$�v�,��vs:4#�-3<���a��[ß��(+�ñ��nh0Y���+6U�M��X[�ga�/۞1=n�����.90��@/ 5,�E�>����ɗ�j{���H$V�:��V\n��5M*ǯv��;Ȇ(�p�{_���&*ˌdP�M_5���<#X��+�J�x@3|�ZHk���$ VaU�v�����Tp���8	R��q��Ϲx3��ji;ظ�Y6Nilݷ���4�!ݠ �#uxdQDž����P~^A�2���~M�\���2gսp�y�����
�(������;slsǀ&�}(��qI_"��B���8�[ S�:܅t�vVW�ǉ�K>\���-X�!�ߔ���۾ΗP���za��y���Aq�l���@���F������!���h����ԇ��Mn�ɥ�~7��"�����OX'nS�*k;өj��,�WR\as�L�EK�b^̝D;(�IhDu�"6[u3]�Bi[���LJ�z�Q��[�eӉ!to�)�Ҵ�7���\�?q9��!�F�	p�Fy�ܨ���9G�B�ل��'��z�ʕ!�6��.?׼ �ffH0A���Й?�km �,�6^:< Җ���=a����c1��,��_�I���R�H=#���-k �ÙO �G��	s��U.r:k�h�8m���9����Jd�T@y�&�QQW�CR��[����W�fjYl;�0ϱ�PX�L���U1E8�%0tk��8a�+H���������#�VHiN�*<�`N(q*1�av���j7C�YLC�4��b����9x�z����I�/U���kI4�P\.Sv���H�d�{��p���w}�3�t�t�@dK�-=F��Gܙ��s���%�((RH)2;�;/ĥ����x"@JY��D�x~n�{�e�B|��� űb�"��hN�Mr�A����;b;�,.��֩�)���2��o�ȸ�1�3�Cv�[в y1�H�8D55���	���h�wsR�� h�+;�,��4�AaR3�����b�,��F��:��B��u��<�����&-��0�A�˻�ݐ��.N�����N��c������~no�S�����i��p�k�`�r�NS4��EA��y�)��^�e�9��iQ)�(��W��I�	fNR|�� �[;�צ[J%��6��E4ڪM�r�0������� ����NJ�ov e��y�p�����kW8��Y���2Ϛ�� ���8�)���|�#z]��aͤr�%���$�+3�!�4΍�-r���*Q(�������b��f���W�������rXj:�ӑ��/��µ	�,���R�|苓0�����?�Cbv?.��������dzl����c��.�ić8S�z�/F|��b��K*�����s+��i�<N��dS�F���hNVIA�$b��L/		���Y�G�08YEE���̕ A 1j�s���J���֯�ܙ�Ƭە��f��뇷#їĊC��7�]ճT�J�ɘ[RS���-��|��%��JNgK����3ʉcq`Ǖ]����9��3�_7q���q�,ޣ�{�2_)IH�2K��=I��Ա��rv?#�C5������uJ������Ǥ��C��c~�Dl�Z��4�ÉP4� dE�� �<_�����tW.�p��b���o5T5\gj9�m	�Gg����_ X��.@v6Uj��9��0�m#.9P����H�D
ϐ�4��[��D���=��"������;��ҽx�{a]rq�H=3�̒���=�X /����j�U�i�EV��(,�ӹj � �c���sB��R���Ƞ�;@FV�J�@��v���θ^�d5��tE1e�������}P�D���^��A}Q������W���z�A-���L���� H�y4瘳�['?Gʠ�h9��{�"����{����(���W�7	��C.?�]���Sj��e7��|��x�m�����OR0�Ǔ@����,y~�PZ!@�lZ�
��S�v�0wu�Dd�B޲'<���8�`d8^ZP��E�x2P>�=������x�!=�� \dړ��*j�L���nU:F1I6(BB�eR�=h�����::6��ԦZ��e��O�5d�-�y9� ���لbP��� tO����S�NPbd.��i	J� VH��C�\3�Y	{�eZA�L{�d�=K]{ �NE%M�K��0OPV��nh�E�J~m@�%�ǋ=���M�R�ae[�S- �o���Hq]¨�&�ڝ�6���熶v0�<�)CaK����\�v|Y���Ft}L{t���Ώ%.ڋ�ϕ�����H� �����cEI-F5<��E���s���C_�u81�P�d���-Pw��(�֭��L�ܘM�hӭp�'�U��C��;����uK�:�O������ޥ�����%�4~�L���JR����� yPׇf��J�S<��=�;�O�����:�itu�W���q��٦�Ejh0�f�vY�d@��'l��
�T�i���Ǎ�ϼ�`#�h].H��3�E�c�_���ҢS��QFqtʵ�ff �1�=�<&��C(2���L�&_����
u���A�=p��)
�3��(��eb$O��U������g��ה�/")3|V�P`���3�Uݠ�����0��^$I��N$g:.��P	;��$�D�"�QPT�=�S��� rnv�5(�V�h}d�ㄠ��]�2D�j?D�[T�G�y�@n_ń�B���5䡽�h ���S�S�z�iB>C�� ��X�(�7��ug��iL{>��Nre���)��������	e���F�e��")�"�+2�l�����]�L�0��L8X��I����<�,�@m��n�}�R�G$�Ҷ�5�Ji#�"�7BSTHJ�>y|������-�8�'��"����D����
F���H�aÔ�M>������v�_��� �b%�Ò,O�7#5b�ǰ]�#�:)�4����F �Iw��6쇃�����ә��Sm�i��:���@e�/b��ħ�̦�k/*蹪eW�.�C��y�k� ~ -�U'�;�]у�"bZ����ݙ8��c	��"iV�6�g3�aw^��#1 -{Q�[�j�jx���(*�Ç��Q��?"l�W;�J*����1��/�d���`��� ��6HOA�wu>k��&��iBOJ�$?���ģjg�	[��,���c 5kNW���p���ëg���>���M��W%ů�?��_�ږ�#�?������R���(H�JV����������U�LțiѾ7��� �3zyM�C�~� ��J�0��`3�:((&�"���2� ������m`��������M��<�j���PfZc(�9b�ѕ}�O��̉�x�`�ϒuؗi72N�wj1U�ґ�3y��ak*�s�uq���yX�\�v@:d�ɝ�=�qz��偌E��'�Z�
e��������He@#����̿.�_ V�zTNH�tM2���I.�3lb�j~]!�����)�l|��V%" �ƥe�t$ޑä1�4���f��%w�,�(M/�}b����(Ȟd#W��D��2@�oB7�1���e����<�s��5D��H�5|Gs+��A�L.'��4��/�D��U�#��<�k$vxXi��֠p�ߖdӸ'�4�k2���Z�j�5�uD!έ{�N�!$�. XJ�ݨ(�����U�#�|X�  ��(��'�+�`k.��w�����$���z�t�Aw�p��td�:�L?d�mU�Λ�n@��'r>#9$i��I��T�� �'K��!HH�X�o 0���
��v�.v��K�
�Xs%7%<�ۘ�/�{�Z#|�K l��!AP��q���q�E��Cf�&�XR��nܚU=�Wm�Y�o/���Ni�|ȗs7�O=��؃��Cn�<����.BKiR���YP^�
F*ي����E3����%���q�c/���9S��H ����K�o!�ͼ���'��(Ű��,~OR���o�.���R
��z~*c�d����0�i�ݎQ����C�э���H�<a�F�0�`p����,�IL �1�&��Ƴ�[I@���0!C e:�:d-��*�em����V�Pu�V�{��+�h�+jQF�^�cU���m��,%"���>�K\Ee6]�=v�#$��3<:��$q��)'*z��Qu�O��hH�����;���Bp甝9�)�4�n�����IƖ�j\��x��S�n��ud]�r�1�d�%)@�kXK^l�Ԑ���m�e�ۧ:������ A��e���fwi��5@�ԁ-���JSf�Q��4�D�Ԟ*�)�H��؟w��+��������/���g����q�?Dm4;w��v�6wIa�#��C�[5A���	Z�K�^��d��ݟw�MqJ������&_OA��	�������c��\s|/�_�A���:7�1��\J�T��x�+��	>�7Z&TWέ���4;B�����UM�|k@. ]1���ۯl�NX��N8X�?�ӛ�۹�5����������#TB$��~�
�`��?o
��
���bq��,���������ʽbn�k����L*f�����aC��]I'�B���o��5M`�FЪ��4����Z��/���ҊyQ��Lg[Qᝐ-�y�?�nqT�&6È*|���1:M6�
=��%�7�V�9�)�����*������Y���b��4�.e¢K���e��c��tn�,~��G��s�%�
�y������ �YWk�Nhwo�o�����e6�k�#�D��@��I"�š��kɣ��.�[�R�{*�K�l��>�d~�o����Ykg��-����@��'L��L�T�D����g�S1;���&�����+b����4���'�a���Xi��VU|�TJ�%t�~T��)������P5[�{��ۣ5oE#��c��|�nH���t�⌚9g�S!�� 
�ja��R6�Ŧ����w�]��ښI5��Z�FUb��_EdóN
�\M}K�-M��@�3�J�#��0wX�_ܑj��q�AS��<���6 �(���]%h�G Nkoev����%�{��KJ�@ҿO��9"��26�~�b�%},�B<>	y\?N-� ?=���V�sAݓX48��R1�8R�{ޓ{���z�]��3\��1��-�[�!�|����>�RO��
Ï3��3�L�NM���T���l��^�tG���훈�lʜ�D��w[j�D"�R��s/�M݋x�o�]�$���ޣAbM���j\R~=�� ���:�c8ƺH�k� �y&XN{����]z<�<G�ے4�x�Dp�(��9(�������c���'
Z�
�a2��ӂPdG��<){��-��#,�n�[�����H���"�@Cv�޾����U�
Q�V_�z�y?�ChM@�5&����"�;+�m���)"C�����w<1����RA�ڱvl�����u3�r(�pt����F�r�=��ӭF�1�Q�mx%�D�+rzG$�Ļ�}6d�ɾ}4<QT�R<U�Yz̈́$��RjCMF�9wP��]�d�����J�e����a�o� �HT����R6{a��?31VΛ��c��yI�"�Cm�'�g,�:�����j]�ְ&a;��)�a�R��.8@�[2��@;�x剔ta�TRbq��-Br���i�CL�����L�(7�B��~�]��WŴ?�#���� ��!�&�i��޳-���D�'s���Ţf1�@#$X�1]tb���u���w4w,@��)�iQl�v�2W��qe(�qR��C+�ߦ'�8{ ("�A%Ȅ��j8�p��`ƌS���XL���w�t�F���v0�:qL���r��N�\۵$��2YpGZ�)�|��h�X�>����͆��%����{�[g��(H,��d0|$`>����ε-2Y�pkI�|�Ҟ9��!AK:w:�I��>Q�e���G1�']Ё�l��i|&���sgXhЏ����B��8�Ej�-_^�	�>DŬ�.������*7b��H�0�eu����ܚg���(�*�S��?�ͪ{�zA
YH�}�W���>�gm�CtL�yT��Xh�y���>�CO�T}��}j�4���(����!���W�~�9�k~�۔�����5|��vH�[�%�B<{&���������^�͛V,�77YC�B���d4o��P��n8�^�3��6�k��՝ ��'�9�~f�-�]"��<���U�Bj�bQ:���;�>�6y�|m,�:��[G����\AqG���]�_H�c�<T{����X.�t>���<{�2 �-����a*}��Xր�7ppq�����|�s(	z%��%��w@[R�5_1�#V+=]m���b�6�R���r�l(���G�jU	�7Gd���#��>@f�/s[�t�˶Z,�\ֆ�����U q�}�G�X���R��d���@7�����v�����_y݌�o�b���WXp��1Mj`��U��1���+g�Q��Zx��WdkՖc�����N����U$t4K3�K����^��=K�E�*����sG�k�O/�]���yY�gR�]wnk��hL[ԇ�ds��^si�h+w;�d9�W<\��u�L�=��e?���m(:#&"�DO��oL��� �`�q�'�T�tQ*��bS!�������hs�ߋ�"_�P�eF�cJ2 @Z�;��܆@��2����ꁉ�A%	
�m���8����:�	R;#i@0n��h 
j�$2��o6G�sҳjf⫙e]�����Y���>�H�H�;(8	Y�xB&�i��|	��!W����H���0�Q�r\7����fw��]B��V3e2xߥꕹc�=��ں��[�a����߳�/��_T��9˶�Hh2��a����+ƃ-����g���ב��gu|-%v�?g����m���^�bcbdRt;�P"�2T���Z������S5�@��h�!�`J�V��A�x���P9��5�&�X�^u/p�p|�v1�N�˚�д��&��g��w*L���}����o�M&�3u���u���1�y_0��Ϊ�r�S^�^!���ç���Bi$i��A��M������̲h��>�M�9>fʛ`WZ���>��A�6!�c��!B�йם�N���T�����:C��ps�t�����.us��]<��T��G{U`Ņ��Y�cަ���u�k�
T�+'���+��RM��K8 [P*��2�M���BP�G�_����R���G����Uc3�$%�g��C����Z��@]c�Ke�m���ݸSx���Mpc��%ԁ<�C��*_/y]��UA�y�+*T-�Q��a���t�J)7"\������JT�&������$Z��F��ld�9'��d_�@�~�F�] �֫�pe͕�<j�J�z������'eb�'��5�OƆ����j�e
�چӽ;L�H���@�0��׸+�l��(�r�|߽9��Ո�E��wJ��8�q���q]�3�����	Y�	Sϥz)xm��=�)�N�JZ��]�ɖ#��N��Q��=�[���ർ���N��Y����!H��R(�������s�C{�%x����8N���U:�l����w�T�,@�ٸ��D�y��
�IF�>�rh������;�~+�<�k����O�fy'{�A�PjN�W��ۊ���
�(!�ާ�B�@䍩rv�냄_����g�$(/ G�7�U35��g0����=�%�؍L#)L6b���;�3