��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�i��a
Α1S%� �uj?�L�3��TLei-3^5]E�$���,�;�^��\fǈ,㥜��!#���`��^%�؎L�>�b5�1�c��+}�����S�ձ�8|�0 ����sc� ��h�p��e;b� Q�EQ�t��/Q#�'0�����V�r�F|��?�kH�썓읽E�nN��oh�RÓS���Ŧ��3n[�t<+�`�[Y}��$fnmM~ɕ�?p��U��M`$a�I������x;<A7?�Ee�)����ۏۧ|"��=�~͕��>�n�<���K;b��?��p7�R@꼶�xY�зߪ��"�+��AC&����<�	\8z̾�����9�t@�t��.�S�ـ��Y�L�kx���y����= �ҷB.uB҉� B�ʉn3}��8���L����H����Vx����Y��4��Pj8��i��~���%R%7�_f�68ص���ӺonXj��2��19�Ci6Q��7�J�Ҥ�$e,�Un�*���Y�t��%�����Z$",�Ы� ��!q�&�"#,�<	Z���q�y,���߿��o�5
�0��e;�/;;|�(`Qc�g�g���eį��a&e� y�����]8|�)�mɯd��������W�^�5ϑm��){���?ޅ�k�aіQ�R���s:�'aH	��:9�넔h���5�~#�5`E�,ؐ��6�l�0�g
O0�,�������͓O-�* y)�[�(E?�j��l͛��+1򺦍�4!i(_�+��|�pL��SMD�(2�qy���/�N�����R7.������MO��&�7Y�����S/��!����s%쿰�yo�R��F�,����mDƨ2 �>�E+ҙ�寤��%��X�f�N�dK0���B�0=67�d:��<�#��C*�?^2X��+��n���1/|O���u� I)h����u ��[OSa�I��mu�Q��p��2���9�.��^�l���]�'��k�ſ�����=��g�g~�!O�'�=�p�Y`���C����4�)Vқ�bg��Qa@�c����:e!N0>�-9��A'� �&Fէ��U�D �	E�g��E�?�� 7S�����޽NCT�w ]�%Ϫ>��^ZD"`a�}�a�}u<�����e'v_x̆�cf%�#���(��������q�J(���
���sf6i����t�͠����ZP[s
J��up&���JÓXukcI�]
"�7��hŅ�����v��س���sXǹ�k���G�����.͂����b6k�x3�?S�Z@��X���ʇ�9A��C`��3;!L|I����z$f��z�u��4W�H�U��0(�VoZͳ$�㙣ۤ���k v}�B�Yl�;�b���vh����j4g,����c�8�Y�W���C7�KI7MK�\kA1j��������� Eo����iۣ2���N�J �*������t���c��>05��0�x�	��>;w<�F!Y�%�Bw�0�t��:�[�4��%xK��`Ui����]�[N1���mX�$�����>f&��(9�}��z�z������a�c^�ڱ��Z�q��O6ٱ���б�q2�D�c�y�����)�BuZ�9g�?�mǍ\z0+�}D^/3��`���Un ���N*�V�L�ʔ�
�|��g�Z���
��(��0��п�m�&f�7]����%�2�Н�]=�gb�P����I��E��gV�t%���Z�9l�x�"�)"���u�R��w;���7���ir�U�7_�g������lR_ǌ@���MJŒ�f�(��Lӟe2+*[��+{��1m��#�t�C��~���sq�&�~��׍M]�{	%LL��V�T�tyX˶�]:�4K�P�}b�̝h���GR]����e������r6�0�ޜ+� �Je�N�j�;�'#{*���9���dݬl`P�: ����c����������?�]6�gծ��H�I��K��.!֦![�=q��� ��YG-���t[��<̲W�2<�k{���Ox5��L��W��i��E���iv{��#{uݧ��~�c9�oP3�l��pSi1�7��?x.6�X���C1tߕ� h�&��Ԭ���z����u�;��ES�J[�ʳ+`��σ���)ɉ�	�g(��q��Dܸ݀1��v�i
�w%�Ƴ�����$������!�e
��0��IöO���v��hE�ktSӆ�0����GόK��|�,����_?׎)-ul[|�����w*�f�V�!���#�_$�M]���_��NYL��������#��މ�8��s�FF�(��}�??-
l�t����_[���mn&����m�K¾l_����3��FMK{uŐ�Q)�B�ʵ�x�CWE���(���g).�H�jI�����z���9^��F%�P������ZQ4�l��PGYihх���g�Z��c�
��oT���}�4~;z=�����\�mqYe&+�"�=]8f�`���NK0d��,
͔�N$Ln�gr7��.N9e+�.%��R��lJ��<��:��H�7LUJ~��K�F��'�.���hތ�+IP�]��%�w���C���Jp�AH��i\KDuFkH�+�"��)d�Ld�n��)�jzg���\�v��w՛:,�LBF�kdO���#�O��5ò�C�WC�F�Q���\���ԑ�����Y}jڌ �.<Ǳ�XL���;�꼝C>�dC��%M� l&�}Y���_�Ʃ��|�����q��"� ��h	*�
�30���W�Z�5.�g�9u&�1{<~@�]�%���d\PO�:���]��w���Y^(5���3h�����>xc��I$����[�����V�;8�/�d��23FrL�R�Ū�إ�,���,	±{Ö�����D�^b�]y��D�M���ųP���ѕ� ��v�Ί�,$��bv�%}��w�a�ir�#�g_��'�J��O�ꪙI�4��h��}��D�N2���/`-t�dV�@��!��:{�]�����2^}�ΦM�RU���B�#��FR|��_6�&δ��}<��zP+1pE�z��h�x`e�v'�昶<�C[v�m�E�̪wc#z�;2MLpy�8����j�%֣��!��_3{T>���ع�S��OL��*4��.t�������ҙ�:�',�����Ή/
�����5�1�Ďn[�3�:;Q�߫\�����I�$Tj��K9kⰴ:e\�����R�XI	�	������(�!���QO��	H��gZ�~�V cD�Hv��_��S�p̍ەPw�98�`^%�݂��~�'tʨ&��n�I�B�{������s��&`"&c7�>'�&���"F3αQ�Rz߂B�X���_����i�y��PV�^2����R��/�դ�
�*&!_�'���(���i>ؕ������	=���ș�l_˫����� 1�i�b�P�(�Kk#
���(MԐgP� ���Z�����S�˦�E�&+ڎA�����}X+�Kް�QWf�1Q�m'�׏ �_�chM�cx���(�}L[��2���ds�w�>��rvS��[�W��c�{���(T�i�]N�m�$�>���]����bY`u�Obd�������9c�6K�3{��ٮO��)��)�ڣ���i���hg��+� ���̓��܌�0�qY���8K�Д?�	&�ګ���O�&�I��YȀ�a�YY�J'D�xFʒ�R��@#����p���
9�؃��b���$L_�{Jm��#��+!�'L�Z) ��p��E��Ĕ�O�N2��Yj1�T/㗽=�[�����:��bQ}��!��2v����_���锑�.D6���Z��{�T�q13�y�DDw��4V^s�dm�#��OjzC�CH������E����OA��w� �НWm�i�"x����1��Ԟ�[�CA�����8�(%�!8l/.�i�� �DgNNs���
�&�
�[��+�BR3(%Ԃ�QU��f	��JR���9tTG�}�RO��2vk~�etv!B\4����ā�Hg�j���K~�Ew��� �Rzt���֫2?3D<�d��}6��_���c���)��6k��>�<E�d���ܴ>@཰��y�a�p����A"Q�����Vt6=�!9��N��ǜhC��ݑ�8�\�Ϳ�bl��MC�a�JP��xv�À� ��B��U���j4s�BN8	���?ś�#{o�.o<�Ї�^�.���;0�u���z����]��2�E&p��"R�r�/lD��ޮ2?cq[�u<��۷մ��w_��CG؜(P7(^h^��uc���
���#��Q�wz7����?�˖Gt��$n"Ҕ�\��CM=t z�jq4L�@���S��_+����v�@�p�Q�6*XZ����;Xb�:�@̛�,��lg|�wY�{���	y�'��'�� P�^x�he�2&z��x>�?l*ӚL8Z��\��?y@��Z�6�@���kb;�d@"d��	k��{2�z�%&{~X��"Wm�u,u�:[5�?R���a�F�v��M9(S�����*��#^�~J���|�7薩2md3k�3%J��Rc�_������Uފ*)u�qEyB��C� ����QB+�<�A��g� �X�	�[a��B�Y1�s�)�L�.��o���#�U�OPes��O�柃} ��p�A�%���X9��$wd�m�1��:�F5���"`0a5#C�E/�yQ�=�`�g<U��F�����n�$�;�"�>nϊ�6�kB���%C����ԕ��\\
O��P��Q
�$۲E�E>���?ӸT�(�u��R#�=�����r��M  TP����x.�IR�<K�K�v%5IR����D���J�0T���I�Z��3�"=?<3W�����;�z��ꀁ��KI��J�.İ��2�>��*\H�֫�Mn��>{�Iج�D�+�J)s��"5��j�(e@^��QS[P�6+���n�ݖc�9E����J2.�����Ry��<K��#�N�f?�`�t�a�b~�i>�� �w�MUc,(�eKq��i!�3��	[?��Rg\�]���M,Ka\����[��s��B��j��i~��u��MS�cdK��Tf^L_8ߧ�ۆӱYn�uP���)ھP
Ǧ�M�3ϼY`B.�.��7ǘ���8������d�iPl��ݩD�L<�<��5fѽ�ȕ��	&Mv�.1w(����[�ǒYf �gʌ�Vlh�+����e<��8YdH�_�<3S������X��
 �u�oj�]e�(c�C��ӃO�h�~{��^U�p���c[����}~�UOvO}���{�BT6��L�j��Eo� ���$�F���w���D&��P:�5�5�������!3u��@�fP�{��֡�n&Ǟ��lݖ���������t�3�17����� @����2�mb����z�/Pc\)��3plX!Eg/�G3���O��<AZ�S���N�*RM�2JרH���s�mti��)j�<��>Ғ���[��f�Ş¥�jf҉���>{��7n�E�V�Gx��>B�����E��Ɗ�$�9:�ޓ���@�2N"�#���P��fiV+�X��v�&�?��\Ԣ��C�7�~�}�qdh%��͈m	����oV�9��[?�-���f��/�T)Q�s�vEu�5�ěaO�.$l�{��[җ%���p@2) L�I{L���{pD.E�'3%r�� k��W��Ktc�
�톟���ځ`~py�;f�t�뾝�ނ�9U�&����r����5Lq����f}I�M�D�t�4�$k9� �p��Ψ~ ��������P��(
e�����'�Z���^ڹ]�S�G�
����U�������o�Mx���Z� �w����${_J�ڤ�QR�7t@�8�p1�*�bW��`n�O�����]��Y��J���gA���[�f�Oy�zo���2o���\�{8�jΞ{.&�Y�'��jv ��Ą�M���3j��n-�5��~>S��VL�����"rއ(`.��x#���,n�(0��n�A8F���_�Ar5��ױ`o�p���|��2�P�Kl	E(�����T?����3-�`]/
�lMt�E|�bF��L�6�5ND@^�G�nV��LT����\�M�5�;�kl$��k n��4Yh�l�=|�F8�7���D?�>�	;�����!(5���@7���`��Md,��L=���p۰<{���4�&w�i�ё�g�)s��c�T���s�$�أC��#��L0m���0��C��!<��~�^}q��蘨�]�W��R;�����C�{w�H-� ��/�vB��[�� ࿗��aߵ;,&F���|��Y��Aq�N�>I�|s��ӈ�8۾ p-�^$+�����t��V 4!���G��
'Nx��׌]
Tx�.��Lp�S�$����ߎ���22�ς�&������C(K����eW���^��g��+�j�� t�#ݥ�QҞ�a�#�:�h%�x�_��	�,{��٪ԜF4ъa�>��<��xf��yF	t�	�Z��&qD`o���3*��fD����M��/���[��hqq��5���n!C�ltt91L:=�[<$��-����S-5�_�?fj�'M#�-�N�GS^#`�{W	�JoV��O�h��N���bz�"纞[�]���)��ߢ9F�cϛR4%c�J褺�m�<'7�Yb�$�n�~A�~�i_/F�|��{M�g�y |����%֛j:���UD�T"0%U������]qJd�S��{M)�9�@��u	�舱���V��Z'�'��χ��u1�Ν��)�RJ�&���I3#�<�&c�,ܩ��<n?w��2�]�p��<nލ6��'���W�ͩ�C��0c��~�e<&��Ծ�#HL��];�5~���A�e@�h)� ���������`�D�ݺ!-�VQOH�4ե�~�=D41��{Kf]��U��T�*��m@:�2qm�f�Wx��\P=y:t���0-��-J/jKt��z�32�Y"�#u����|g�����Gy��m��V�{�EMq���t\��J�#�h%�ES�&&(��ȫ_��7[�^���S��ӊ�ɍ�r�=Ґ�h2K4��CL";���+��֗��)*�^�j*�f�E)�︲�`S���N�S��uì#AdXT��q�1�p	k�� �'����� -�h0ξ����� D��X���
��\��3V���LϨ�)��3T~������~�I9��"~��UF�4��k�����%�	�����Ʈ�� y��0@&�,��M��?	b0�angW��j�
�s���:�~�o�C�'��'��+������W���~����k���K	U�e�a*��1B�d\��-�_���ea�^B��������,Mԥ�vw�&����l�^v�E�AF��2��˿h���9:��1�����Z�dP�o�o�[O�������'�It�r$�`wf�(��4����[Z[�����8��S�Pn�.�s�U��d��$�:0�V~�P>J��G#��	Ó�+@��sX2r���n4^,_�B����b�}&��!{8�u�?w
�kѾ�D�d<�©2�`�]8�f@�廝���jf�y�2u����"�� {m�H� ��L�Զ�S���P5.�����
�^;�]%�ϘA�-�% 2=Y4�:iCR}~_�a	���p2�;v[��\�H~��{�F��l��f܂�L������^�3��g��{-dY�
�z=W�I A���J_�I���/��h���υL��̣�w��2�\�9���'R~t�,]�l�b����>�.o�c-�U2�5�]g1�3P�bo!�����Z�^�%
�5)+2k�6Ɛ��,�Y��]�0`�z�jLH�b4$�59��Iޒ@h��=:[id鲮�6��z�Cn��-d��]�/�����`����x�A齃cv�2�t��,�a�?BXgX,�q��1��ii��l~�av�P�]c�dqK�b�_w�ŀ��=E���,��8�j��|�wd��.ގ=+y��p>2����(�A�M�*���Y�����Kg���#0{ƴ�4��,!(��=���
dx�������h��z�j��؁�&�̳W� x��3��D:�� K��,�����o�����J�M�%�v9Z��8�������A!8��,�Ƹ�N�]%G �e+&��x!\f�L�7���`P�^��al��]�V��a��i&Z�X)q'y���������74͒����
L)�Zhx0�u�|�
IV�6�~�.��.q��PqA,!�|�.ϲ��o�P55}�a��B���XOV�r[Єw:����?|���
獑�gBt�2&�Ͳ�7��s�j�H��ߐ@{T���;�PR4e�.����8������ �k��o��@���)6�9�� 6	:�hKp%�;��OރW�.b�d���}��@��g�z�O[^�w�X2�D8�$q[��_$BۘЛEA��)��xw��6_�x�JK�o�'rЍ%��Fn$��&x�e��Bޝy
�\C��Ĩ�	�;��ӵ��Q��o�H�O�9�����Q�հ������/h7��M��6�B��Uu^�#Ͷ�q�~�3���5Ə������@�p)'tX��d,�dƺ B�u�"}0|���m�=9�&�j�!�CuQx��1���Ip֪���%�����԰�W�z�l�8n�*g���33O6E��G>�����9���	��0kbJAR�8�N4�l3�?�Uȿ����e$��Ҟ|���;�ZE�5(�v�R]�g�y�)��q�a�ɉW�K�8�I-���I�FZ���B{+�?��\
��֎�ύؘn��D�Y��#��~�����?��\=N�fh�4M�A;�i�;@����]�&�:MU�U������Iܦ��CC���P$�^�Dm�t�G�a{ʝ�����~!U��O�9�Q��_x��ze!���z"�5�p5X~��:��3���[��Ș;��rˤ̡��K�Ɵ�[F��������N�D������
B-�+�vO��{� |��-��%�;��k�k����C�e��ލ�,���J`�q������k�/�l��]���� �����D�Eh�r�z,	.$g���,��%\֜��sݎ���~L���W0K�d��&�OF���iLU5�!%���b�p
!zz	CF5���sr�b�Z���ӷ�]MZ��s,>�8�f�=�D��}fdT��eI��2y	<�a	b� ~����ݛ�0=�΄��fQ�K����lċh���t�=&�5vfȄSO�~̥�ހ�

��W�����rY���� �91P9[�F�������Bu��-&�ͩ�*�������,�H~D*���V�I�2=<���@�fF3����P����y]�*���)�yf��Q�{yV��ij��q�M��9M{^ӹ��u8�%.�7JC���F_�cV�VIN�L��,uԁ�,�<R�3>��m�u���J|�S;����Ɉ��5J�p�DƵ<w(��p��Fܤv��}I:�+�/��A�G�Ŀ!�}�Au��vZt�6+=$��,�	.r]Դ�΁�RK:&ޣm,Q�굊(Rџ�mi	�036O�C� \�|�j��^X ��ҲۃVP5-t�sB5ۀ��`N���7���>n���3Rq- ��1���P��+���^&S	~�!�D�h@ZI?+����BZ$�y��;1��}�����O�3p�m�
�6�]��P}|t��v�Q.�k�ޢ��K3�5����]`�S����@����D^1�kF�L����w?&���V6?2���t�ɖ�y���jnt9��A�^��܎=8� �hG�?1��� �sl�Y��������-#MM���p�h>o�l'��Wߔ��TX�������Bu��ow��ovĝ"�V�$
���E�r!I�S�(����"�2����E8�%]V����Y1��3�U]	pYo8�#`�Gj(y��r���9�xxG+�HWh2e�ʔ�#���^
*Y�����e�y�V�Epa��'�� �wW�^�����gO^���B]�*5�o/r��OT>5H�p� �ErY�����,���t�F��#���#���^�0��
���KJ������j�G����T�v����+F�a��b�*�s֒/av�����<Ң���OI�R�c��+���S��Z}@����u=@�	���Q]f䈮���e��c0D+(�I���)3�d���ǌΑ���T0�Z���u�+b�Jjv���U_��z�_���w����'s?ʖ��J���K~�w��,��~Ǯ*���X�+e}���ߴ
�o`i+�5X.pI�f�PJ�>�8.e��w��ٴ( �e��܌:Ń��Ӭh�:Ύn	��>e�_��$L;���N&}�%u�7z?���i�P^C��(�\��j��Ğ�Q��j�������?z#@�������WK3�l�ۤ��ͭ3G2i�rG�iJ���t�����of<�-��+K`SUЌ_{`t�S"$�g�y���<�R����:�94<�}�r*n�=��D����7�&��⥢�:�Ж�Y��s�l�D΋���F��/u� ���f�00M��縔cVs=����5	$�lϥ�����(�u��˭�l��<Y���a���!l\L�&�S��F�me�F6����֠&�ᨁ����D��pߵ��B;��Ȱ��i�D%��p���]#'�٫~�IRY�|�u�c����.ג��U-\��܊w�� �
}��&x�:��tsK�_�5��[�\}~y,`����t��V���]��"]&v�7��T�:Z�HB$�A��q�����z�K���D���aT8V�I+���'1}�#(�un�팽���Al7_}5����}^���c�(�AAsK~uY����G8ir��5��^��ȶ.<�p���_�h1�����P��B�e�F���RۙW��+�p���C��W7�ֽ��E������pC�)exq�<��D�l� Ir����4X&����5i.���Q݊� ��c����u�9��C�_P��?_-���^���B�*t�@³���zt�a�1���������e��+�(���v�PX}�,mU�����Fg�l��W�"����a����ʔ��+PľЕY�O��r�}�@�����f�jWT�?�d��?w�)<4�a���Q�#G,��1�r�����������j����=i��q�{=xK�l�Jw)�M��{��Fa������Iҍ$2�c��$��cU�m�N�ɢnw�Q�UW��nAv��e�um�JM���%S�٥rm��ɓ��n�"�d��TK��,��>J��0�ײ�-�Uu{��[��ՃUn��U��{~hBb
�_ݥ�g�L:ߤ���]�������O���/S1���D�n���<J������2�;�N Hh0�I�8 �kѯ�n��a�I���@��5ڪ�+$7�����9�䍇�P���^�)�k�֞Pt��8(�%�	�z��䟬vD �ሊ+Jf�/�~�4���g�rYH�TA|DQ�M�N?Sc��a����?B
y��_�F�K�~^�6�DD@_�֒ڭ�4���Y���/&��[�}x��?>�y���]\��T�S���3L��1CѾx�(�(޳k{�dʃR,�k��l�U �����7��c�����g?3�^g��?;D�F�"����S�y�gG�y"�J��a�A���!�=�i���Q���[�ͻ�� ��!lh��q!��KDl�g�������j�Nӵ����B��dp
S�[��ew��?p&Į�C�VE��}�@�a߯�cV@gNW����At_h�|�KЦ� �N�i(� ���b�8������߾��]l��*�lŶ�q���^�v����#N��Qn��7(>3K�GS���+���������B�/5���I��rG�sD妆8��O�F��&�)��=����8��.c��1.���ƠUHm.�!l�c𩄘��0p��*碑�j�G�!�I�}�
MR*���T=���M�=P�H�<�Z=��9x�H,�X6�{�����i��Hr�QmDHQ�L˽p�5��3&�\�/oP\�Y�fc��l2{OJ�m�� TH���I-j(����K��p��H?����Nt��l�ɡY���!�g�r{eIx�p�Yɵ��:GG����u�.)���p��SJ��������?[��B�z�ƴ<�O�	����W��%�C	aIj��I�\!�.X�3 -Vg%�ď�GSFA���{#)G8���W<��<+\ɖ�iXE��=�)��C�%��zԷW0�.��~53��Q�TzdCi	�M�7ZV-NV�+0J�+��.kN�T�So�{	P̣̕���;Ǫ�)yV���Ip�8��gIښ"�.�
�6A3�h��4��P�睕��iYд-�O��3��Bi����~�|rX��k(�X�#�ڪz��9Rw�[@LȢ� �0T'�.��!�@�����v���}5($V>�3���>���
yj��4d���I툶:d��R?�%H��C��N�:Wf�)�U��B烚s��@���*�T���j��+}S���0HJW�4{�<���U��Յ�JU/�A@9�*�Ӝ)>��NeP� C�}t*r��S��3zI���}�@�f�����w��H�?J�~��;�o�~�w�05%��֡u��U[�O�f���O)ow�`�L�)`C��P R
ޅ }ч�	��~�G
�r��� �C�OE�O��ёK�o������}ZL^?�eQ�����0�e��r}7��iQ2z��ډ^1`��bo��&5�i�|ߋ�h�G�f��֑��� 1�
��xwrP�+���s!>�� ��\��$���(|b�����n�W� ��F�`]��0���.�?47���6���^�~�d����hg���9�t�s��1�>ʙ���=Ru�U"o�i6ܛ����7��vԛt̋2�8�
ke��O	�=����Y]P�P�m����0
1Q�?�yl}��Ӓ�������4�2�z�{~s�^���@���o�����o��[\���/�k���8�}��9�����t�`:�.gx̎"l���E����1s�/�m.�Q���UX/?��h]�zp{F�����2v.,�(������\G�7�����l�_�6Q
��I�&J9�Nv �`���,�R�;�]^���]��Q��HT��	�lQ�8�G��9��/1H]e��)�:����ĭ�$��F�da�b��$�z�KCA�HriTA-�'�')�c���L{� ��yy�C�H7�z5s������r��E3]Z*�k��%|x֌�W-q���O����/9�?�����^�ºX�e�#ӫ���U�3d8�������L~��IrOR
V�$-�M�Ƀ^N�q��٭��,���_��GIB���J{�4�ӛ�>�����/��'��~^$ 	�{C������\�3D�RiF�#�Eث0�:�+}�R�j�H��W?�������K��N�`	�D�� ��� ���L�d\�u��7���R8sXO[�T����e�������c7;	�A�z[>5�:��f�+���(��5�R�����@� �څ�ga;&f��?~-�;Z��! �+4:��.� ��Q�;^tFh�!�ۂ������RI����4�����
��d�u�e�,��<xZ�6`�<�*����B�񵶂!�|<q�FtO�e� ���cC���%�I͡>kRD-*����&E�AlB�Xm*+��ϭ�; *   w���'��_��c�͢q�&xxIg�ķ@V�͢�������5A��8Ѥ����M��(�^Ҏ�>��u"�L}�>/��e����׼N �	h5��rC�
��L��Y�:�'��Ho1�Qu!>��y�ש�!���uh���L����j����M4c8 "�aԛHD��$i���J���+� :5��0�EZog�����"��m3���ʁ ��![�q�=(S��SB5�^��$`�kXW������9�S��,���+�z��Q��B���/����7��S�-j	�G�ƶ�/]r�3��(�ĭ5*-�@C�>���u5�R���S�d�=�������
i����/�D�|�#�ǣ�V\ц��A��ƚ��g�'���j�h�S�b����^*i�i)��8��a���L�מ��`.���[M��|�Q3t&x�������ݯ:�N�Ǻ���U`��%��W	G-��Q���y�IW��ڑ�fJmq����<f!q�/(E�z� "���Mj91](Yζ����;p��m@ܨ���L����)��ӨR
/�}EF @�J�3Z��K�f����ݝ��:���0��7�g\'Y$����Oʐ�T5o�O��p��Ѧ�x}J\E���4���ۇk�=6�M�L�(��gZػ�pu5�*�(�ʽQ???��h-��}~e�V����ɨ��iΨhk��R0E�p�!�����D[��lh�>!�/�9D]jKń�AZ��I�~^ +���Q��CPn�(F���<^-�3 c�m\��]K�ŋ�˿Ǖ��A1UB����M�|D�!�E>з�*.��vmٙ�����i�[�n���|Iz��9zĐu��3���qY
���_��DH���&v��F���5i�<�r�6���L�1�:RsE��2���.�.�q� u��,+X&������n?��A6���Ύt��0~��0�fa�v�z��D6tK��hmFU��?��3�o�Y�k�)q�eA�9�ߘ- �-��Q�O���:Q�d�Ow�o�LL�D&y�2^�x���"���p�ҋ�K�`/
�Ϲ�vc̷j��n*���;bBV�'=�:��l
���
Ɗ�Gx`>��B�F�)[����+5��7y�6�EV>�̙��Q�R��8�Jݯ��9�y4=]���%�Fp��O~~�c��0��o0����x�>�n��spb�Y�Bt.���?�kg2�W��m����X��Y��i�N���B�5w�\+�P5v*ד��F�~�t�(Ȇ���RA�~������n�3��윜�C���!:ЉO퟽M�]�����eo�c.�o(O���dJ�ޒ���Pm�4�7��쇟lB`���
;��\r�,`�AրӤ�ya���1�����F�"!�u/"*�*��;��s,B/O�DJ͹mE��(ȄN�f�����B%��wd2��� �Ե�O�"S�em�"2��_��m���qS��m���k���%~�zb�R3�~��k�kܹq���°8{g�0wQl��VDgY�|7x������c���l�6w�s_�d��E�ʜ�*	��I$�������F�锡\��b�`]Aq����
_:�)x�/�}Q �e��9v���jL�����L޴P��cD=��)�Ｆ�/�,�\��e>�g-�v,�j�����;��}��q@�����3��8�[1�M�JF>����$�^{���i1��M]+��$�7�h�5�2��ת���7wyى�[<�n�[�x(����	��6�����` n��)�P��k���u��
_,��!�����H��SK��XE�������������\ӓ�#<\�m�&�s�Q�dF��3�7����#J�-�a�-UCcc_,�N�eU�#\�����U s-�{ov�.ԩw�:ī8P�g;9I�!/�9��1o��;)�B�J-�G)Z�G�>w������|@T�Fiu0�]6ř��M�5+S,o�ךd��m����x��׽���].ݛ�Q!�j/S�io��)�|�x�b��	L�0ϓ?0�H'�N�[{U;e��gK:��X��k��_�ZN��{!�%G��GPz�S��,՚�(��(a8W=1�?��G�뾣l�'C;h�E,]pR�Dk����(NE�4:��,��'cٞ�A���ɢ���������X�]ڷ.���g�?�$�p���6�󓆫�� qM����4IH������Ć���8ٟ�����͗_�X���j9�L�c�6�^�d���Ϸ��M��ھ��������԰q���^��bhb�O$m��	���[�e� Nw-��u:?[*z���f.��Q5�	Cک�ϦtD�:�M��E4$�1䊺�f��k_s˕Œ�'�f��D\[<���of/=���#_ne�:P�ѝf������e��ެ���?H*�H��M�mpJ�P}O�W��D�q�WMӪ��q1k�j)∛aB��2����\�޴����Uq�SP�.V$�"Ka��N0.���u,�W�:<a�_h_�/+Bb��[ ����-!�Z�����>S�Oח�����m�N�E~�ʰB�w/�<z��p��r���Io�C��R�P�%ΐ�&��=i��@�d��I�>*�l�X���XI�ݭ�qa��twc���B�O2��26�y}s%If��_��8V�r�	i�M#PB2 �"��sш�\��w6�z5�&�,�p>4��lq�O��KF��J�8bD5���NmC�����SgJ媊��������_�D�,܅,Mo���׮AxB��\Jԕ��nR�$���sr�pbM���z���ͮ�:V��l�}_�V�'[R��/�O���Y��#��z{L>"Q�'�N��(C��s=����q��XzRGH_�8/x���Fd��n+~<�)NWE^�*O'��Ph"ֽ�R�g����ߔ0S����'-�O%����J����˺��}o�F�~��*i����Z^C�����~��cmI�D��0T?_�f�a��Hu^֭:�-�q�PV�T;��&n�AlZ�񁶓��hxu�Ī�q^Q��a	)Z=LK��Y�ٴw�J���Q���ʵ��feiJ�����ȃO��`?G�}Tz40��=�u1 ��7�DuR_J�sl�G�(��9�Ve�u�󫎼goi����CȮ�$Y�U;$��++_�A���F�ۈ1�M	�kH�v����s�Q��=J~�SjW�}�ǵ���������+�l��l�:u�FP-9�O�yI�pY�����ch
�vP.��׻V]���D��c�����:?ӮY�gwK�ɷ��&�8�TI���`:�O���p[�X�[�"B��F�x��W�ؕ����R�U~���{3�ta��mv{���ZLW>��'s�t��Y�؜��Mb"FI�#2)W����KNCd��*i��XV��?�'I}�	b�A��+T�C}"�ƻD���%<�������=��mYce+Eu�vR1��	bXz��N%R9�5jL�y˟ ��d�O?�g�YS�m\'�QX%J��8jV�F�4�D�/3"��s$���!뼮���㑚S�0�|Zi+f_ObK=� �ҙ>���8�6��q�M�<���F�O�������[c·�;�eL�}hEI���e�o}T ���p�N�8y��X���\�sY�du��� ߅��3�PC��Qɞ��|j�?������[<)�ⴜp}�,غ 
/��4i\gէ�T.�������`ڡ��� �i��$�L0ƀBI���n)2��W�y�UVܪY×J<�i�Fh+�c��ea�>��&N���,�8ٕV�ڬ�)D�E��O��i>ۏ��,�7*�WKm��P7�����i�@�ocǾ[1Dv��I�U6dX="����ѯ�F������?�8p�H�Km���1^�4�<�2�ze``=�i�s�ą�UƢl�9v�iѢ�br��R @4��u���c3��P|4N�
���c���ҍ�y��ٻ��'e�i�I�&҃��P�ae�%�u�=~�XOg�������F����y��/��r	jU5�ĉ��t����L�	���~,�l|�澎�o�M*�f�X���yX����7�z�|巳�>ct�l�Q������*�����cv�#�L2�!���3n�W�F���^�&i �>
�A�Ae\��"���+�ȑ���n�����J'V��	�Y��J:I��"�����l>���V��<�:�<P���qE9�ʕ.,N8 n�1�IV�����16K*D7�;��ܪ���x��2Rc��G�zHa��p��N������ ��n^�ǀ�»p�VBʰs�O�ġ4&��1B��P�S���40�N�^�S�>�{Jb=�x�<d������.D��F�Z�d6�!<yʦlu�G.��FB	��P�EΕ�U������TL0�e�P4��hE*����&{e!���;g��liaЪ��c��&�1Vw�\���+�(� �38��&q��'�!��5�ܑk��"�r�(�IZ�"�T���[1����Z��<��H���c�����-�����G�n�QJ��X!�'pQi51������8�«��V�K9��e8-UڨK7���vq��V�V�/�$��`aD]�`ݛKg���#0���g_�+�"K_��-�Y^X��̆�.�0%V���'�����汥 �mТ����v�t{�D�׾N�R�uI��*ꃛ��V�Ġ7v J8�~�W�p~
�}��Cz�P
�Z��{�Q� l�F^\�Q�����W�)��<T���&"��b�o�0��eS�#;�v��Z��/��]�K)<|��Y�P�PJ��� �4��9Sa�4-h���<���0���P[K�`��~�CIR�(�����k��]�����&|2P�;���5��ۥ�[ɥ���A��0?��/DKpݖPΡ�'{V!z8��E^�Q�C[�fUr�8��w�`��3h�����$H�W�-�?!�]����D�Q6��C��26�F��4��I�+X؂��@7��!�����]��^�#;Œ;���hQ���hI�	*h@�ta��c����b<
��SZP����r����7��Q�C�i�-~v�R��:g�X���k,��*�bơs��0��c$[a��43�������ݟey������uH[Y�o?����;���qÛ?	��dkE�g9sh��}�T����%���jQ\F�3)��ml�Ʃ<�6�wփ��i�EhR4{�� t�hn�҄�P��dk�.����}��Yt�M��E�ڗ�	2��%�_�t�`U;����*����·��a�u*���|�;��FǢ;b�:Ah
l��%���J1�3��H��o��?yJ�đQ��10����ۡ�R�C��d!��A��Λ���v����J;c��Df�nf~�����i�\Jd4�p)V풩�n4��������ңq�O ��[g�琉R!bw��$��!��BD3�-,�(l�7�����p�5�M��_��-Z3��ɉ��R�5��*��7h�=L�_���`j�b�@��W��{O�P)���aq�Yx�v�����xm���^s����DS=O�k��\�'�u�j�*�k����O�Iz���sU�M����R�]Ũ�E�)\c���(I26� ˵�������\1�8ҫ��A�	]�e��}2�zT�ٝP��iD��?��L0	�㻯Rt��nn��U)��)�,Q(���I'��0�t�M� � ,���3�`��a$���G�Ұ���n�\�㹿G��w�s6f�H��]<�Hu����
�o�dP�,�b�AK�Mo�`��埈֕F�EąP
��{���L�Qx˻d�lG�3�Y�.I� �n�JJT�>�O�ʲ�ag��LU�E�Yy�(l^n�CT����\3�uT�X�{Z�3d14;<��`���Xu\�Jb�$��i�Fň��h��ۊ52O��Y!nus���?�/�y�'h�ƪ�o����ۢh�(�W����>͇Ϸ�ؙ�(��X*�Ϯy|.��������`ܻ��L�	���r�!��8�װE^n�V)�������MՏ�-��0��q���_��
6�*�f����Ѿ�_�'�`%�j�$�}+|� `�qt�X��-��K1��k쓱�ו [E<F�l��R�Ym�Z~ 2�Cے�{�|��,~]Pl6�(>ad��"4� }�`��ԣ@�F�����B�re.����x�P��3��_������o�c4Yա�-H�٬g���p�tކ�����z�ѹ��N%�ӋX���S�x�Ddw}j��Ҟ/d����\� ��BsR���3|@\��3V4p�׵��<xˀJ�G���=��j�{�s5Bi��5y���"��I���
�~ޯ(X��!((L��{c-;� =�b�i���XD�Ǉ��+���a'D����Ĥ��Z�yg)`O����D����S���pit{�t0
����)�� ܍�p�?ޙA�+(�݋���<52���"�F�5�Q@Œ�G��9�q����A�~2(̐�Xqu��e���o֘x�ب��쯑�+�:�H�������;��Β�����>��o��oȻ8M(��r�9���b0d-	]Z'qb�p�9Oy����(�{>X�(>�x��z�q�\̓�E=C�ɿ�.v(9}o!��ڀ�O�hn� ?�;�s��̎�§��*�\5��E.�}����	h���]/��q�ǋ�t�?�q��)�0���NTԲ�)Ivƥ]֪*�h#��3͟x�_/[g�6���+��B�k� _�7ҧ8�W}��zx�ӟ�>�4*P���髢���O/���=�`���I�˅ahǯ�$��b	=*s^�cW�ޡ��q2W7�����jL�<� ������~W���Y	i<�
��R�2#��,.�ٴ7S�����8�l! ���c�E�W#��^9P,F ��n�@U��/d���>|��f���_����r��@��bK�IF�S�����<.G��T�ŭ����
��k���g��?��e���k�]Æ���j�U�)⦴��;�&;���� ��X���PB�X��k}`�dX/"*�[����^]aͤ}��=ϞB��r$�͈1�^��C�k@�0�Ht�O�|*������L�/Zʭ��3��P㢤J�<�s��:=}ȹ��&hwq��	,���֚?�:i)Ç��}:Ɩ�q����0�*�!�/,�k�)։�O]"�}��?�CR��� Z��Ɓ�MG���$���F08�\�O�?�u_��N�v����EyX��M��N�)�����쇾�X��p>yI����#��0P��F��tx�2��_N�=Z=M��8Я��iL��B0�xvc݄ފ�V I�1���2�
Yd�����W�膐sӠŶ�d�dv��u�)�o'�#=$>ndE�aQxE`]��I�]�&���r��ꄤU%O��ɓ=H�p���-�]�P����u>o�=�=L(�|o�����Su�ĳ�ԣ2N���U��p��^��bFs��4��Z*�)�a�����x;��S뺷���j��%dh��c���/�L]Q���)l���8IE���G��͑v�5`�\#l�ߔ�J%�9��_g^U邓j+�ɷ���=kgjAZj�]����,j8����2�c���+q�Ձ]��W��Q΃��cf����M� ��`�b��Ȝ�L0,m���X��ZB����,�E�F����s��Q����f���I�G�*V�3v��®l�W{*O,��O�.�G�ژ�+�)��KGuu��ް᥇�%��VobbRx#���v���t��(��uGL�V�������v{�Z=
\e�G�7}��ˮ��&u��q�໌Ϳ{��GX
3R�mEA��N�����U�g^,���o�ZN"ε�^XvࣳR��z�̙L>��Þp��?W�����=8]��
�&�H�=����#�ޑ��h��m��x�,��1�W�F��_���'pC���AD�,w)�[yG��n&��M���O#%'����=�fD�����m1�m������b�I�-F\�I堵H��/Z�����d�S4ꉶ`x��1��y@"���etX��u��m���>2��qÄ�G�*����	*h�F(��*�EVQ��T����wL��#��~��`�G.���4wZ�1���M�	�O^�(�vT-ɒڰ�M�951
��:�9Q����#�	�����wTK���T��R(�K���
�?�G�=�(^��9��~�aW|�J?��	���Qa �5�,OB�>���,0R_낈-�I�>��~�+Έ4�?s7�$//���m����z���ʍ�R��~���_]�D�ƹH؇��ӑ��;b�m��d�X�D��{��;���6[�/�@��t�J2W%� d�le99�PM��_�2	�u�M|Q[���F�_�z:t�k�����yL����RɸR[co1�2~;�����]��pgb:�N�
O:TK� H�.����x��T
��sC�W��lL<)P����RvV�^o��al�o�2���5����ß�!B|�<�,_/{phҴ�ioI7Ö� (��0�0j���:Kt��t~am�8�>�;ӻΘ]r�e�.1�|�&c�����%��(;��e_��ے'Y�׃eG�Rx�ɞ�.CEQZ�w\�30c;pIaK�y�H�H��x����Ci������;1qD�x��M�j����q�J%1޺�f_�e�H2zb�����m��݃E���<�7_/M3�b|���R�# "�果��c�붘`]�A�+Ժ��OA&6�.��nߣW���/K/&�'�BB���_��C� �2`4J� Z�':� �P�fM 5/	⋼S���B������pDii�[4T)Z��k#��̐����?9`���JY���UX����DK��9���[�}�#Nk�>�R�h�8���-�o�3�iDVLXz.�oa�&� ds�����TgKj#5\9G�w����+Ⱦ���<�񹅿ms�L��Љ3�\ ����[2�9��!#s�IjD"3���P�n��,A6�0��עᚸޭ���L�a��ֳQЭ-�+(���J���b���w�uݢ���rPi��7h���h�
���Ƭ�~�6�-��x"*�f|����k	5�e����{�{LrA|%�����5I�3�Ť5b�Auc�o>z԰��.��<Ll3�Q��fʽ�yNs���I�s�A��~<-Q'je2��[ �ᶍx�+��,R,�'V�B��вꬍ��@��-��2�ݺ�9�1Rl�a�j�}C�$�+�f�?@�/�?��iϾ|jV�)����tX��Z�>Q�ڷ���셴�4�g�R�ي��U'<��\��D��9c�:$ R<B�iG��^u��@�"�︨;��|ME��Q=͎t���x�M%_2N��n��۴�Q�R��lV�����ʣ�l��f6V�̬������?�wق�Ƽ/,���#)9��p��s��\������'i8�9����ǡ\��=A��A.0t���(��9 �Q8�稗�7�"���`�����T)�n(d�>ϲho<�� �-�sdI�Y� �k+?�ƗWIS��I7��b�T�fS��`
D=(�;�͖wV#(���d��Wv�����ψ�� �"v�"��A�t��7��"1-eB��@�Q�g���O^�	ƞ'��S�����I�V#��.	�4��M��cd�ǀOl�ôE��l��e�Q�qg�Ȑ�Gy#�ѵr��]蕫�q�q��� ����~��J�����j�,M{�A���EyE�#xh�+P��]�&(j�n�D�c��>�^	+�q�0�Jz��?t����!�J���
]�-�tP�.I�x��C�y��jϯ��V�.&�9��7;�d��� ���\��?�)��� �]��+0 Y�R�𑘢��P�P����HN$*����-�᧊�H9`x�������Y�e�M"E��qn}	����)w����/��}c��!?��S2)��M���O�/agR@F�^��E)���P�y�����;	�����M�r��@�!"��QOg/A��S���6�z�8-�L�j���[w�����w�/Q��.�(��g��c���)�x�(��lI.En��3�j�t�D��R !�X<3�s*��c@64 C�RU0��s�_CD^�]p1u$y��0x��.�	�}!/W��a^{�`m��i�(!�He�˽/T�&7��XM>!A�0/�_��H�sDy�/GIj�_l&��j,���v��9f�F�c�bjJXI��L��o{�*�̜�����1;��K������NZ���ť�"��U�����]��zZ��닱c�@K�I�uN���Yq`%���zOT6'I	6&"V֙Ao�J����P��/χ��":W� �bV��Zl�w�h�Y�Y2�Z��p�]�W�k��d�t���ˇ�>�)��$�h�v��T�+kͩ����-�qbe�7����	
��u<x��+�'����{"����j�{6p��,gl�#0T$yN��g9Ӊz2>nD�!��������I�y�8���s�����rA	rf����������/�+��?.~r�c����N�.����i��{J�y�B���=Q:4����9{U陮�N�qK�����Ͱ��EN<���]J�96�"P��	�#��XR�_������v�hp��f��o�4T��'e�0���(}�Ё'�~���U����4��КO�K*���!�>��5;�2��!),-2�kb��ȥ%� L�|D�f��ab�1l�Z�,�Q�Uר�v��gy�4[��[�\v^qg!2W'������V�B�i�/���Z��;zZM&�l����?�0�Ò�P���XO�\wlV�=�j����>M���kS:��d�Q"AJ�NQ�0:`�ߛ��	t�'�ޏN8�;���e��w�pH�ݛaS>)�<����xG��Y�c3�g:u�ƴHr�����Wݗe#�D+D��e[�O#P8#����H/���:2�`m�ӎ�����{��1��ߤ9��&N(���I�f���m�{�@��n23]Fw���d�,�ԚU����E�˰�x�؄6��������#��
�6ɀ����y:9ˀ��' /��Ӑ�j8�Kz��O�ӒN 3������*,\���ϷZ���w�rV�����A/9�S +��R����L�_����e�i\�˥Ũq*�MR �٘S'���k�Xl02��L��������3�����K6�ft�Odo=J)5��Z߀�m�0P��Qd}��-AeT�ə/���*I���Rȫ�zW���$�A���
?z_�
���?u�K�9\�b���Dɴds�d��x��R�&��4Iﱩ�!<�IR#����a�WiE��Ž��E�w��?<T�P/�lJ����k���Q�p��x�$*\�\�hXW���!�9��߄m����vp�S�x�h��Xz��(S�q<6���(Y���h�K�-�S�i1� ���>�v����a$޴Oo�!�_�	v�Ҏ��$՗gc~s��F_�v�|���zb��6}�h��� 3�q���A"��)^٪.Y�x�:E@��ﰿ�P����w,���5��V���J��U�Ӌ�s�<ۄ������x$"��!��<�5P:�r��#'D����!�R�AH�$����k�����U�J+P��3v��2�K�Iaد�F�`P���%��l���RJ��j�c�	�!E�-ţ#�J'8
���l��9߱�.���w��bT�T���/p��3�"�5�Q�P~I�-3���������i�����5H���|�KD����k���4@��"<�9�D���>�R���Ӿ.�@&�ȅ�φ��RuIp�:����ɜ+�3g�~$�lT����j�io�_�4C��,��tۯ��k_17��tϝ��:�`	�����)���f�
,��O䦿 �����7U�9��w`zO��=�}�r�#��	J�V6]�3���V��\L�=��o$t8�D\���Ҽ<!�g^�=��ٵ,%���/��9%��n(��*��"Yr��0�!��3�N*�j̫Q#�_�gd��^�8r뺴Iy,x�,4 s~Ͽ�V��1��Q����۸7F��|)���,ċ���G��6�����Q[��H��/Ø	h���9��΅a��ʑ-@��+@܎1�	��RQ8��Bx,�Tj�����%?~U�g�R`5ǭh�^�����~�8�e�n��pҏ��F��pڭP=l�~ޠ���H��^_�Z�JRG���y����O�ł�֢U��)1	��U۪�UB�)��d%�V���������Z��-VX)�6����t�p��<<9���0 Pz�K��Q���e�/1�lhӆV2��\�DT��ilm:����m����"R�(T�	}�x�a�OBܾнf�M�+PPj���|;�:��{�;"�j�	�SK�$����Z@���)A{�'c�[P��((��ǲ3"��s���� ��/����d��|\�҉4)1y�LDF {5�~f�c:�	F7�m���%)��o��R�����\�4�M7&D��vᐓ�>}����z���7|��'n�h�U�U4���;����S�q=!ֽ�+,ᘓx��S�j؎��3�'>���f��%��b0�d�6k���/v(����u���4�iB�e���t�xu�Cv�-����-�|s�ۗӿv�~;����Z�@7j'�J��1�['���3R�����M^�*D�*�T�r6�߯��.o�**�_����*LQ&\⺾c��>NE��5�z?mq�v�*_ЈnE�«/�^�l���3���o�����^�F]&�f_�]�M���4ق��B��C퓎�=�1��xlڏL [�o�Gs��q��K��J8��jv�.��Yt)\r�+�%��j�Ko���G����g3�|���\G�������^U�jk/����m���b�{�+.�M����6��vxqΘ�pf��^vg��͡� Z�{&pW�ǋ]T�7�Tj8�@�����&�d��Q�Z��bHe����'�m�z�|���݄_�1����d��bΥ2Z]v�3*��1�ޮ١wG}�}���ª�
����� ��3�d}U8 c��>��m��p22L&���+k��c{��
9��υ5�V�P��.@� hi�X�#������������	�O�l C.Wa��Udk�v��"�ެ�R�a�D�+$8�����M�zg>@{IP��t}T��ŝ�/z4����,�e�CP������y �c�l-�gq�v%�׸Il_���!]��ĒP~���wG%��fz��0����!r��U�kO;����G�d߅��a��~_����K3grL�$�[��('��3R��>��Rvj��MC���rԧ���j{�-���-b4�ƼPvE��.,Pu�����-ׅ���Ã|��D�9���J�����+ǩ��~�d�=�^��!}��e���)�L���qh��s) �^��(J��lDȸ�*4ܽ���aw;Uo?+�
���c�)���.�t�����8�ǂm�� j�IW�5��#K��.�*�65ދKBȕ��ǧ.���%ts�_���|S���A���=��SЙa�K���Jmȶ�
H��/��5�?%�}p��{��r���ʏɐ
��x�ͩ�� ��L���^P2T5���1!���̕��ꬶdc��T��e�B�5�9 �ɩ>������B��KQ��X9	b�[�y,�l�o? ��a�A�\w�����*ϟ'�m���_I����n�����H"��ΐ�Z=��6���h�gA杤	8��I��)tx��RA�O�Q2{S��G�91�O~�fL!U�>M��dT�}`��ܨ

Y�YV�POD���[��#h�dm��%�)�p2���c���X/�쇂r	l�B}���Xd'@���,B�gm��K�䥻�	E�ɉ���6��j��FH��-ڷ���ѥ[���fJR�j�3{�K�Աg�>nE��eP���Qr�kd)È&�ylet�s��0� �.5P�L�,��&��>B���-B����wL7�h��*I�ܲ��z�q�ȝb��G�)��U��8���u%��J�۷j�s7����:���ˏ��rN����"��Ra�'-M@=�5���n}�Ί�ٔhr�U#Sм�5�^)r���FNY�j�R�/ZY�1�~�.��u�(k��u��k�Az�d��kʅ�S��o�+,Ou=h���5^�	8_(�6z�5g_���x�����óU�q!(=f�S--�����0t+����8��d#���gt�%m�D�=H��iڤgӔA"e����%v�偱�Y�"wTKeG�~=>��+l�k(��0�#�m=� k�eC�(E�,�:U�[ϙ��s��3�W�0�i�(����|�մ�c9L!�jj�t�Hؑx��逛B.��iA��&=Cm�V�*�L:����������rAu��;1��������4�2��	�8���A���½S�5en�}�y!_K��R�N��U����g�do�#_�C18bY�%R�-��s�:����_�hpR��(A�Wګ�2w�_�+���U���T��O��(�f��߱z�T@�=��A8֨�Y���!c	ߛ��V��Z�:,9��1y��H]��[�E��i9�%���A��!��j�'ۍ����OF��B)V0���El�J�J���Ϫ�k�U�ǎ�D��S�]}�q�7}���4��6E���U�w-�E
��Ť{�͔����-���AT�Jɾ��3	\��mU�c� ^�2\�3�z61O��k�zp���B�����Sލ	���8����s�J���OJV��K�e���=5���5���,�C�5���6�Iѩ���;�	�]������N@Ľ�S�������w��ѩ3�bR��=s0qd�2��t�*�h�k���)�O���c݁�}�MQr"��� �'X��8`���j����F�#�*��x T���Jj»�g/L: `�0�:,O�)=�V��p�^��{X/�Ŝ��H��\��w�)��ۏ6�;wL�ޟ�X/�2cG��X 7&.���y6�EK伅
\F��%�'ߔʅt�E��|���B5Ѫo�ʉ!�)��|�-�m��.��ޣ���WX���
����f�:8ڙQ$��O�S�ӻT�Ť�ؓ&ykƱA��t�o*�%]&^�euBV�:e�Dt�wW��,,�Y�p��nV�i}���yb��~���|L"B��a%EY@����Rt@@#�Zi�S�-RV���X?W�D��N�y�������C��*���F膃��57^��̚Ez+}��q7�{K��ah�DGx@C]�<��M���-a���[;�DF�3o�Azn��j9k�^�-�k9����_��"�cߛ�֙1Df����=�OU��V���j)<�� ZUDb2����g�R��\����os�g�V��]��ɫdݗ�f�;OlKV��y�?�N���j�����8��������~�٬G��`է�8-"�dS,�^�����>�1�T��i�$�EoF���r�ҭ�9����{T�ԸM��o�L���O�D�i���t��+�e�Ͻ�"��kklƉ���Ѻ��|�!�~>�!u�C����߄����.���0l�w�q� �H���H��% 	�ީ� ȱ/�\:~j;�PW���-	|A��$'���~Po�ג�?���ZN1+c;ZK�6�]��2?LK��0�����`�Kn����p:�.��5��۬�Z�% �1}�|I�2s\���
>E9��_N�C�ܞ�ӂZ��6�O�l��d�2p�=S`�-2��qn�/r������Jj$s�}��vٗY�<+�C �,��S(Tŭs.>��k���Vw�bu',��i�L��5������g�x�|ۏ6�N����y�f}�ͦr/m��}������<V�a7�y,��ϼ�L�_v~X��I�����T��2e��Kp�F�����}#�7�ި���,�J�w��_�j����C�����X��F��מ+dj�C�l��<����0��L1��$y�c�R�o�i+����RY�}[X���[~�e�(A�bB�!l�!pA0��T��!�jՍ�Ϧ =�4��-�x�C�t_���
���I-��*�[���Ԣ�����>�Om%���n=��TW*�Yu�\�:�b?�\��1���G$���il*�^�������e ΩV�5�e0A��$8����D�Ӓ��{�I;�a.�3���nG�];�s�kS�c-�ߠ��8M��F f�zc�h�7v���7��5�W�*�Tp��xQ=���]ci>08����������@��V�6�U�ϊ�l��~�9]R\�B�)`#Z���sAT�*:
�[B�MI��4�m�l��g*�|\Wg$3�W��]��YR��$��R���ɘ��Պ/�MkʲŁ��L��ż]��Dm.�%W��j�+E(��s�����2�ʊ�Ϸ�F���;�*�Az��@V�ѤX^D�
l�}ȴU�,�qށf�$+1�.�P���2'�	��Ky4:����NV|B����8!7�d���4R����UTNjj`Dh�>�v ~>#���7a�1z5y-����L���d���\�|tΏF���{5q�<ڦ�vH7���hk�*��Dn��_�Z鹎�H%��Z^�n�F�!��`�bN��G&\����Z&�<1��:1:���m� ��='�۷�5-�@^:J+��p/����G
٫")ݰ	�`7H���m��� ��߷}?H%؁�h�aUe��2� 	9
F������@�>�^O�(����	~�E?J�f���VV>����n������Eg�5갈`�?'����(��\�"l�0lh�f�D���V�ek����`5�� ����jS���r��3�9�m �0��_�l��GF�0q���?����y@k�P^q��0`6��4p�����$iN�\M�����#��MO,xs�������9o�A���=A����%��t�4qќ�-/����1��(J�8p��يAy���.c�f�ꆔ?�����8
x4���!��%VUZzф& 
�z�"4cD=�;��*l�ҋ�0 	���� �Vee�C��z�|:H�u}�~�܄r<:ИٕS����S���~�����(�Q;G�F��D#�~����ֻ����'!���·j6�X�ٴ}G��<�[x��29J��,��g����4�*����o�o��M���'bT3-O;$��r��5��A{/���jA�XZh��g�vt=ŏ����i�������|2�@��W��k�U�=23����n�/��Z�_U���)��=A�"�fC������J�� �&�m�u��v9��^��H�D=+�_\z,a�O�(hp�F��^�?\�k�=��H�&<3�9ܖ�>Ү��	샂|�d�ĺ^q< p��P�/�ɿX��]v��!��qS�P�p��<-� I�+�����"�$���|K��1��T�^�p�t���Y�J`�R��5wI���R�x��!K��O��Z=�g(�����_�}E�ͻ4�w��7\G��,1� t����R�;� .rF�oe�l���FS�
�)K�\o�,��SJ�Op�"�)n��àlU��6�2��9`+@%�(��c45�7�ލ��T��]zE7׭\:Jڄ�==u/�Y%O��-n`@]��N��Ij��%����k���UF�%N��/�!֐�I�V�����6^b��S��G����J�mHhCA�O�5�q�?�5�sx���䎿(��� �9E�sj��bT�G�}|9�9G���x��c�_su\�댊����z=��)X�ǈ�=��ol-K��n˾[�[8)�d-z�w�,:�����|%�c	4�n�`�3������O��v@���$MB��oI~�Ԑh\,���l?�?,��l찼����in��<�y�1E�����F=g}Of�nE�c=�9 �	:���E�m�A&9�خ�aڂJ���-�x#� 7���2�� k�>�v����D��i���V�����Z:>i���[��0�q�Զ�,��͎F���F��?�֖P�����P&d��%�E�W�C.��P��pG^0�����J˚6�#N-��ҲI�H�f᧪��V�.����x��� [Թ.�&c%�͒�EzMz�39<�K]f���4�yAl��^��I�3�C����ڃ�@�nA�[�����S=FM/�5Km�^���A��HC����􈇳��0��>�����%{� ��wqie�% _Y&���X���x���ĭ�?����t���I�ܪ5w�H�� 0��X���JPr���K��e���5�ˏʾsO�c\�+�AYd��w'm@q]KVF���|:=s�oբ��_�tK�zQ�Hvz�{�JI�lj<�	�#�H�I$x��ăMehY�	�|	��00~j�W����R�Z;��̒�ˏ0�?@0*��#)m|�h�q���D|R���z�����yx�_RW>���YrR�_���7!��!�\�M��KbV1O��W�|��D
�0��h�[������y��%{��7HQŪ�q(��T���B��7� #�ͯA:ux�F2�� ��M�^��+T���ߛ��~Ǟ�`��2D�%l�9���cEط��7)P���%�l��As?�$�In�}N�f������N�盯��hl}�����JM�����4�]�R�^h����H���lG�ę���&tj(ߕw����慞���S72����qf��?��aj�qm�F�C�o�]0{�)�zDD��֟[�2���R3�j�2jJ�V���$���00���8wڋ��,O�n1�SJ&N��J����^sB�(KĞM�h&8��G8�wl/��NgŌl��
�O̭1��O��5�ݼI����#�F���T<Σ:��n���~.^17>�������C�y����A�톰�%æ����/�Ɠ0��)��vma����Mm�?I�$'%4n�@��Eǝ��Xe�f	���c���)�XLM��sG���]Q< �Ɵ�r�y��Q,8J;����.���Ž����B�L���R
��S6�
hPU���G�h�R_����7 ʝ�LϨ�H3"d�/���>3̠5�Es�PV2ծ���}I���Ã;D3T���%?%L���@��NB�$գb���	��(���N:��ucva�~Qs�S�nJw-a�{y��>��	 ���4��kɏ�N��Y�� Q;�ĺ��f���;M���*��.����*�S^�!p�`�(�����6.�����dy@���.��Op2W�DG卒��`E�{B-���ظ��$#\i�X�8����95���4Q3��	M�0�z㗥�r�����8.�B�僐"�*�(}�*d:�)\���G`�����28�R�M_kFyִ�%�k���[����#�㥨;8�j��M,�ǜ@�Gv?~X�YA�_�q5����`7���"/0P������v���v0��
�۪��¾�(�����@����M.�f�s�+��M��&����V7s@�1Z� /P;SkǠӳ8[ӯ9��ޛ����i^��?��^�G>j[�/E�@�1� ���u�nz�V��5鬥�3��DHÍNI�A���deX�Oº�oZ8�tV��ϩ�*�H��
�Hs-���mM?Cg�oO&y����_f�IJ5�!�{_mm�pc �m����M���fn1S)WL���:�v܌6kʫ�o}�f�b�|C�z�,i��^��T��~Y7Ĭ4_��g[��7�U��;Pw�p79{���k��K�#�0��SwǕ�8���%� �����(������5w69/e8��2�k<�`hy�;�ߡ`'�\��bG�Wڎ��XQ: �R>Y����3i�3\���ϝ��:]W-l�T�(E�$i��I�AA�_�Tj�]�����g��kn��">0!�K�	u�s�����=z�5'o�����΂ �1u/}�<�H�q8��įP쵶j�v�o�x����X�İ����!X4���l�����$�*۹����3KU=�Jv��d̞�l�Y�K�5J��N�s���]�Åđj����j�!+�BT���~ܸz�NϖN�ڈ��+:>&B5`G�#[X=I�f%O�+����*���G�H��u�Y���	�cF�����:F�2!�@�y�c~�?��x�dIWw�!����#�����r��:��ňlDSLxyV��p�Stb��$K\���Es/?1��j����9h����}�`o��}�9�Pq��@^���y*I�~� 0��Y_��r+�ó*h�7���V��[[��!�#kH��;WO�)��V�UL��Y@��_������T/�\�Qo.��S��m�Ќ�6�,�
?��b@�9#؜�XO&h乪P��4�?S��ӥ�峴1&�2����q�A��V����#����#�t)8�~v�C�9���j���:�1J�8W x��d�Tb�Hm�Dy�yY��߫���Ҧ/����A���U/%g�9�~o�F<�2%�T�������f���x�٪�j�б���`O	�Ij����;٠D ڃw�TB^��g�=�6V��K9h�g�E�r�E7�
�X���;�ԇ�~b?��
*�b�;��d�4MkB&�*�ď����1s��GX���HQ+��dq�1��x:�+'5��=t��2���!�R1 �P8oX�Pa@���mu��Ƅ
o�Y^��m�E�����Z�$�0$4W�6f��
8S��&VCW�W����еQ��_ѽ-�P�}ʳsx3?�+y�)�����$�+q)�N�����cs�Ms�˙ju��sl���o��@5���U�'Loq��Ɋ�z�����'�Ee�� mS���;�G�9�qi�A���@�}��tD�qx}6l��?`*�3�	1+��6^���RwM����N����<�a��_�ڮ>�,)j�x(ΰ�-)o>�=���V*���| k��h"�h�h�*�P��	b؄#)(�e��x�Q����3�ϵ��;	���N���)�g�+%0`w��dH��W�_1�7o�����G&J���A�M���v�L�Kg+�|:d#@<�S�����Ԍ=��s]П�QM�����T/ˢ����r9�_��?�	:�d�$Ba�0�i�U�f�M�1��GUz��Jn�%5�z�Q�6ӥ$�(E �,�Ԧ�mz l�`E�IPL�/kT@$پ^/DxI�ZX<]4�3IhvW��*�)���5
-KZ]�&q!O-D��4�m���{�?ɉ������@�q� ��I���"����t=<6"�]�8B2��+%d��!�w5��dN�쭨݈�j#X��|�u��
CN��Q�*�Ba巋���U��.�Qr���|�dVIzͼ��&@j�"/�� �;$��!�o�Ɯ�(3X��Uq�]lsKV.U�H�(
�*xf��k��΃>�O��΁��jp撲�.���av���l����K�=�,�k"z'�M��U��#�N�8�e+�t[|;�}hV�ʎ��{Nl3�x�	�?����+K���(ߛ���/�YD�[�h��.5§5��uEaI��-�;d���Q�L0eecۼ�2�.�-k^�҂ܑ��B��s�*��J�����e1�G��_��U|����C�!�?��׬x�X��W��oo��:o��"�8,�T=#tJB�m��$�؏S�|\�A������M�-f���`�#E�Q�Q���x(A��o��$�Y3o������� S�G[̼��=O���$3���ayTlb�z��׮1��[��5����~����/��q�_�턂_�os�Eo>�'΃xe�����^�CtJᄚ�3����5�����
��	ߛ�s���j���6P8 �/�`����l�ǰ�	8#��1Vˢ�|*��)�R�g�?�\�(��kC�i�n��#�AM+����l��qEP�BS	:E�I������9������:��dŒ����-Fk$/��M�\���b���u��V|�$�jy������w�Xw��õpCj�\��녷��oÙ:�ɹ1"j��=y�N���_����VaMO�%Ǖ��A�[�r�ߺ��$�b��5�h��ɬ]���^�� L�,��	�rP�� j���R\�������p"�z�j���g�D��������8Z��A��G��r��6��dȑ��6���X���
@Eb�Ў��t'yM��,[���m�*֨3�O糬�f"�Z�����yh'�^R���_�� ����[�|�[QvR�f�w����b�^_\� ����4�s�큵@ƈ�;R�����um_�bhGTɰRb��I�,�Νn�t��|])���ְ���!7�C�FJȖ3�u&����/Qd�� �lQ���H�{�)�/s����|�!@��R%��}7�9�'��/Fj��Z\6*A?�����FuS�ZՐê�N?������u�),�oDk���T�NL|����$�_�4�U�?��M��q�l>Ш{�S�DR��aZ��3Q?��>��/`Ӵ�����{I�$�Z$�<m=��/�=Οc��7�9�K���3]�7��ϏK{GY��tC����{F����+����h4�Ѫ�8��?�.
��w0��1�F>���cҨ@߲��_�P�?���ǾѻL����\.Eqq;ɼ8�i���F�;�R Yb\���^5����vu����'�]�u�GL�dj�̓?�d2��E��.�|�|)������P�9ǿ{Z8@u�{�|d�yD�eWG���*�;ҿ���d������C�X��Ɩ@�;ʽ�G�/Y�=���QO�9���j�Q��M��Z^Z�t����K_��������v�t}�����D����j�����١�{����!����`I��O��aR���$�G8"�U�� �Z�ᤳ�9&���ѩn�'��{͙�U�9l�?�R_���P�ۣ�<���NS�f	 KXX=[-�o�Y����8U�6)�>����	�.�T�s�"�ч^�h|7�3��%xa��钳]d	N!e�'r�U8���0�o�m���>��BxL��av����\euxP�Y���ĉN���~�|3�@���{޸QQMkv�t!���4��S�d1���<.����֓��}��K��z] r��lS�9;��(F7�%�!acɚ���2ex���o�Ϲ7 LwYYTJ���k3�_h��A��N�^Y:GJiOD���te�e0b�2��	�K�Y�f�eQ�ශ��BTw+�p
�n����_�<ٳ�,����F8[���:��e(F���.7i����U���7h oEc��B)�b0�h�)���=��YY�K��O����b.��	��!He�c����)�=� ~yj�@���N�Zb/քN��N�r�12&�ٱ��.`�G������^6�0��m#&��"�lx�k�{�9\:��Ap(��y����_�F_�-ڰ������Yяk�n�3��7�z�X0�e�k~�zEH*�J��r�2���v>���K��6��p����p3�nb�~�����M�,��� 
=����Z��X���ǎ�xǻ2m�&��eַh˼���J)�\�Q(ٱ�s���綰�x~��1�lHiP>�����@}MpH:��Xж��BL�龫�y\3��g�j�*)-��b��@+	�b[�v���IT�ͰI�Df��D@c�ڏL?��;P�Ӽ�)��=?��&+��{vc���gpf��$� $��r���7r��=>�����?��!%��{��/�F�..+��o����I��b�E�嘅~)b,Oa��.#o�le�z{�,���Yb� �U���^>���� η�y8o]e��'�����ǻ�H0�kʷ D�-�|F!��n_x�lQ���m�J���b��U.�u�[*�*ӫ������i:��Da7�HHQJ��/��LJ�`�:v9���A�4k�8ai�d��B�,aX'��o�?d�D�;k|�f�$Q�R־�H�l�>^�Z��w-���E)�q��@&�(�v�='W�>���|Q^|�BG"�����8��;��=��C�Z}�;0���l�[k���w�5j��T��bs�?,��@��-�r�}����v�i'�eP���[��/��,���[7��b9���M�yDw5�Z��^�g�$�ml&�_Kcs s���~�׀# �5
���[���[;D�����1
�v9�UO5�X��4�R	�?JŽ/�t�*�m���v�������qy���T�i�X�O~�ӡȽ��Ac��[�%�J�s��g���EG7S�O�X�X�C<�n난��k0�䬍>�Ӏ".��c��5��'?۝�`>��"�@_���X4Ώ�|��E�+6�!��v�oqZmsg�5�&][�ǝ+��Դ^i�~?>���Y�ȹ�%Q�i��|(�/Sђ��[R�ē?˫_�G׸��Ŕ�Ǥ����4A?�[i��p���9�)��ݢ����b�����A��%o���!����D�/��L�)��w�"�V8"ڵN;Ü̇jŅT���O�8`,���Z�+�t�k�_M��1�)V����� =���h
�����/U8PƤX ��9 Ύ�rܪ/ �fݗ�d{s�U�v��/���qF�&P�;��_��w�]ǣ~�)��j��_OF�Q�f�Dosn�PΉ? ���{v��`vt8�01fQ� UV��:��UQ��Ǫ(6`DNfr��st$2hmQ��vP�K�P�g^߽Hđ��_��+NCq&����1��;>ou!���t]!��0������nҩ�i�����얄.���ӷ�b�GU��!�U\�U��6�u���m�,׫*���KB�A<�/"��d�P�N�|��z�ҊT���<���܌^��꜂d���α��I�L�kc4�%� �'�??���ȯ��Z�:����k�a�d�����_�I1�-�` �V�m�d(�T9#�YLJ�X�]�E�~oqS�Rr�V�m~�2�l��3��Y3٣�����R��ZDqZ\j��,�3�+·�o򘽟\��^~���p�rx�,��Y��eyɘ_eħM�ƟL`�mj��1�M����y4�f)%�q/T�_4�u�I>��fN0Z.Kc1r柭)�	/���H�y�����l��3�jN��@��y;����������tҗ�`h�7q�y�����Y,�!�M�	������W(�s�y�O�$ɳMD���y���	�Ʌ�İ�V5���}F�7�`�e��ˁ��dl�&�׆}�>����b����.���Ᶎ{ϑ�y�q\%H�la��E<ܕ�ߐ��%94�[��K"߉��n�*M�Mֵ���Ji1ذ��{5o�:5��
�ݠT�y,c��\��wg�Z�����B�R~�oܷ�w��*�t�ɖ�r���Zn���c����U�X���*M�A:�3f��K�KܦR��C�<�c~}�D�)5�#��*����%v����	W
�3g��hIޮ�!��2�������}�X��@u��o��k�3�"�|��nP�7�w�/-Q�`�dd�0�5��W�W��_�z��O��I&W:����`����/�1(T�-�Z�2?���}~ax0�ѫ���H��}�U�	^t?�	o���ҫ�>,�_��p`�� _j�#ߙ�����$"�[m���{9�mͅ�f[6���MÚ�zq$���Y~J��:���8G: `t�I�_^��=�����N���zm!>#�L}��nϔW(8�����`L�S۴�Q��f�h��F`��;������;��V^'���[��\�i�6�=�zwzټ���A�@�iD,�u�wCc�Xc_Y��ٻ����.)�_X����W+��vbEq���8��*�ն�y�w��IdK��*d���m�e�GV�'H�o�~�4�^�����o��J �eFl㗳�C�=4���%���J�31�սmU���g�#�^���.�p�/U�C����b[��:�&'�ݳ�*�уT--r��+���'�.]B��Y~w���G��<�c&8�����
�8|�f���f��&�.�N ��I2Ay�w�D )����V�����0�e-�,ܓ/Be���hkz�9�{���q�̖��ג1���{�^�|�-�lS� ��,��s�>���Nd��f�K���fPKX+	:U�,0]/�P@��o����f�)�Ĩ��w;�D�­p8֥��$�����D��uF�F׽~�X��Zl�W�3M�ty��6>���pY�<"YX��UJ� H`�
(Ê�gC	�q�^S<�Z��J�*֗� {/���r����$�uP�"/�V�F6����ɐ�k�����A8�γ��.�wq%fn�G�G�l��]� �����rwzqhM�mD�#Vy�f��\�Uji��I/���ת����6�Ԭ��N"#ŗsp�J�bF�A2N��e����=��g����,e���S�(�$)ezē���<A9D������hVFQP�L����\K���2�3���-�g5�V�*ˈ������2_ust�Ϋ�c���1�,�h
�Zy@�� �����0䔻e�>������fR\n���Y\ˬ�M�b�r�2X+��zn���﬈3W����k�]&ױ�-�ւ0�a�[����8�����}m���^�<��.����@KQO�a�:bT7���l�ЃB\����پ슻�l��"�����~<�5���[��n����|�piT����J?>�Ȥ]�4>Bq�(<�����Xt�ƽ��;Δ��˅�'���d�=$���0Z6	X�QT1�1e)J�u F;��5b������i7�,-��b��%?�4`��S���ۗ�c�Ya��̆>Ñ=�aZ)׫gegL��!�������˓Jj.oN"Q=Y�'»��2 T8jyjs׳a��Y�6�B�_픃�0E�SW�^	m��������̜(�a}D�P��ӊf׻�)	'F��
�"�����Hs֩w��:诏6�$:Z��ϙƯSs	:1;)j���Jy/7�>{ԩJ5�AR��L]"�U��G���.��}kr/�#�Q��(�5�PH�l
�h�&�BF�梽�V=��߬2�P��O.��D~�h�D�$�Q��f]�&*��Q^�*;#��4��R��}H=�B8��
��j4k��=��G΀�X�ye,3� pŦ�OCQ�7'��k���J�1\���N�8�>�,{
D5���(��y0t�� M�90rd^+LIх�s��"���Y�:��;l�d���C؂���L�8�7��p����1d��w �e�$��XI�!�p@���]+6��G�͂��g5o"��T����蒮u�y�X��4���b�Xj�kR��3�ӮTJ�9Q�����ᆇ�0=)���G<X�C����k�Oe[$0�O1��>��5������o���c��}�d�'�+b�v��V�/�%�>Շis����俱�$��$5�͒��:�4����wn�ǎ�ŉ�R�a��Z񆲡�L�f�pIt�A��.z�Rh��(K=�r���	�����������֨�R8س��l���Pت�����_[�G�!+
�6`��K&����P��:,���g�V���U�p�F�C��8Uyo$!�DE��<h�ż�!w�~��K�D���	rF0���:T��Z�A?ї�
������#��(ЀBܲCJ��=�é.~+x��sn!�"N���="
`K���i��t��b��2��l�v���bE�f�x�1����Ʈ��f�-��X���n����b,�xVYbd�D�]��'FFBuŲ�CP&��,���?$�\��i4��K^'Ć�Iܱ�w���lZ ��p��{� j��f֫S���6
ҁ�l�>� �C����R1 �vҔ�u�z�X�TWo�d�K)3?PT갢����ʮ��%Q��+����§a��v��ɸ�C��͆�i)#������/t�^&W�	�A����`����fo��*��-���^LI��|Qv㙻��ͤ���dN=���9�J�7z�J(Yt��B]	Ig�jz�����߈w�o�{�9]I��΋�1�`s�;�)���s���>^3�dhwˬ�/�d��%l�h�/yUq��R�]�Bm�P�
NN)���d�
�G�H�>��ǝ4�.�������>'}�/��p�w9������L��������I�55S��{u1$9�B����a=b�$o�ьe,��Ru�?|���a=�*s�c�ߎ
�gE�̟����n$c�D��@�{0��������t��NiK����L�n��#��v�P��k������6}�"`��&�Ӓ�f��焹@�L���,���G,���°�k�+�λT�}�R���9�
�sM�rG�8:�H��5�Qk�/�rwb�1E�"p��>n�SC��q#;�Kj	�rڵy��J��[ƭ�T�FtA�1�`�����2@���'+9���:��
)�>�����ԪF=�V��2�����©���8kJ����N/�l�ɕ�?���DY����9�O��K�Zÿ�L�;y��j���и�D`��<Kd�
�D���x���x��QF�$	T������p/6�X��ĸ�8=�C�,V���7�
�}|�tߕ$�*8�k�O%v=l�/a����3�k^���S�8=��X��n�(��������1�	�[�p.�u��д��1�)����s���ܩT��t����ʻ���%W�G��;�tuh=�8�[�1�K�YV����k��Ta����}?�Ȇq5� ���3=e�+FB�C�|)(
��|o�xEϛ��2j
�=���l��A�b�[���(dlCG��%�q�i٫��=�ty�={�`uS�en��B&G��E��?��3�|�ߗ6�ϔH=v!�Փ �^*đޓ�;��Te���cS��͉|t��/-��8�_�bOئǜǣ&'pٞ:�@��s��bt��_>ߟ�I���x��9{����]f�{�k�GT)/	-��p�����L>�P᫵�����B`�,I�1�-?g_����A	�3hX/I,��x�<�v���B9~���v!�O\���;2/���0_�~�%���}?`����t�Fp�E8����
��\,�>��1g@>9ŻzgzyLp�-{6p+H=.J�Ϡ��FY)(���D�x`��:ix��E&���޳����2G���G�N�c��\���x�R3��:��<���2�*@��z�5���&���b~m�S�d��[�TݴY���w�8|��g�nޒ���af���kpW�g�
<��W�GOͮ��w���m�_D��tA./}Y����{? cȬ2�1'�>�H��E�����}b�o�sǡ�-X<B<Ou�i_�PϨE����k������,�t����i42�֕�<�������+ʹ 4�SAj�溾�^����p�s)��P�s�P�j�S�Ϗ���ERn>�����!s��x�����ND䌂p���������2�����!N&�_��yLpL�u�'�gi/�'<f �3��\}Ud����o��ԍ^����Ǵ;(���N�a{�S��@��<���	sV�@�(�,j��r������]�:@��1�;O.�{:��Ea�O��^�ޥ=��9d�7z�V8-��t�&��� �)��E��c�i&�~)i%x��|[�<}�(��� 0�W$���);8��A������3H�Q�F��08p�ތo�M%PYh�D��W��g������e$�ϵ@�FN�P}�Tp����!PJi@�|N�Dsď��>tgS�c=$ՖK�-��K���2l�r�t�A��e��=6���"�:2{��K��G��C7T��r4Q��:���C���SW;'%h��=�ƏK�Hl,��ɫ2/:֗ײoC-x�y<0��:"����S����0�5>Y!�Z�5�k�[�s�nt0���o��\�
u�3�o�j1��~/B�rE�}-�i6�2�@�uη��m:ϥ?����'�\E����H.�粖�\r]�;2�]@.��@���.�N �6A���:�>�O�M~��A�\���	��gɴ���M��v��`�3���UJ	��c����)���8����h�m;��q����4vڑU�g.�ӨM�m~0��D�~]��PA|qR�M�q�-o�M��:��u1�+|5�e������ד]���C}j���N8�yDm�#�y״A��MIᤱ�� {fP����{k��$��|p�12~w���.dDr��2���W�����;������)��qt���R;�����0�����G�(��]��v�>����[����dCp����¯���8x��z.���|���#��W&�����Z<4-��
f`!l�h��g����t_m�u���
Uz��K+:9IMU�6E��L�+�oN�/��_���V���H�ѥ�P	Q�C���/G�nN��C�m{J��%��N��և�%��C���jrߊ�G��ýP+l?�joģ;�,S��Q1�_[ �Y}n&r�^\�D���wT.�; �T�`(&����s����=�hB6�=V�0x-������Źb�HP��c�s�֜<1���4���6a�׫�(�}�%�g������2��7�̡�%3Dw�X%�D�q7?�%�;z{Ү�����ە����|�����H��B-�w9'�ϝ=�݆�o����� _T���B��f�0X��hw[&`�~�-��3�ұ�R��D�[�d�ދ�p����2��_�ȹm��;p#�y���Pb�Nw$8����jd��J>��g�t��'bE�^.��G��6���̍E�lU��y�}��ꪟ ɞ�K^�ϛ��p�+� �fd�X��G�>��y��_��/r��u�~�K�H+�A��R7 �<�������(db�zN�F�?�>�¢:yj��D�o�A�3_�����B8�b�:/��{�c�_�3^�W��Yl���:�(���b������:��V� Ý+�'��Wif� S$ѿ�C�ї�\s���b��n.����"H2�R=X�$������;E֊v���Bo&Yu,����/��� j�I k���P+V�J���;�s)�l�#
K"ˌa�,Iz�N�����Gh���wn�&���B�`���+e�%$��q
7y�G��*�;�:G�d��vr�}`������ۅKg��>e�8�����O�_�#KQA̐B)��e�� y.ڠ'$���.�<o&�n-cd��c#���U�m}��s��C���F{��  :�ߨ�\ݻ�����쨡A�k��i��w/�`��ܛ�ߍϫ.ۇ��F�mX����Y�6�(���x�[�8\��������cO�m�H��/�3�tsQ&�>����@�Y*�>Cp'�>YB.;r�R>�<���sn9���W`=G�h#�L^k642r�e6��g�I?JA0��6&����9Ɲ�9�p�Qߍ\�j�4+�QW�|V�N�Dj���#��1�]'s&Bk�6]�2�>_J�_�d2�����ɱ�i&k�� �.����3��L�DW;�XՃ`��a��t"8
�&�-��r��� 7W��֗鉰��U�X�~F���6��@�q^����9b���l���Ћ��
�}X����;7�+�p!�#����Rֱ� �0�C������!"m�V`#�~wBɜb���O%Z��E"��9���?�G_|����is��i�"�jCh�7�XΑ3U����q
��d]�Zp�K���ݮ6��9Z�Ǳ��8�<�����<�� ���ꜰ�g&�K�.�����Wu(@a��'3�����/Y�^�L0"���d�i�o��+!5X�z���`h��*�X'�����<6ּ-�k�Bw��F��}�r\p��w^*��8�iH%��Η�	Ӿj�tyz��+!��zZl���}JX����E3�z��3˕��$�y����sB��e�(�a���V�N� �]�\�����Z�(��O4i�K�8�0� )j8`[FJ�����Qx�MO�J���@����"�~RuH�EtB~c{L!RMiIO��я�f�k�c���e�Z:]/m�=S84��v��Hߣ'[�����/+d�m$���`
/���LǶ�m�Ut�����v:�a�*�ށ����v(����	�0���E��U����* -�s�S�+Y�9U�6ǋ�ŀ[�Q{� �,�����=���n����\xc�WRPM/���SF�w:N+#z4p��g��L�{tA��1�"!D�l�X��?�ʃ�t�z� ���;���	rW_���(���*�(5�t��*����l81�mٱ��!�G�#��њ�X9���D���\�]�ޖ�Kt5��b*-PH4
�P�L�v������o��U����l��o���2�%������ ��̋����T�)<�V�H�]������NV|r��2�
߹�e�ذG�^���T�I�@�A�&����C���xA�<�8�֝�処��aj?�zL����"�(x;�Lx�H����sU�$���t�$OF!OЕ1/� �w���%|m:�ۮ)��6o�!�J�'
�y��,+k1�b�^�aӆ`G#b��w{��������	��
��$s�0��.u}�z��y�wP�q~�roVՙc�.̭x2��p:+�4�8G�D���U�h\�gn�N�Sld?:�����;�#�A��C���R�#t�^sm��*m_IDn+�%�x$Z2�5gh���CJ2P�ܨ�S��j&o��<<��$��4��É}�Ύ��b2#8qzQP'^��>>�M�}�X�x訢�I�O��ytK����զ=)�-�k���|�!������]��g�(mn@���r�Kl��eY��9$��t���o�f�_����8X�at���#��,�D�v�-�'4���Q֍��v�7b9|B���	KB��\��K�Ѥ�N��ۛ � Y����ә���>eoa��Ёd$}K��V �|���%xi�!�����y�A%]����V�k����3,�#~�I��(Bt�L6/� �	cE0?�l?�k!N�`�����i��G�TI@jE�������lCESƔ9�H�#K�R��X+o"���놦;|��^�b��C�Ne<�`R�ĊK�3�H��Ԡ����K߹��TZb��r����Ҡ�ʥg�F<'o�JӬUؕ�P)��zÍ`������3C��,g�MQ�Ϸ�L"]�`�F>AF�=L:dah��o��6��A�X�=Ν��%x�Ǳ@����
�%��|�;Fu���8v|;�.B���A<��i�ջ�+e |e-�C5k�Pgp�n�t�#�n���{�3��������ߣ�ve͵D~��M��i�
����� o�)Fq)cb��>hv@$��l^b�s1��=eb���ʑ��e3��d3��J(��A��+��\����}X_hG��aBz�Z��,�P�T ���m��}�Y�v��G�)w��#�ݵ�>!�c�$�0KkF%g�����������fi#��U���.�48	�m��{��:m:���%L�S���	ėb�_C��i0!��>K�NA���wrǷ`�s���{ʉ�7�K�x� s�7$C�c���*�wG+_�-[� /y��~�K���q�S���z��6-"��3�Q�G��Rs	O�t��L�^��"��ߺ{0���m�H[�Sj��+�����]^����R��:X���@*<Q	��˾)gf5K�!S?�W֓A%^��~�	Q�ś�"F=H0���'�����
`����D�Ҥ��̱cvQ����;�@�܅�_�m8{׾�1�=�2�};N��k�B�B$�.��:%�I���Z�ӡTN�.�<0���ݹ��ˈw�xT.Qum�x�l��ٯ�L�_��/&��t���m�2VߚR��h�)�ᄻ5s�[��b��]�F��������W��S�{J(�`�3#�'I��&�A(�
/W�_�b];cfѫ�^�����&ɋ*t�6�r���z��7���ԃ������B �X���µ��.�0�_'����|�Z�\^h�4>�4d�
���z��*'q��7�A�L���O����<����1��8[�:�1�i+����g��q�T�)�rj���$�J�}f���6N'���|UW�P�}�
�=�
O�8��kD�}�_F�U���\�i#FBZ��9�"��p )�@�I�����৮�ʹ��$N?W;+(yL�kZ�ЬN�ҋ�%[���ݚjiH�c��1.�/҃sI%����\����_��ϯ�2�/�)(�y��R1��]�~�P���?��"h��1G��o�ExoHQ{M��F�;��M�F�J�0��zn�3����P����r��@{�5�Jz���ʇ�s9G�����_�,@n�:ǉ��kX.��Z��?�4rn���C�t��]�]1o�R}T�Ω~2�.�=�h
�����j��6?�����G�wlp�ݹx['�c�&��U:P�N,�"�G�O�� C�V"w��{��9�8�,~�*�y��}�t���RY.��2�&�j1�度���DY��ՠ2��bL6 ��`L�`ubx�ߒ(��i��9�K��6L*���Byo�9�";¤��듖�����y2=��r��Ya�qw��^J@�H\���taT�e_r�Rô/!}��U<8~Ͼ���,�����������������k⤰���I�\���5���;�r�P3�����a���
�$�?�:[�4����Q����
�<�V�2�b㍶~f��<'�y�����]ЪOݫ��cy�I�7D�w�nLY�mNϚ�(ME�Hr1U�	x�כ ��-`����V���)���0���������!���	 kbփ�d�_�����^�>O�޸m���^���K������'0�ʑ %yu~X�&�����:Bjf��a��u:�?������N�+�?�Iqp@6o��jP�I,LWԺ��'8��_�P^�00c<�X�呟̝H0ؾ�3�H��Z֥��0�c2 ߔu�ۗ�-��$��������2S�k��g�t�#'�ٽ\㈝�,L�
��I�]�F߃en�r�3�>1\=����a�Q�E4藚ė�ԉ�̩=p�5�V ��i�a�(�+�H8U��m{ܕCH����|��ݡ�\C ���!;P��*�V��
�ņ)���M��Kϡ-}s����;������1B�&NR�cw㱍�y����oKüg��	�t�kM�xp�>|X� �x��I�.�YI�1r|����D
��GA�e;I�!7�|���2d�����HX��8�O�UocȮ7�]�pS�pB��S���9V�M���%VN�t_�re�a�N"T9� �<U��_���4��m�5XU��.N��&�����4�G����]����R���/~��o��1��ba����]+X\��j�)����p�h��@ ���^��[6>���h+fl6+L�.�������h�G�]Y��qY����φ���A�G�^?W�Z,�����X!7hyŘ+�?4�t�,�ر��-&g�e�Y�-�6�v uG��U	SZ�~X�F�&��}�k��P��)�DXPd��Mݟ��ݎ!���_d�d��d=_w�sM��:���:������ʪ;V��ޘ���l��L�g�kd)5\yz���vzI�mk�J��T��䢓a�*�@i�;x��V.��D�L.���I,��-���aU�a�������/��q���� ��5:}^p`���ډ����Ф�	z��"��#c�N𓚺1�m�*[I/��5RК��b8�j�l1:��x2����k9��P,0���bІ�^-F=�S�#� ��w��*��w�ǭZ߼���_q$Q�7,93�9��(le��Ҧ��iZ���:<G�{�?ׅ�G�'�tÞ��m"%c�g9g�� W������p�ӦQ�rچ�ҿ��,Gh+^�W7�K��=
��A�!k�6q���3g"���u$��|�%�����B�
��G*^=2尪�H'���יX�P�ID�\.ӋK%q���/`�!.~��;O\���T�I�D�ي�B�w�k���{��[#���<QT?Zq���vS��g�O��o����j�����p�r,����dǟ*��;�=D��z<�ha�T/��q0'N~#�u;�%A��8�E>-H��R��:���>3��.g
��AW�8�n�7mP�̤��ť��L��=� mS���/&5��D�"�Ob �G��{lg�G�*���K�s���_q����#5`�# �OЕm|�����%��!����K}G�)���k�A��8����J 2s�`KD�; 9w�k��%V���+�NzV��[�ɩy�o�	W_�O;�X>�(��R�d�f���܇�$�3��{�]����^�N�-���u/�kI��������}�A9�i\'�U!'V�6dꬬ�闯� i�U��}֧B��\���&s�6�^�`��^��ma��-R �װد�晝��K��\��X쫩V��K#�_I�R�u�-ґɲع8;�����? v�V���YW+��]�jd gq�ü6_����yx��^v�
�B���q��*�#<�
����;�����]t/*P!ޑ�� ���Pb�y��+�8 )U�s����n�1]nP�'TΚ���u90|�������_D*V�80��e胄Ǟ��f򰫽�@Iv��KbG��rM �;�UF�t���*�qa7�=Q�qU֒���4ht�V�W��ＦӰW�H�[/A��!�΀N��68����k$��\egu#�F��L�}�tV�q�`��N��M���������Sw�x��+�$a�u�~�蛯��ڥ��w�.�l|3��FH���֙�8�1Ъ?~W/ m���ҐE�cE���J���Lf�	O$YaE
��v+K����cQ�'a��ms1Z�.�,�r�||�`gB�8K�G�����:An��@�%ݞRה�h����-��a(� �����|�d1&��#߮�[lb���RP�I�S_)j)����fAd��fb�ޏZ�нٞt��� e!3���Z��d�?�O��̉����c�̈́���R��*L��+兪�82��}(���ԫǹ��z���Q#[����)Uh��|ѣ��ى1_8��]�x�t�x��t9�>~5��C1������؆TI�
�7�)�P��Q��·S���P�d���s���0)>v9O���V�:���>5W�ޱ'�����¾���V�������ޥ�ϒ8�W.Tp_^�ͨf<���4���|�,����x����)���+:���j��ZM�,կ.F�ޥ����0�Xy0c�-���Ғca�۪B�]��&IA�m���w�H�>D�🞣�poHR�&
t�m'��"�=�UELL�$|���k�P4��R:�#o�h�SBW!4����ˍ�@�l�*�D0o�W��`<a�(��om�z�_߀~�t�����Q,Am��k[_�Su}Q~ɐ-�e�@>�Cf�=�Dǫ�۔�����Ϫ�� ��f;�o�
�qjj<���^OQ'�6������[�N��ng�#y$�{�BFEU!��_��a֩/�W��`�E�3o�P}ldd��qW.���(kB��`�8@�����w��,"�⍺�-OϦ^K��/�ƅ���^�a*�F�R���./��8h�������(R�44	��#��aWF�f�t#e����o���)�������c*�||����(�v'n~ڄʠ��m1k�fY�R����]�,~����J��;�_~�P��ƇG����v'�_��Z|3�-���[@@`
xp�M�ǣ�b6�$J����v)���v��r��Y'%�*K����>_| �(��e+i���ew�a:+��'5���tq7Gm�:@��W���l$�3� _VL��/�o���]jU�n�[Ɲ��6<QуP�4�i՗�C�T6�h.j����U_6Uf:��/+۴[uu#���^Δ�튍�ٝ�y�xRT���|�Y�.�sT�l�����G�A)���WD�BN���xs�	�C���#��4���/�l3���_�!(�)��e`\2E�3y_1��i�w&C"VY�(��P3M��;�����1p��w��m~I���c���UMh$� ��t�;z�}Ѻ2�4Jê	���������ѧ������Ǖf����nN��2�[=�L�E����U���
���<#.3|��6wt���3���0�eX��H�%�om6�̗�T9�!�-�4��`[b� ��������������o���� ���牝��?�o2������'Y��8s�L~�mH���9��R{5P-�:ʱq)+�*�Bm�Yq�t��¨1{�~���Fe�نu�����E���WI��8ʒ+��jC���Cw+�ނZ1�Q��e�a�,N�T> ���:g��e�#3�)ǃʶ(�Yξev�90����A��^�V��l)�
���J���Ɍ|���W��p�L�<���?|V�#G�+3�hܨr<y���Q����Y)p�^��wO���2�I�B�t)o0:���򫣽���xV\��q��)�8:�v��| «@չ�T���NV~+�������<�d�Z�����-VJ�%�{c%I�޷��-�@j����"))(�6d�EE��h@��S���n2��:z~�Xz����ab���
�?�R��]R;.c��)>J�%�*�D�B
z ��>ޭ�VFꢏ�zL�툱.��麸[�� 3:f���NY���?`�r�
���t��Ӣ&��-{���]�2X}3j����w86�$z��s�ۨƠ%�/���y.U���d\mw����a��`�$ 1�p^U���a�4_�7�"�����E:�yY��ZL��Q���i<���X�~%4^��cA��Fp�]JC�W�q�-�q�^��;K@�e/dV�o�8�c0	,{�Ll��d�� �1w���8�0W넍���9̨�wg��y����b�����|D ?7,:�{�w�-&����g��~?����TxI�{��%�L��LM�N4"�l�fr��g����(6�s��������HE�ݸ�J�#�T���f���m�+���y���9�7P$M΀p�{���HU�`U���|?�M��Ec1׌[��S�8�5�@�?�m�c���LuF���O����@_����=>���Ǻv�ܞm7�^�`�{'��^�+F
";��/2�����*z"6	�̤JZ+�8����������Y�q�oҍd�?�w�c���-d�:��L[���2���l��9%�Bӿ�H�aŪ�v�1�]�RZh}�fF�׉(,�0�IیA�()�m\��Z(	y!�}I�w�����4i-��{,�\�#��>�j0�1���>]���h�rX�G&����lWh�~�D�����ٝ���� � �#�d+x�^���뜿VX�������d���7��y>65�@�!,���A�Dy7pAFf&��ׅT��i%ə8��:+��(�7����Ů�"��m��:Ԇ##��,ub�|�Έ��A��B���fk�*W��Ţ𒣧/v(	�O4���2!�����wm���a	��F��kf�/��
F���4t�����0=��~�_&ȿ,\H���_mC K!f�V�*z�����*�1t���F̧�-�4�F�뚽�
𘿃����A�2� �x���xO�~�.�D���O�ɖ�{�9�C�5�w`�mj۔��Ma]�t�]\l������FA�& �7�V���U`�>���}���|쨩A/܋82���&��� �� ��)����n<ڄ��Q��I�V�+}T�S�^�1c	E���U�Wd��@E�ԉ��P��e�%J3L���RT2��q�s�H˽,NƖ6��x��>��f$6��qdq��F3�<x8v���`լ����2Z���* ѽ��vt�vg�����ׯ��Q���`�A�#�E���Y��S-��[bAEέ�}B}�p��������2t�<��Y�r���14�ON��(��]�s	�1jd����'���*���ĳc���[�x>��u��@�Qțb.���Z�ة�#��n޺L�
�	�8z���nG�����L�b����ꑩ��r�S#j�ÙQ�׹MD���^�Q��S�&GF�C��e��ʓE䄸צ<�ed�$���#�f�ZI���8:y��`i�3�v�oE��Y��q�Y�~�;h�:�����R��6����Pk<�6�V3c��;����ЅP#�?�$�[���Fq9���P1���� �y�N0�IR�V�Ѭ��B���|4-Q{�*����=}��:��.�+8�,�-����;�#EX�@붔��,v����%��wc�Z�K�ܔJ`�(L��N��<�Y".�?��4������G������'�C���4�,�jRr*�%o���G� L���JQ�=
��\�Q,^"-�%���D��0x�D�]�[�Z׎埩|݀ՕW���2,n��X/
�\;��L9)��w�yIo1�Q�����L�Ěb�G[ЬH�h\h!E�L�CT�����/G#~O_k����&k��e�h�.PW"�i�������$�;�X��~x��m���)��᭻���m����gf�3T�Bm�E���C�:}�ǿx3���]��O(O/d(1�FD!�(������,	�>�]�:w��}=&P����blV8L��2�k\�p��Q%�ZEc�5����-SH���1�1�Ǎ��t��aS/P�t��,%xt�=�ޢ83(��<�|��#t�u���wP2�>ֽмca���:0sR�`�|f���x����ƙX:@���v��3����T�g����y�����M;
]�`�ݭ��fl��$&e�g�ž����k ��Q�k�am2�mY��W$u��b�a��^<�<��L�B�3A�*���Z�K�wG�G��>Ia$�A/����9��g%Ѹc�W+��88sL�:D����bTb��X�r5�c�=�~�K�2F�^�W7���bC��]��Z�#�]���x�	A�2C�����M6�yН&�p��T����t�y4t�bފQ�*�$	��=��KE�}(|Y`E'�QUv�`���c�r�<j�)����;�k�]�@�l��S���L�}�U&Ʊ���k ���g�����x���㑹
(���w�s�����.�n�� W��C�?�H�M4��o�I/�s?�ᨥ������i���x�d#��x�Q���?�0 �6_�b������=��/'x���4���~EU�.�� b_���;��տLY)�0����$X�T���I$�'�1w��O9CkZ�yJ�1�٘�:����1q�Qwᣃ\c�Do�<he����	�ݛ\��>n���Lí��B�/�p�r:U�Gi�\�(DB#O�l�����K�ܠJ�r	���zF��9���a����]�[늭��'�aOؾ�4�Q}�aM�X�vC3�<���^܂5� ��5j��ƷD�OXh�g��ڮx��mc,�:)v"�-��h���)�~1�v�$2x>yb"h����u\i�r:sf��B����R���Eyؔ��z
��a}��;9��fepI©�]X�+������.zl�ۈ���D�`@I9t,�G�{�<�����c�%�!󥔭�k�=#���D���t��"K�j�ØŇK��e�q��h�v�]΋���4�N�3�+���έ	צ��[�
�k�}7�����Uy�� ���v'	�eS�r�tQ{
�Ҿ�	������)��cKS9B-�h�ϼ��_�����&uA�f�];�Xѕ�xM��x^E�xߏ����&w�,��Y-��˫�}��ެ���'%��n�`�+zB��̩yjC$�5v\�x�ٱ��;y���f^��YQ��A�c�����%u��O��@��!���۟�T+ȍ� ls�Uǯ#o�9������b�[�j��u��gi�Dq{,�gG^���Vo0��h��*8f=�g��͆&�|��?_ҀPyxة�eoO,WmF�k���_o�:~_)��gF<k�����)�3�ݶĹ4@�X6�l4m���|���Hazd�{RT����=����O:�訤2k�S͔Z�]�����E�&�����Pc�}�mjȿ���oɟ��ѩ���ϫ�����6ƱXY�Ý�}vf"%�c�g'�Ls_7�n�d"^�I�I���WK���4\K�	�уt�_�V^��o��EZ@�S&�&0ǁK�[L�@�/�B��z��rR3iܘz�4I��<"��?��y�+=&qSPq�>�rѩF�(X\��K��ԋ=q�O�<df,2kc����H���j��"-�^�>��/��gR@�~n���K�AE4��8�p��i��X�����W#ψ-x�����ϩ��D��C��4xI����i���ظ�y�U��m��$uU&}�H�b?� ���X !F�l%�w+�`�()!��֜�<��&]H9G;_S�UA�q#��Q2W��(�Gҡ�EW�L�]��.�3=�-d�Hpu�Ω.��+El7�9�Sy6��Dd|3 ����D�|ѡ�B ��ҷ[օ���auh�+���4+P0k�lO��L[���0V�Dvgl��n���u&�@};]/'�SW��wt|�JL��U�zH��4�˅򤙕ހ�D	V��5D�ϳU�Ȳ!�E��.T���%ZfP	��,�t�G<�Ij)2������S7H�6ނs���.=���f*��Czĺ���\؃ri�}��qL�|���f`�����sWs�@b���t�[�l��_\�k��zS���+e�E0���'={s� @�ш�|߻��H�$#8C駸�w����뀼��(�{� ���2�dS�b���� G�V�D�T��ں�(��믟�/�QS��q�����O�]v`2���a��N�����$`}��A�ZA�#�W�ƴu������w���� NȎ�0h��ӄ�5�^�/̵ڼ
Å�v9%�Hl�}9�>���� oH(	�Eeß#w�U���&|��A���|j.���oxz̜i�5ik�b�{lE��C�7.aV9����ԯF�ȓ}�ݤP!'���"�8�bݐ19[���ؗ�EW����ٖm�R�_7WD.qc:�_h��{ÐG+���������x1��J��?��Y Gm	?`.�1W�C�Y�1�ҫ���Q�b0�B��|{��($�'�8��E�$�vG8�@[8)�w�=U�Ej���:NX�yJv�O; ��-:��"30iO�A�_Ll6��9^� �ل��o�����7�ql�F�����A���AqW���oMyץ�k��w��TX�UT �e3M��=�8�#�x �o�-X��p��J���-�p�4	�X��[#�ĕ������9�w�/�na��
�;�	���Oak�QV��Y��~�����/�O��e�i��6�`�t��F$+R���jPn�Gb���K��[
��^�HZ����K��e�8U�d!xE��ƌz�Mz��.y�+�wH�y���\`~W�d�x�k���l`��CB�a��ooIHB!+G��\"09�W�B	뒫�s ��J��Ԛ�^�}��v2.�| �wM�΃�~3��j<ߑkz:��!e�d��rͿ�w`�(S�N�`��ҽU������ZHp64�+��m�Y���h�ϬN<�?y',�lRZ5Q������~�cxŜA0���W�d���U,��j͇jP�%r[�̡��t�j=���m�BܹT��o��#�L�h>��S���PO �g�Wn����Q�:,0��;�)�����a8�#v��a�%i����*�a{��KȰ��,�I�|u�t���O�;��J>Y�s���}C� �62�4��I��U/(�YΙ�6�>*��w�r=k�79��Nd�M��Rr ��=>3�_2����)):����o����kKa�����W�5@2�!׌dM�6���[Fd7���l�p����߶�����:��)莰*�1(Em��M�c�����"�3J�r���
�'�U)�M��c�������%.�-�xRo�qT�ߒ����ۿri�*�V��5gΟO�Đ���������a������~C�a�
`+�\0,id��{�[����� !Ty!?1�fQ@���>�dFlF����l����c}�ӱ��Bl*Ӵ--�'�����ǃy�"ˏ��4�D��56�Q�����V��Nr��������r8.=�?m��
w����L!H�-�pOD]�}`�v�&Vՙ-����^,>H4Ii�ė�s(�������d�+�L�EiD^8�4r�݉�?}t��VE��-��%��WI��N���1�ăK/z���0�*�&�F]`*tk��0�6���l/���j�YF����w��.�`���&�r��z 6�m���=ۗ�;����@?�90Hάkd����xL9���+;)8�'Y�9)̾&�����R���KvNd���@dk����1r�������̒��J�h�}��,�=Yٔ7��s)W��e�ϖ���)e�=�g�ꗸ� �P����˖S��"�t]���|���Cb��_v�/}���D��m�����_�k���H���J(���C������+f�$��J��C��\������Gٷ�p+%�l��+��y@�hO�i��2�l��O����֤��Q�6Hٗ�͘��+�C�"�8�Aқ`�4^�t�#���Dw?��
��4�_���s��#�2�6q�����ʃA�>��*���8����� �zTI��pf�:��k��l?oř�>;%�*�,+57��[�nho�����%"��_X<���l 
qT ����~~�wW)�Y��A{ b��ƪ?�(m�D�\�y`q�/lq=�+�c�:�-iѡJHQ��Xc�9O	�h�) Y�4�F�$5��)K�V���ř�e�'�D��'�ȵ�?f1�k�?�-y������L����
��+�T�=�����i� �O��9�Yw��r���.�7d.�G�r��]�R��߉�������'�A�~ɡ�u���^��d��u���P֊�c0� �>�O%n�M֡��O�M+�����uB���3s��G��v+'����'�A�c��tuk4ӯk�ھ�Զ~���ǣ�\���J�	��[��S��ޝ��)v���� �Ǝ��2ͳ��j�~M�MF�t�N=7�O������]�M'dV4�T�D]H2t��:R�����:�)�/���f^؂���hy�*	��x���U:�a��](�yZ��b�Ǥ�Q��*Q��38k��Z���_��($����^��N�΂��-��u-��Pb�$q����`O�n��ԣ�s`�Ҵ�u�G*��M����0k������Ӟ׶ۼe���.5�u��V�ٕ��Y��v�7xhj�O]�U�Mg�!٧��1�@��F߭7z`o�{�}JHlN��>��+���ТF-�.��.�O:J ��B Vv-q�)�+��͖��Q�W���ܬ�b�|���T�VhX�hƥe��U����5�?��*���<���(�-����"��r�"� u��Uc:)#F��\&�F�*����3%w�(`�3.3� ����N�v����E�d[��]P�A�Ʋ�n^��|n<�2m�І9�:m)�d'tY��K���YíƱV���,�Sȗ�?���Q�K��'.�ø�r4�F���GT4ђ^�@1�'ƈ������f�_~:t�{��M�
�I!}7��Qko畬N0#��^�u#�?��2��,=���H���Gj�mz��o�r������H��vTrԼ��Σ͹+�!����	��V�Y����H,QT��BO?�G+��=�\����v�8����y�] ����7�d���VR��r��)���턼ĳOA^����0�1�j,C��.����͵�/!��XRss�é�XRљ�����ո,�p�	������.7����)�\Ȏٟ6°k+i�:��A|(#�z���g��ՇC�aj�*���Ճ�!�w~��44|�sς��^�&'�כ�|��3��.{?�`l*P�EE,,"�<)��Ͷ�> GT	'�/�Ȇ�π=�j��q��CoU�k�՝�tޠt�n����l�%�P۞k>;Jtk^i$>�AN����%<3�/��N6��L����D�$W/�s�8�_�13<17��og}�Ͽ���A�_����_�6�OB�j.=����À`�V�O��g,5���Pk��{11�p��I{��0a{���-��.8܈N�-ؽ�av�AL�GԚ�#T��Ιk��Ց1:�԰�������߂�}�o���?��X������u����:�N�5�Г����1//Y�ɧj��P_!>0���u+E������ё��tʆ8H�d���kq/�Q"v���az��鱼���O�n|���<��w`<��MJ�@�'�*�Cn���勉g�vʞ��l#�5�$���'%�RE:��Yt�Q����{;]���B�����܃LĘ�\`
��
ɇ�X�w&�4��17a�t#�����G�(�?tƱP�/Fpd�8���y�af�V�%��a�1D�C�rշ`b�u��L��~7V��S�Ċ�ﲨ�j��]�$b8���6D�J�l�K�`�w������ˉ�-Q�#��g�� ��.%󉥗屷ۺ�ǆ��s	ͰU�3h�+TS��͏S늵Ρ1ڬ��T_\�К�*���-q]��}�r�F�+q�y�����}����E�4GL7%��@��M���?�Z�ݖvL�f"ZC�QX���ُ�`P�"UC��bk�><�jRZ<e��煎���מ��<�͟����ŝ�	=6���>#2�j>]��pe�[�=���M�U�T2$r�w'wѮX��9�;a�/�d�F�@��Ů<���/\�k�0���#�� ����,dܢ�ʶ����ѯ���O�R��gR=�����*���d���`0;�/����R�m��ɿOQ,�
,�G��O-������=�#��@�|c�o�z���X.��o�r|�F���i��Y�S�X��T�I����]�-��X������Ԉ/�ۃ�*�⼦f�=X� ��:`s\0<��ԍ�z�A�Lإ���`3Kej��GUM8���$�D�uj�;��Jb�7�"�b3�BwxT�]dsI�����C�|3����:�e棪֝�RA�)Ѝ����_A3+Z�˽D�㒥�y��/C�~N����T�䣣%C��\X�)�'LYaU�~Z0�;/{��v��{��q.n�}����ĿW���i�٣Ӌ^���ן� 4��܂�]%��������wmWV�#p�G� x���I���(/�R�)�{�t����$I��`x>Ҫ���xY<g�=�%�y�ShE���âZ�ߘ���d)�`=�Gj�$<�q&�<-�D �#7������ƨ�;Ɂ�lT���L�"k���(E�g�v.����n��}C����p��[E⩉w����37�E�4��aN�0�[a�_��
M�Z-"���6n�h�8�GNb�Ћ3��A� u�P�XCZ �/���n�U[��黋zĳ/Z01�ڔ�⿭sR��zF�W�]�-��M	��S8K��X#m���v��s����\�E�$ոsa��D��{t�Fֻ���3�`�n_ƶ5cW`AEA�R���2���@V���a^����N����#cok��m��`���f��i{���f�C�_	&Fy$�M�HG"��)�\��ټ������k��>�B�@ 193��nn%	��� va7��?`Wt�<��w�)�=iڊ?/�d�m�+�����dvcS�I���#T�#v(��Rb�G���A���ٌ^��v���4���P�/Z/Z�k�3���,���1"�|-��os0��=��R�'�Γ���2���v}j�T a)�2��	,�VL�C��?���u��IG}t����P��<![F�4��f*���įf�i�D�jJzo���*m{X��� �v������Ǯk�9�}��H�J��_`BY�%��Xc���J%Ȃ �g�q /�g�໺j^��%HG�EƱ^8t�(���IʍC��%��&�[&������s�X�����̞x�_�����\]j�택#�FQ'{O5�߽�7B+�F�(���ن����g,.��L�U�$�,��Y�&,�����'�a3�l���r?dq��/�ނ6��6�7K��$V~�:��b�*�*g�10r����btS�tEzD��<Q���^P��C����GN�q�(c.�}��JE�a@�IBheA�z^�`�W�]�ʨE8����'�)�z����\�<�s��������y��C��A[H������x�EU���6ܞ�ݪ㵖��!���I�1�U��|���f�.�&��w%�gL��^o�,:]��d�ٌ{��as9�V*Iv��e�e;rt�>}c�������/_�.�_��9���b�����q1pQ܄)��j[+.���k�U���BKT-��ʛ_M���)Bd�ĝjH�ܐC�V-C+T��C�����W�b��e��$��T �Ϣ����Op�:M�suu�]a��B4Ȱ�J�}�Յ!�ex������ᅭ�|����R�U�� ���
�J��B�������n$Y��T�;�t���^�];��N�p��al��dU��Doi��H<4�B���
B��~�#�@Q-R�xk�E.�8Ѡ/F��؏]���`w�����˭�<��m,��Ь2s���#p�m�}��3$� ([[qTm�ms��Ѱ�����Ԡ�����p�u�l��W���Ym��s�T�3 �%��j�<��\�"���>��#��^"!^/<�?��S�)�u#�s������qKO���7���q�6_��ޱJv�d��W�%z?�%�TH8U���H�f�bdBI<�n�������&�fe�`�-�nAk�!�!��u�Ӝ��m��K�c�E�L�'�`�D8�Ge�	ee!'Md D�R�#Pk�L�}׃�X�ɏׇh���t��3�Lqq��̯�Y����(��n:�,�eU�U�&���=Z?�j����>��駕�w`�^���,r��l����s��;Z�d���?o�W`���á��)HoJ���~[����l�|j�to�-��afOK�N�i�^��GB��(#�4�)l��?p T��J���Gk�61v{�B��T���#fJ<���JB�F��W\L�J�;��%�5�ɏiǿ�jQ9s��pz�v8�խl����˵�v��(ym���Kx�rĦ�̶�%.RY��%3��$���t$�~ʭ���/]{I���(?3>s�l�A.s��'.څA1�&�by��X�w��&b��q�}o]�e�����V�dJ��`��۪�T�R�غ���$�+�~c=7��f])��tn'�Y�w��8���<s�Bf�ŷ�]�Ch�g���_/w�x;I@h�&y���>���z7���kl4�b)m[�5����U͸'��wY.����ҒS�
i��C~|t�/�!�l��F|��b����o�83���W���gbM�|j���E���+�f�!�6�f�Ey:-�`�h�;�~]��긠�g��Tצ�1譞Z����/T(n�찢Z+��-8� ��Ifi�FQ��H4��a��nu������V`u�Vj��s�j^�@��S�H�j���Wp۾���^C]�Qq�-W]J%�wU�7�1�)��'��ݷ�E}�O����t9�����[�G�e+! �a�s�F�qQݹ�hI�2B&/M�7�%_��X�+��uP��i�+ϊ���&G���=e5c�z��5�]Iqh�u��H��~>]���8M�G:�ʜ�4�,P��N&5x�Z�U���9�v�S��zr��B��xߛ���.���;�9���>b�����Q	���rg���4��V��~1��`�G{��hq.Uȳ�ID��0,���m�<�@)��ya����[��SPA{�2����]j8��ցiH�,�Q�f�D��WH�C �g�G&s��la��I/�~�$���S�V�>m��	byJ'h�{�~��� ��U����P~�~���0�8>W�'B,d���xO�2�3,E��8�mS��q2}NX��0�!c,�xr�����'imIe�0��x����sI6�#�����Zۖ��'�ؖ�0[�ꑓ*��B+��1����l��=챗��c�3�:
<�)p�l ���)!��M��)%�M���Wp��@h�V���A�=��WU�~%���Yu�Q'	c�R�T �%�>�'D�Z��}�`"$��!�Cڻѫ�P�����woP��|k��"X>�0�O��t|E���K�.��m���.KDC������ƃ�u�����]�"��$�|�A�b#��-�޹�,�]�rA��j��.�{QD�Ժ��|�,����M�����n�D�����b�ٯ���;�'�'QEǄ�7gq��RԨ�����z���x��4��Q̉_��ǼԂ� ^s���ӡ��.���N������o@3�H���V�J��W��!6��C��7���⻸�Q�Vo��������T��P��+��@ �U4��a�������(Z|+{D�`�V_{UC��&Q<]�ٛJ����n��a��-�s`{^g�i�h�v���,r��*���_R�1�/��r��*��)D]��i�/g���L?�"�rm�ϙ�dL����]�-U�3�HGc���%��ߐ�D�E�BnZ�z@A�������f0F�#wMBQ�!����[!�J钵�]��'���el���نҚ�W���$5A�Y�����z���.])<��&q�WΒ�c1mZ��
��%��upR��4ܭ��w�� ��)�g������c�W�R�0��tʟ��S���ȟ0L�G?�@Q���:{צ�1gő�rUU
�U�������*��ډd$߿V�,��1z�q�ӄ�J�J����A����P̈%�5P��ۥ~ߐP�~����fg�.���]Wϗ�
�|_9� L��Ϣy\{�����񿽼�s��v7s�tJ��i�}�?->�k4S�a����2Y��k$�|1/R��f����]S�,�hw�F<�_R��t�����03}��f-�P�F��1�ۘ�%�!Vm�t�v?�X$��r��t��0j��JjD^�gy�	���}	sxAT���k��?$����B�a�!��ٓ�FAؒ�am�U�z�"��?�QH�m]؟����9p�f�
�#JƱ��E�,��s������=W
Ɂ�O�N)sآLu�k��j�q��Z^O��W�k�dd97�	��S�/���[a�"�� iݢ0hDs����������<�pN�t9�gqo}>��)���r��D������lB���cޑm,��^���Rro�1�3��/�(�d�.��Z�2�}� h$��Yn)��G�:��C�%��^�J��/�'W���p_X��ww�uF��ltJH�fg\��z��g�ì�n�P�~�mҏ��8iKIAZ\Ut-V����Ok	������,MK��ӈ[��52L���8�Q@T���i >u5��/O�o�z�L���d_8�zځ�I�����@Q�H'v�P=�
V����g�~� ���G}
�o�h�>�/N�ׇ�Sg�>жbru���ف�,�ః,ax�x^FA�_G�A˪(Z�ȳ�h���A|7D�� ���  9�Of����d�U��Ȣ�8������w�o_��	��V�#�7n<](u;�/g����#g�(�l"�f�;���^�s�F���"oC���%mdy)Ф�:����_��BBB�@���DW�`�L�D�V���:���0�ams���@�K��q �8I�7��ΔU�]�:.s�2�h*�>&�M��<,�
�{c��'�:h@��碉1��K����8�W�G��l�iU��Ŷ7$�3��;F��H�?�������u�E,N���0b'1��$��Ƞ��I����W����u�h�Ҭ��9,��ԩJe�t�\�>q���}��"2)Jꡲh��Z]T���"��k��C)6�"�&���=���K�v��*���!�v����H��x�Kz\�/:�IB\uۑ'�D�Uv���޵�{��Z��v�NG�E	L5�K�q�Y�A�߆$�L��a��^!V+�:W�T2T-j��1Ox:w�������d���ٵ!�i���4�PbB�	��>�$���N>Y�U��*�
�]?�c-큤�����uJ[�,�-/��y�YvxIP���Yպ-�m��P�7F�v�EH/�
�֒	�ZSǇ%a�QbW1v^�Ļ�L�Є	��˕�c��=�O��	�N1�"�!u�J��Dc\�=�����'Lp�/�dY#�I�&m;ו���)O����o����-kh+p�f�Qof�	;Vq�}��ԉ��b����g\<�X�	����75&�ؗ�/�:vC�X�b]��<�Cı2���O�ދ��)��ݤx�_ۇs������C�yd���Od���i��~�G���\Lna�ˍ�g��T.V���QҩC�}�� oٮ_��D�ˀ��  ��=Q,��ѦRO���(�L�¼�2��j��¨_����n#DE9V}�T��8�z��C�:е.H�nS�:��o����%�I����dV�V��<����$�4�w�����
!��+�jE�:6�5� ެ�ޕ2�1��//���NE��`)4�	
��kt�O?��5Bh�~!��Wh�8�Np�w"n�r�>�񝎻���A!�����/���2��ZL�����|�)��ᰠ�0W\;vI�"ߦ�q���X�j�'re&�������Q4<8���n[D�QK=t\�3��&c�'1��˺]J	���?r����>nm��V�E2��Þ5\�~��R���%9ef����MB�h��#\%��1��dlKi�A��e��(��6֝�)]���*.���m��!��Z<��q������lZ,P���L���ߥ҂a�,\2<�B���6F��dg9�nK�6��"]8s�x?U��~VT���X�X���*�$��Wr��C�1����NT�<����rhZoo��3�}f��}��f�t}M� �������`�E����g�d*c�k�,��c;Of�Y��Rb��M>j�YF{�|Ñ�^yd��3��/I�ۀ�~�(�9kb�kO,��1�� ,0�#��^#ԍsO�Ev�K�,EH� 3r����|cw��!�4�q]�-3��r�C�]
ߝ �ԒH�#ъ�t(<�-5��ы��
9N�~I5)��2A��'=�c��/��Q+1�"��D�4��	�m�+���������"��!\��7��v�`�E�'(V��r��h��p�S8��:=0'H����������pRA��X�H��I�2��"�F��γQ�ʸѓGݶ@q�>04c
��w���%L�^=������SF��f\�R[d~��[]�6ǒ�;��&���Cd��gؔw�<`��U����1�W�����-�Y���?ۣ�k��\~^Z���9�Q׊�v8$3�7�_�4��b���'b��G�?@��(w{�~m���D�G��%��G��B�.ь�C�{�Ú��cnR�u�J{��.�gU��3���,�����
\/o��`�5�<�4]2���w��k�3���P(�^��nO�G��u��@�ǅ�˪?�q�E���w(�1��Y��\y�9lu�����<8��<;�~�sT��Օ�$(Zn�J�'f�GO��$2lF-�n����U������>q+mE_6SV�B���2DD;{K�^���я��X����U��1��x�0:5��U?F<Ƭ��q6�������Yu,��u���bm�ӯ���!���y��L�X�ݐ�$����r�a,ɯ��ge�L?��mrY/�������R��+˰�M��غ�@��ٓ��^�1�����"x��p4�C� s0�w��Pj��U̐�6`Dw
 �7y2@>��-��,�wm˗3X��?��ȵ9�p���R7�9��=A�e���:Y�e1O8�=:��}�2|+~�Õe���0g�ΪoDgE[CI�o�4����.��ǭ�q�t�sP6��x\Ӟ) b$�}���C �,IWD�O�6�9;�%��iyhQc@������(��`.&��	sf����� ,y�g���oZ�C��,�I�@v��� �_�|��h8Ї$ǿ��q� �g�Z����s�;a6�Cށev	�D���׃P,l�w��7ě
��j�V��m� 1����q�by��K��Ħ���ka�Z�+����P}ٴ�[����⓬���U�;e �nnu˙^����w
^�����}�>̍�����{���<��cw������fC'��n9�F�k��-O�P�� 4qtV��AgU���V��G�.X�;�\.��`��!���(����[*Cu�V�X����C7vS���]������#<ƀ׵]�Z�]�8��x}!j�ީW�P�0�[�詬@4�q����sL�'N�EU���[��&�Y߸�h��%����i<�ʃR���X��E߾�{��.<M�4U
�l&�Ģ����XW�(���1<���/��ڢxSS�p��S�*g׀���,BH�4 
����bO6�A�-�g-a�Mb������>�6#�ff͐𚍑d%�B-
���c���l-C�6z��Y
�*�@HHU����gu ��p&��b�zϾ*H����tۻ"I)��)�-���v���@O��Q#�E��Scc뮦�u�qyх�R�$O����Ρk I�^ P��t.;z�)b�CK��*O�ߎ�Q=���Y񑻀����-ʘ�:�I1+4�v$��60�K�B�7�g�U���P�\s�^{��><�tM���Խ/��>���N�a�tq<T��fZ�7Ug�Z��Rx���?�N����3O�m3��p%�kj��9Q.޳���g�ܽ�ܚ���{�Gx��y�1��T��9^��4-؉�ZP4�^������`}k�fu:K~Y�'��ߨY�����pY��-�VC�� ��!��]���;w�%�o�Vl ���%Q���c<����PK�(f�� `���
��o�����������R�ML�;�*䯈�}�wY��3[/ �n�Y�E�j~��| �Xn��f}�� b�HVP�}�WY�p��" �ф��@~���9o]��G6-Iൕ%��9&��s�����l�Ziį�
4ӭ#���sڋ���\���B�&��������cᖰ�kW��z#n]N��k�:���}��е��ݣ�Ю��ǆ(w�Vp�^5}�q�9e<|��/���8e��]qZ�8�-��	�I5�G6g�Y/�6�D��0�Wt���xڦ�"�l�coS
���l޻g5[���'t������-�~�n�C@���CV�n���"2U"���,%��m�ցEt�'�u�@s�4�����)���ew�TO�D�)��&�9�CY~ق>Ï�l�sխ��#\ɼ�g �;�%"��ߺ�թ]�~L��}T%�Zf��!��E��{�?۞�Hε�3��@�l�|�41�
���Eצ>�9��>�f�
���������X@^����x��M�rBD�G0�ʻsK�WEt�����м�bN�[����q|	.�,YE���N��Ϭ�`G�"q�~Eh��@��'U�e�مztܘ�;g�Nd�;����r�2h�X�7�U[�oG㭝Պ�^�Q��uQ��q�8gS7ʧ=����xMR
d��j�I}��.5�"��k��'A#�3RiZoq�}鋴ppķ��7v�@ xG[�H�+G�{���'�kČW����5�>�'�����K�����֍�:^0�)yu�5�Lf�V��2|��N�sK�mv���5���y�7���w��ak��d�b��my�&{�|P?\��bѦ�ڤ�	 ���s��f��w�W��$�Hf^����4��k���|Z6�ޏq����U�3;�~�[<2:�k(�J(��0�6Q!�e!IN8ףvx�ErlRg�9����)��N�r����M2���w?����[l���.1�#�K
>xP�~官�΂�>)���<����O���Y�&��=\1f4����_�&�Ȏ�����,�Rʥ����\BGm�5�	���xPm�NQ� ���NBdD�4�����'��Z�_
0�p�-���"�dT�Ec}�b-%o������X�M�+e]�Cv���������g��/ݱB�T�VN�w^juk?LI�
S�Q�[i��>ׁVa�+����=#PG� �����e��+��|�-����ʜ��J���s��A��V"��s'��8_�.X��{8�����RO_O�"�����r��3��l}<\f��2ҲMq�
;�Z�W8����"ȶn�&-Вߘ�S�x#"��H5m�]�f}���@Sm%�lx�0Pm�
��`��Xb�����x����߹U_��=�,�B��T6�� h�s��ş��}�J�	XP*;ɫ��,��n���M��=C�6���N����v-|�X�z��.-�<iER}m~X/�`eܥ� �9���]Ԩ��;�Y}:to57�T5������R�MY*�e_�$��L8�i�~���)�l��Z�6,��s(��c5�#z��C���ˬ`��m���2)��m���ϔ��Q�nr��u7�p��븞2E)V��S�H�C
35N��j�y���M���!����b�.����j�+��;��&U;��2j@�wJ�NY-IZ��r3��0s�}���I���)&���N�uK��Th�ƥ�=�)@cb8*��o�Aю�P[3��L>���n��?�k����HC|��Lh�&,X,�rt����n"<!�jGe0>���s��Z9�Ds: �R��v�W,wʦ���cc���dU���PR���z�\�R1��O���?<��Ft}rx�*�T��w�6��ö�W��>^���䥒�MYt5� ��n��}��:�-���(@k(��H�C�)|<��v��˻M�����+�!��T�b!�k��ң����.� \*c�J���k�+�J�����v��Ύ i�(pP�r���ѱz����A+���/�DmZp��]��v�K(�&T,��P
Ud�<[}yV�Aɑp�)�"-�B��;k��q�Vn
2���P�N��rX�A��n���F�v?�P�-��B/>P���7�c|̓@���#��$�����{�*a)y�^�l4�� ��$���;0)��.v��_~UDC7x�d]t50�h�E��){�e�<{[%S�fd_G�I������P&3Ԍ�VAݹ�!�W�W�*f���ŋ�П����tL�Q�<�[M���,��F*�Q3����<mh��ݍ N�p�n�b��N�]�-�*��=���o���[θ�,�4���gZ5L�v�Kao�jeF�E!)��**�,���l�a�"�:�7��I��/�Յ�T�3_a��b�I�1g�gQ��q�����@����I�(��n$���82g7�0R���\}
�i���ͮ���T�.j0�q+��
�.׬u�HՃMC�{Ej�.�w�3����P?�����q[����>�Q㸚[��P�Ԓ��Yhؤ��z��D���U�2��Y�I���!f�ʇ>0���b̢T�k]�Hȉ��*!9����wDQ�R\�wHs�*�#���V������b�(�B����d��i��5�J����Ӵ��;�d��}f������[�txGeM��c�+Tҍ�tz�!v9ǹ�B��}�NdFz3HKP��3��"������(�`XAV���E�ɺ�U����0��1�af�K%c
} �Z��d�����	�Ug��͵��P����*[G'g�D�/ކP�e}[�g��@f,
`lGC�d7��F`��*]���PE%����#��(X�r�92`�P� 	�
�U���GżwIO�H!��Ɂ���+��M���\���ޑ�A�0B���J�k3�B�Y���l�AqtH �[TK��
ha�w6��寙�Pv!�栽��aԉ�����&q�f�"��;q�9̮�K��N�쀊XS��U�x���eyU��Ic��ǸZ��2w��I's����(E(Z���U�w~��"���}�k@�;�R���5���FA7���<��ZF�.���.����FyU�΍1��ze;"jv��om��ya�i:X�Ff�OmN& ����/?�]� ��^6;J�d�Yh
i]������&q9D�O�@��C��M�!V5锢��`������ey
���G�K�ޕY���?�4b��kEaaZ3�û�}��c��6���IN�62����%B��_ټ�LM�-EL7���Z�UX����_���g��\������+�T�e88�?Y��`�ި2����f��G�E�؍8�:�!8y/j1�|��JtZ.�#�D�:؂ O�(K�@6*v�䕋��sx� �N�X�5��n���&
�N�\q�(�0�.nq߯ ����&�P�"N��@�P�����/��S�m*p��%��<�D�*�&�0����o����o�z����k�r�/���z���_��.�H�MĘ���Z5.���c����ޫfS}�9�%o��>>X��M�elk�oAw�@N�!L�H�|D0�s՟���|���M�#�|.Y�茷�3��n ��9�d������t:˝>u��Q�
��EL8�(�B�@t|
�{VYE(�䄓h6���y��5��Z�kv���tim���W���}��UĽ~V�^!�$��c��e����g>�3��{_�]�_\��;{�?�2�Zc��o����Ete釤��N�ޖܸb�ʜ��(���5�8ͫ����Xj����4�[1�&R���v�SJZwF=��Cs�{5���͘%ш\��w�M��ޫ ���ͨbpolI/7n�iQCJY��F�az&�&g�����y ���9�5��nǻ�[K�^ȑ޷��,�u�Ղ�ޣ�y}�7�Q���2P�X���h���Y�^�ph']=�!U*��
��M{�&m~���Tg�A������dFvU]e�<	�ć���rQ��>�p��8F80�Di�����(����گG�wnV�r��d��Û.���b����C)�:�z��r vq)���Ԋ����nfغ��NS���1y��.�N����c4�>���z��`N$~�����մ>��2iq�c!w/jմ��Gy+F�t�.�r������he��H��̪6b�e�}��W�z
�՗����a>����>H���*]ڣ�ǲE�*��;8���,�/�)�B��ڊ��*3_n��6a3� nys�G�+q�
�o F˒7�?��JG'y��Ҍ�	���R`�G>�Q��H�8��i2Syd2'���k�~ܯ�7���-Ћ��1�y"�8�[�-!r���y�νmu�ʒ+��Jq�'��]KZ�i$M*b'�?�J�D��<n)&�i�[8�]FiQ��s�\Z��:�W�P�a��¤��w#��6)4?��=E�Y�gn]ă6t��h�fAh�G��/�����v�?�����_��7d�R�r]?�\ۭ�3�y#E�93h_,˜L���8FE=pcuO\njl�/���8<N-/B�/-%p���#�������0a�:��̓u��Gn.����oN~P��,�&x��1�%z�����b��p�/��i�/
&,g��	w5�H �o��=���P�k�����N��#TS�>�� �S:�r�����]���52�{�~����&OH�^���2��@�}�� mUѓ��Bj�\E��)b+	=Rn'�[ ]IHK�ʜ�*��a��]-�%��bvk{��ɭ\Ť�7��?��L��AWrl�{��TY���e����J�<u������Л�u�`æ�o�fd�u���ܨz�;�@�^Z��B�x�*��6�:10.}
��xA'��?������ƀX���{�����+��_�>�V�΅͹V�%����h¿(����5r+C�0E�jj��RVZ���u0���F��jXi�U�H�%e�f�9�ȏ��H��ټ�Y��g]�R�i��g�N`�����֬�Br�>��l�@~T=�;���<'l�M�[�i�ͷ��26b.l�VH��e׺ߜ0v�ׄ{YF�Qy Ȁw��	�(�2�`�=t���2�\�7�ٯ?]S��f�X�B��gsӐ���ۂ��̡�~�Ë8A� ��X��xB�<6�3l
����g0��#�6�[+<���G!<r\��]0Ѭ(�
Qi��ૼ��S�`۪��_rB'?��޻�R������=h����Z~2�?�/���Ic�jj��	�W��JYH�'<�����L�T�l�)P��_����Ԯ�2���E@  bC̜S��V�Le8�ܶ����C7�cy=��K],�#�;�`�0�#5�3� N����V|�*rb:��W���(�
R������r ���ӤV��X���Ʀlg�K��3��[�J${o�KH��\Z�\���QSV[ᯗ\)�1%�N��I|�����"���>���\b�!�ߋR[��l'ȟ���6L�8u�N/G	n9�`�xqP���|����w��n�NL �K�����	���O�gt*T��w.|f�7��^0���,	�}�^�u����� `Fpoe"���p�J����-�㫋I����~�#b���Q�^t5��Z�r�u�B��,E5��j�y�3����/%�fVq)����E^��&��q��8�8/a̢r���ȱ&Y����+
�)�!X}Y�C��\��&���L�� d;,�G�����\6���{����nX��&�V�p9O eCAZ6��;˙��l�]k�.�%�H/�����lb��ͽ�\սu�����	�.s+=�ջ��7'z�"ꕙ�4�$ �x�;�;��1�;u�l��=�x���{��D��dB ��boEC5Z������)?�1k�_醍�m�`6�A�A��I�t�XG!��M)x�M�"ҹ����x(j����>�b��GvhҚ��u�V�r�y�N��MJ33VvW�C��ZE��*:�8��B���7�$yCxQ��g�o|�L�ZK���_y�����g�����c/���tHA;��cM��V����(��+Mq�,j�X�~.2ɪpr�{���Tj�E��HH[�l z��O�Ȅ]�W����o�~�R~�Y�s9j�R���X1ik�^�ӣ�([Oml�:B�~���Q�Nl�Ji��cz�C@���Շ��^n��1_|�1�ʇ��~��~Th_��ce"��f;�v[%c��o!��l
��.���܁�eu)`������6&�̃�+/�DD�D@-��;�g�A��2	�'Ay�/l�|	5��t�F[��<Ҟ�2.����`�,|�.�$�1>�s`�yq��raFuk��.�&��ZC|��'�T �:Pו2]�{w����%��nvW�nt�(-�^E)�Iؘ���$�}	:I�֎���5 �[��L��1�,Q��U�7�d+$�FL05��_��QA�Ovpfۀ@��K��{��1o]Q���<wg-ܒ�uub4�Ǳ;�&œ���k��W(�=�+��;��C���#&�/ﰘPJ�1-;�:�������o��)� �Wg�#g�����@��`�w�vN��?)ъ�~�~SwmȨ0���Z�GnG�QK�b7#�&t#��*|Ň��O�u*1����X���mAp��V0x�:R�#_�v�9�E�|#=4�*5�(��/~�}D�^F�d��U�����f�C�9�nWW��{.MٽN����$�U{*ر׉�oE޼xX�? ����)R$�R��״����D��a;��%�b�'�d�_�8�������gVŤ��x�����L���!h�Ӊ�����5h�����$�f4���f ��Yj}��4uJ�+d|&d���r/�.&��)Փ,؇��΂�P�[ԭK
�ũ��)���A4`�Qʒ��tt2�މ?�܂�<�pP��vޟ	2�r�x�Ȏp2�s�p��m��f=�6��/W�f/��������s��:g��^iH@�h,��N/^kHM����J��s��5fN�]��IXe�NI�"$C�� ��?m�\�ֽ�_�L��gS�1r*TߠK��8�"����ۈRQ"��ǨFD8&�:!~�,F�#՘��� �v��d*B/Շ<+D5���U�g�I�A�=����+��>л��i�f����澶^l����� },�(��W�G�#M��+{��ۘ�.H�T��" ������� �Eǭ���<�bN_Q��C
4�gyV;��'�ޜ�f	Z�T�y(����p�o�i"�o��� ��>��x�#��27Z%��BS�bD01��".�`�\un|׉�馩E�ɾ7���o� %}��c)-B�<�BH�Ž����g�Ok�}t_�	
�'��g0f���D�(v�z�Nz1�������}%�!L�s~�$1@Z�b~+���g���--�͈��b�d��{���Ep�&�5�{uv���k��=N��U��v�i�}	a��ښ� �$��D�VF��z3�������¼v��3���#�;F�G���P�ᇡ��^I��N�?�n�>+O�&;�>'��V���a ^�*��˛����u�Y�����օ����I�q&u���HI�Ix�����i�ѳ��I�l$f�n�V4=m	P�|��������H��g���0;Y��?R��	����#�f������2�5��г�+L����;	���B�*M���1#p3$��R}�|�Qy�hM�1�ƴ�#7�X��3#w�u���}*����'4N���V;9j���y�c�;+�9�2��/�B�W3'�}�=^�Aʡ��CZ�H;UP�s�Hp)�ʮ�&i�s8�bJ>���/
D�D�N �N�9J�X4�{�]oh�y��[Ï�&�΢ϯ�F��{O�*.�j"�I��BȌ���Yx�M�Mә�TG�\=H�m�(n�6RǤ����y�F���M[�Cy�A��O)��9�v��Ce��f�mϢ+J&� \�=}�=�J�$��'AuU@<�4c8��d��^2X�#�־���q��^���͙e��p�8����%N�����Qu���U��&�ե����I��}_����m`�\��s���}	��>��\L�����IFj���{+�(u!��	|��O	��*Zʭ��D^�X5/B.�r�V�m�X
<� �\��:P��×��t���sϾ{��;rFVb.�\�8J1�T.�!L�ȅ����G�d�Q(n�X"���1���)$�ac@���q��,� P���9��K"��f2��{��#S�_9M��x�2E���Jjp "�?$�s��>���mCiH}d�f���8~檆��t3��O[�7w���@��P_���vm�o�D�s$l= <�!�eQ��[�-٬�D�����O*5�.�g�[Iy�
���F6@hݹ�$��سW�y��	-P��xy��K��F�.O+~D3|�0�'zֹ�y�f�}�x��baP�$�!��[���]��瘝H2����@��i�dCN�������uۍ�/*gb}�'����	�-���q��:��K�bҁ�����Vv�O*3��jX)�\����Δ��y+�V���q�b<m��_?�����5@4Vl����9A���mȧ}�-f��w߃J�a���M1�K�G�bŤ	3��G��b�ζP�P?�3�0��^4�qp����	��+j��{��+(�D���[H�=mrw�U���V@3$�[`��cl�������8��˻2�历{V_xx����b��@��`w�=qK��9>~b��������H��2E�Ū;�EQ���Co�-� }�ZN�a����1\���=b�֐����R�Px:�P��+D��o���<��I�G&Ņ����yf������;���:�(�<�6u%�ʵ��.�K�U����<�v�S������T"�������l�Ԑ�Yݑ	� ���f��+��̎cS�Ya=�&�9Q<��	���%O+5#�����+��W
�����=*d���a}]�����"تO��W��P&&�(��	 [��e
;��������P<0�_<����q��� f�&����8d��l�	�@�Pt䡰�Y`�Ό@��,й�_7C��nt�C��އڹ�Y���$��ǘX<-��C��R�jS��Y9���)��З@�v�t�I�R��W8�x��5�	��S
�qi"�ƔfPƝ�.�)U+�GثMP&(NG�zڒ��e�!�J��N+��߂z��6�V|%�y6�:��VS��*_��G��`�.Pܪ�&���;HL�4��(Rhu����0��eN�٠�� �'Sq�1�W�w�0�PI&׫|W��H^
�%��d�F�_ϗ����.���zRl�Ɏ�Vyu�(S�'�)�i�c�!2%��Bq��@����B9�ƒFT��s���T
�ӵ�F�7�(�b�����ˆs��Lʎ���=oy�y��s)�!��Խ��j�B �2��s����m�F��?����3���R�����\# �j��7�C�+IŜ�i��^^Qc�6�!be¾E����yLˎ����䍄�!��5�0/����<D�y�ӆ���NX0]?��^�b�w��J�P���v�ۙ<�^�|�EO$�wL�ȋ��U��)�vjQ��ܜC�3��߀ލ��Zk!ߓ� ���8�54?|?��|
<���b"�-Q�*�F77A���~ �L�F�c�Q�Z�o&�QG{SGR�t�fj��NK��	Հ�H�6U�������Ǜ'
��_�N����J��Z|�Q�T�d]�D�0�	�/Y��]�+�+U,�����B[/�d��{�z�����:�����<
�<J�gn��,�A�>�o�Ί�Sˇ�*פW�Y<�|4�$4+:�L��QC�҇3��5��w%��������>��7���Ϙ�g8�Zv-�B~�O�}
F��D��]�>@� �-{T��ix�[��۩�oB��^^���g�Ӥ�u�6�֢wRHB����(e�Bɔj}\JGo4aq�Lh4����|�'?�㯬�M-�F!D5�����V3�u�À�ۏ����~��_ZKґh<x��
������g���#�9���W��B��n A�o9;b��Y|Adx��Țd�&�Z
L E
c1�ɣ��XN�r����.��He�s�Rx��'舔oM��QC��У~��L��VZ�Q�Vc�> �-6�4���I�_=�4�6�w'0�D��^l�R��j;�a���z��;�NmdD���Pw��n�ĝ赸���QUܝ��Њ�0^��w���ڶ��Ge?y�#��{��~ǵ;�7�cĳ���EN�w�l3���ɔ��}A��K�C�}o��KJ�ݽ�"��Z_���Q�S�q����ƘPutzCiD�b�x�gG�wՁ���'q|B*����BC�`Mys`���v��G?��z����ad��>?�ثz� T�l�2҅Ì�;�T@&7�e�	}?����!����*h�j��~hЮt�Cm��B��Ŏ���+dE�3����
8z+#K�Nc���zFq�O�d�4�6x�6�xM_D���}qrȶ\՚���LC�f$��^З�\�k@T�̀}(��v���,�Jcx�v��KH�{���1䔍��'�2.�+f���Ҁb5Ƶ?T�[������Ѫ��dW1����HyO5�
$��b����:XH�w�?μ��UO [�p&�oӧ���d�`�JNֵ�z�pD�9U�AL�{P�i�	J�H����\S qj^��W�.��K,����}�B�ñ)�~[��:׃E?o�t�N;�ԩH�U�Bx�0��~Mm��l2GTC[�BHU�K�=e#���A0�a�Ԟ�?p��a�����T��ۡ/�'�����saSG2YW����G53Wj��5�$_���q��C�x���G���{�y�Q��:�G����Kߗcԉq����«�W�-熣��i57��5�#�9+J�b�n���-���b:���ZaU��Zp$�����Op������9Ͳrq%l��A���*lF@p�+����5w&Ș�)���4(ڟ�/��r�d�Ϻ��]�@b|��a��+���vZN=Q��u�Qy̥�O���\Јֹ����`w�_�����}�X>��x,5�8ד��cB������87��ƴ��igw�����B�[���8_��i�Z�u�H�m� jM�B��(6���������)������0`r���􈸈&kɿ^�y���ky��TC⟯G>�� ���?B0����3`w)�n3�1з/.�|�d��U����R2��>�P0���׫<ϟ`7'�T��(P�B3�����*3c>f9�5 ��\������Ң�
Ӫ�Au"+�0�·y5�X��Dŏb��ɟ�؂^m0t����		$�G�U��	I�^�2)���ׅB�Ǔ�=��JW�щ�vN���$��S��0$_8P\�y�)!,DB ����Ao�6D����^�F�}rN ����0J��%�P�p��~�*����c��-���v8M�ᕢm�aop���z���n{_��R�f.~��H͠ز��.]j��'�����h��5O��JT���q��4�L��YYL���`�)�hF+o����1�w��v2.�g
O�R�ld����TȵdOU=kq����m��h��5�"��Xp��H�w�hh�D��\�@�OMG�+����I����Sޡ�l�t�p럅�M�0���.��w�y���m_v�����Ą����U�,����ӆ�~[]�e#R�)a���8��F><Ԉ<o^����L�G�1��3(?�~]�iy�]�\�gP��'G��\F?q#��N�"�ѫ���,��o�kg��=����?]c�~�����z&(����i�sG��#VH�gsڿ��6w�	j�<�	j�yr"�ܖ�����$�d��,2�սlYArݦ�w�Ch���Ŋ::G�Ĥ���IB�X�;M��2Q�qD�R���� B�q^X���?�-=�*��@����*�o�n1\+��%��>��}`��Ӈ�j�jd���}b%/�����Z_��Tm-9�&qd�f�;ʠ# _���O�BE;L��JC\\h��6_R
u��%�fB�j<��cѤ~B_�#��x�%9!Q���Z�)/�����M�n����hQ^�r_R%aR|���u�B����k�����P�؅Z+��T.���G����,��˫h�����a�j���ϐ�z4S\=�^���9���+d*(�K�.LI��3��Z]�� ���o��-���5��f��ɠ�j�T&ff�ؽ/�b��:}M��`%J���N 8_����a$�[)������;L�F�.��a�<�|@�1s����_TKN�À?���P�r'�� �����x}�}P� 8�%M,�z\;X��MUc�Y�f�_6,����\5~�� �p�V<�$�Fx���wކӍ��w�O��n��Ґr�Z��)���m�U��ጕ~и.�����P� tٚ��BL).Gĭ�̓�4c��/6��"��}�ЖZ�� �ߵB�E�jܔ?K�?�5�E�4C����˯�i��]�,�e~�o�ͫA!�k"�rh�g�A�>y/�O���8���<	R�iՑ�6��^�x`�$'*����<t>��D���m��Q�<-�g�V�T���+)2�,� �:�p77Fq�T垮U�X�V�-�d{�����"�$Cx��/�Sg�L�1T�~έ©%�:=��FJ�͸�V�	����Y,��(狀�Z�E�
B�ҋ��_�ֵ#�ݭ�r�T��U��j`iQ�N���t"}��ܙ�oź����G���L���֟���=	�k���_o*Sz%o��y��b���7�^��ua�����a�nyV̦�7�j� 1����kf�P�Q,2?a�҃�L��^Tǭ��@�����Ъ໩֚T%�'ә��A>9���"��4�c%�lV,����,a1:�"�G*3�nm]ื�NP�����A�\�g��eL�=aڻ��u�}�
���B9���R�'�9GRr��6S��*��[�2��~K�&��zs{�P2%T��1�]=�G�n-&�4��g�C�D�	(S�T�aN�D/���o�~�=��$�8�}��⺎�!��e�9����'�ڥf�nv|�k�Z4�e�hD�oA�or鬎0�3��hI�K!��!U�H����q
d���h�#���J��VJG)����:~���a
jY+�[��c��`<�����o�g3�uG�T��[�)����(mZ[u�t�<���,�'T�Z��Pۗ��a���$z�HZ	�;�u�B��ϕJ�'Xg{L�R*��-�S�\���Y�maW�`%�}<�0�~��L5�$��G(��o��1����Z�>� a2r���_�=�6!�6��s+�4ƆN�p1�V�����<��g��4�\##���d��F{�:|pke|��SzayZy����I�x��7}H������z?^W�ڤb_Α��w��j�t��e,N�i:RLDB%(�����v�Us��������N�c*>��y�1������}]���=.��|C��%�e����S�r�"P�u���L�Q���ͷh���pG�[od�r-N��K= %�dȖ�y��3�A�(�2���2��,�(H{<��PoN��}(�^BC�-�W�Rn����Y��|��{���=.�>D}��Y�Vbŏ�y<Y\��@�Rfj�i�a~�VR��P����b���Gdif�ji}x/u����nR�.��7`5�1���|�r�Rm(i��?�]�V����տe<�t�k����L����-�B	v�0��|Ί
T4����"es�8})EW_�(I�iU��Q��4�_���n�%S'?�jd��o�O�H���tQ���V1Ր����:��^o.Ǣ
~��i�>_}Z�:"�9)�ͬ2+伧�8��[/|���ZJ�&�oZ��c�t9p�y��ϋ:Hnpr��|^�ٌ�H�J����Ob��Wj�,��������t�[i.L*SA�@|��5�줫�3�b�B7�!�#۰e�>��� ���|Op;�X�(Zo���r��֚��D��u��X�P�2�W���D�!8��чfosk�4֧�=�g�'м�	~�:�/AU������$�;d�� ׆ ����9�|�L�3�pk6e��{_3g�&�sH����洸!�h`a��`jX�.�)����8�+�?�,�`W�T�I�!��M����S7}e��RŲB#�O�O'��ˣUP�~Z7��4��%���h� �'�P\կ�骧��?r����M��x���#�P����ۋ� J��� g��,V��?[�!�)US���e��P�6�w�ϩH�2�TysJǣB�?m�������%`��J�i�5t�����$��w;���iO����P�+XS���(ɵ���;\�0���Ū��� Z^�AQ��A<b��܊�'1��Z��9m��#�y�;�����cg�<Cċ���C��ټ�D�/fQ6����2fz��~�H��W>eMj�!T�@�P��p%�u,�H���
i.W�7K�l��h�,L�}�}�Kܟ`��f����%B��NTgĳ�OJ+����{�Ժ���� >���mD�#b�m�o����T�7�?`�6�Jw�|s`�П�9��G}}�.����i����ܿ?�/�3�c<dw��*��6����#?TM�c�s���m�Y���\eP�ٍ5L' ����8�����>�� �C��(����ጭ���� S�I�Z0%~����G����F��Q���0��]�
�"�i
��k*�\~�$�8E��UX�oNojw�#�9%������i>�J�����r�\~��5W/���*��yYk�E����[����"}y��st�f-;|���>�WK�v`�:� ����E�i��ʭ�Z�U�z��l�� rҟs�Qɶ^�P�)��3�g. �c�U7X�K�)�U����۵��Dp���[���~��=ܢ�sby���80\J�`Ηc�p��X��e�����>I/�a�./5�S��s2��u]+�3� ��u��J���{��ȶ�&B!2P�@<3G�G�@q���}f[n: @��4y�/��)�#%�^��>��MC���飬x,\,N�1�׆s�퐳�8���n��
NRu❺�
L���fhh(B'S�0f�툻ky�[����o��Uu�!(IB9~$��͹�s����}l0׶ầ{�熣<�ˢ$�T�6M��2n�H�(�C�D�
 ��-�V�'��q{XZ�j�K������Z��"�� ��(�ã�{e��#1v��&|�*}�kD�rK����m��rnP�]���s��Ϭ:I����%stj�/i <3,Ned�#�0\��0�n���"�k��g<�JJ�!9Q���,�%8����e�nF���H��� ���́��ک��E��U�h��9ҍ��`�?B֒"�C��+F��M��E�-�J�B�����:  JIh��$4���潰�������2|#K�8E; c?g�������@����g$J�4a��,.�{��ֺ���=&%�Dz��'ĵkT^���9����T�@:T��P����< [�X]#Iί�$#S�^�ߨ)G��O��NA ��`���5��|�r���qC\����ݏ�_���z7�e�T���Q_`M-�_}�H&����*xX¯�&��V~�Vm�/4z�P��\r�&v|��-'9ӗ.j��3>�鉬��=`,i..y�6{�}�����u�$p+�b����%�I%	z!Ɍ[~d0HE5��	�;��y�w�vLq��3|��{1�e�����|�J�����#:���w��$.�?��R���ȟ�=���4�g<T��2f�ZϿ�j�i���j:1-X�j'�� ��K�Pv]�E>�@9SJ|��}Z��y>d���SݳJ���G�n2�+��:�x�6���fH4�櫖��Nt�m���j�=�bM�=sֵ��;mV��p���L��}�si�I���S�R�۰�`�kC������yZi��@:�V�J�Jz�;����"$2,�����|���W�W�-��?�p��|qǑx̟�z�ᰟP�u���S�˝�)$䫸�,/|�d~E\�db���ʰ�̳�L[��Z%��V���k��0Z��[�F��8��tOT��tn����4Nl�ޅ�{�KF��hԞ�"_��:��p��!�x�+NPd���Pv�2�K}��U���#ظ~��yI=���4�7U�r>���
$�� ��ʖ��N��5v%��z�������QM�"�L��t'e[����+' �4d�c�"t�'�����������|�զ<U�ns�����/n��$�W�&����l8�4(�w��9�I�e$"��^(��^����
;��o��	�+�KPqU^��ݒ�t�$G�n���I��/tt�}w��;�$6ɟ�%�R�W��G<�!������`z�4`�(�#��-;��b��>j�y%h/)YC+�w�Ӂ�������,�n�8ĵ�bڍ�e�I�y���Rf���8]0����߭����s�[���R�lXφ���/���ʇ��|��fC���?NAR	�U�K�⧞��:-�w���+��^Y.Z!t}=����s?=L|�X=���
}���Z��wQ@%���)���8"G���#���¦ɥ:����A��~"�J���.B���
�uӇP?g��CQ4&Nk�ܹi��8jȦ�|rS��?ܫF��z����v�EM�Nd�!��Se'>٭���K�jL+�s��`=� ��=$B�0-c��n9����f��z��F���)fP�"0������4�Xlo9��!�n�[9�?�%��FpJ̻+,�^��w���}��g&�bː�B7�--���'�2�����D4#����D.�}{�SK�8����h3�v��mM�F��lP2�"7���E�W��؊�F������_��q�ŹЖ��x�?�5�r�@p�rc驈�a�yQd�/��H�QR� 6�����[�O��mM�Q"Fj4>94ޕ	���&�t]��A�Љml�O�sL��]T-�y�?/s���WL����h�;FwLn��y�?p5�X��/h*HYGGQ?��D�e�F�^�^�0�cni����,Ę��W��>���C|�'�Df��_���q��uuVܬdn��+������|ER=Yy�u�؅��-�Uל�2K�9@��sj5�s�E�s�v2i�QF���P ���=.w��M�+�,��_<�C{�t��NŇ���uG�4�����d���������}�����ܺ����"��x?��u���`D��p���;�C��i�J��V$���5�$_oB�)�oI�ʙH�}|�\##�Wh��<U$�<T�.��q��N��yP��x9i�j�uϐ�6���Gq٣b��^��Ng���-��T��i�6�ЭߥԱ��T�0a�W$�2�^ڟ�E-�����Z�ɛ���\>���*�`8z<M�e"��f��Gx�D�or�ʲmP6��њ3�o�o�~���zD�a�|fhQCr�q!���쭖��:0�`ՉP
)���d-iDO����Nr��8�c�OvJ{�Ӕb�OR�h���hRYͯ�4��X����k�o[8\9�P\1r�<&b�,�իD��j�5�L?�!�9��`����p�ef���`d�O����n�Sh&Ďcp��
M��,�adƹ���.�N��^��s��[��z='�ΠSzێ�.j漜�̑�a�v]�z���ȣ�Xɋ��Ɩ2��/� �Td�����Cj�/�Z�v�[Ad�o)�u�DK��X�hƁ�j�ҸP��R�?v*B������#�<֚/.��8�0�AW�A��	�u!rќV~
)��0���C�H����/�,�̀0YK��C�����#8����s��������{���"�&V�����BS�j\��Rh0�ؿ>g��]�F�����,&�:Q�!�.f�^-lzz���eo%8��"���a%VjP {����x껩�GO&��� 1�G�;۠��t%�l�b�dD�YSN~3à�91���fl��a{�RS���|{>���,e(���PN���h��D 6��8aw@2�]�Z���~Cg��B���E��Aw�J�G�[��|=����-�8��b��ͣ��&��1h�����O�/t�����m��>�	˼����M� �'�+���8��� �F��h��)��G����U�E�<:Vis_�����xL��F=����
~d�������Hr��+My���H�E��˪�Ϊ��տ�@̱���ØW�{s�,1� ��/��4UX~�����@P�|P��Q��T���W<%3宀�)�o9�:���þ���%�mE���^�p׀�f�K?��do��
,6�7�W�$l��W,.�&�`�m�LF�@�}��1�e�.dR�x~��~x@�^�6���JiG�,�����*W�gj�F�e����a��O<� ���/��a���lk�t���p�~5L��а������G|��R�F�5.�$��d���.@�˱*&?o��ZF2��'��я4�pb�8h�Z���N�=��3p��x5!x�ꖤz�Ҍc���iNQ�P o�K�����E����'�2X#����pCr�0�,�M�!��2�D_�mV�6�+�<��\��`��Y�a�8fE�[�VG� ���L���b*u�1�)�@�I��LW��,&h2@���K������I	��x��2A�4VZ{��T3�xD���
`�"n� 5�=k_/��7��49-�ᅔG��On�/aa�"�%إwcb}�����rn���a�v�t��1��V��EY/�3�3$��w>��CF�f�8�%M><_w����!�"�v�|ux��J�����<BΏd4煚�9a� 4\�j?���$_�zQ��9<�3���tXO��	�ϞO[pFBZ���X)Uc�ڃ���h�Z��I�S�������R|���τ��N6qJ=�a���i-��p)l�gȵ���Ν7.�wP]"
��H|�_e%CL/O�*�i�)VG�"�A7w�ɓ���P���J.�R; �{��|��1q��ã>v�f�P�
�׍��AAL{Û�,�I�
���r28]K�<X�a| S�� �C�������V4��v�h�[������ërUƏp$s�a�*�_sC��mB3iW�
�3p�tGm_1j�+ȓL41lG�Ni���æ���|7"j���az��d���ض��TKhr1d�[�ڋ(`���,����{HRѳ�c�+a�1�-�Sc}*daȅ���9^��=rd��V;� rR*R0���'J!�B�5a��7�uA~axG>\��h"-ޭT�ŕg@oE�!�������E��V�R���atuuy��P����u����|RmS�o��u�2�?�T�J�ظw����鹂s	Tux��ѷ'^�ZUu�D��O�T	8h�7����Sy�;�@��Ow���W��e���:���(�Xm��f�:�`^�����@���3'Kxß�_�&z����V�d�m����G8#X2o�Zr�9|2u�/��������ԣ�ׇ���LȨ�+�yYD'����4�ii��O#l��!�}��I���%��Ź�0��b�6©�擉~:	.�M�.6[�F~G��x�qφ
�m�s$67��R|ѥ�ļs>I�hnF�@�)�=JU�Q5]�Jځ�?΋ȭ�Z�0@�g(�J	(�#%���g����1�����DU��<~����䞃�|k�y�6��/�S(M��Ѯ�u.�:��EpnE��!�U�rU�\�����YЉ����4�׋CJ�e-��:Ư\��%v�L}B�_�O�M]䃓|�v-n;%�4e�vȑ���v���Kd#�;��O9v�i���������C�j����5��5
mY��8c���{)����--��m��ԟ��z�>�{�}�#ud�2���~�s��)?5����$ä�r����i��,�,N>d	�UܜL]_uh���W������z+���cM a�!���,�LAQa3 �r�c�4�WT�}������h4J����:t.�/����꺣�@��d����E^��B�ׇ�ɕj	�%����l����*�9�2��Q@��a��{d��Y�>�������U!jI�ps���w�@`��{m_IS�!k��&R�'�ƽ�,n�,��0S�F	y�z��2���!G�"��(��}�����-��������=˚���K�?�r�ͥ��b�%��#3j�[��gҰρ 
�H�����.3\��S��@��#_��ejm��1�����p�������Hj�ӟUS�˕���f��A�u@Ӎ�\ 3�6� �ǹ!y�A�RO������kh�7:�±0<���i�]� �xbNyx\ C!�$Ub��CwqٺLOm�l����k8'�8��L�Z�l4�Qŕ�v	K��}=:�TT�'Mo--�y}�N��+���鬥6��V�����Z0��ȴ6�RT��Q߹�<�w#q��̿(��O��Q�8]���o0�|�V~WuX�M}z_���E�ة{,�N K6��NE1⛘f7������k���_Ժ��u��m���#71��H����a#}�Aw�;�TI�f�c]ǎ!�	E�թ��nî���^��T�Br�%��4y�W�+2,!�E8���f���9ᵌy�}�z����IJ�"��G���P%="O'#ÈTZ�Ƴ�Y�_���53^U ?���Q��Ͽ�����55tOfȓ���Cc���֡��D�eߞΆ����`D�u�yp
���<�"W��P��R4���wHSD�H��e�u�̛E�@}fd�`�2o���:�[H����!7	Y�x\Q�i���WȜ\=��a|��8*�}o�g��U��S�Ք~��M�� ��`�{��*�R����`/����3]��>�Ga �/Q�a�Y/��/X2�ǧ46::����FS�#@����.ws�0���i33�P� ����A�Y���H־����� �u|�PE�h}�~��Q�D����歈�����ޡqp@WU��SK��`�ȥ����]l/��=wT� 4��˓l����j��$zC�ʯda[~ř��d]��"��"]ᤀ�;L*�'(��Q-�/��bcnL�C�[~`���To7���@��\cf��W`㽇j="���u�L񸔳����:�7������Z�P����n���N��]����sU�u��.�^��]zRk��7=�'` ��M;���"�9nz�}�^��׉~vB�%��i���u�̢��P�>���E�JJ;x�(��47�����"�]6~)�����+r{�
 �c�h����+��JF�Yʽ���٭
�&�cR �v$���%O�n��[�@����F����`�5���ur2G�^�蚊�p�fj0G^>���H�}��Ԥ��1g��J����Jg͇�K9����B�x�-}�̉U�[-Y_e���%��7��L�=�mfbw+")[��WA�Aܱ�I��"���E)�<g���V�9��?_ �zU�۶͢-{sH��Í��]߷{�꼝�2�k�^��33L	�h(#���	��40?��u��H&�4��f��^����h�u�Ci��ٔ�ښ��:�員^}a�Q���"�8��`��~�}?��v���04��!֯�D����b��g{������Rtq������)�(���Z[��K�lt��K��@�X͟�&�j�-�ʻi�#�aȓ]���06�J͠ �Meo}|v��+Q�(�2�3A�V�	����X̒�c�ӱ�@�m���Re�ȋ���sN7�'s�~�,��k�B�4\��nɹ?�5:�V%#�&��{>�:��4���/ƥ��{H��ɴ�a»�
Յ��̚�~�����lo�,���
�@��e�7oeI���*��㲪-=Q��tA	�!�=�N����G!��	Λ�n�v/	E��8{1��ߴ�p���ES2�F�ɝ����O��C���Vw�+�;�?gPU�uXe�_E�`����#:Lq��BE��b$P�H_v4ۅ�%���������n�Fjt"�VZ�)l�X�
c=��]������f��׍����P�5�� �t��A"��`�������<:K��?�	�$z�L��|��z�k��Eƿ�� 5�#�Pv�W��A��Rϙ//��2�p�e�O�B�Q\�:)�L�C�*z-C+��l�h2�P�m8�==6, F,���o�b����:�*W񖂖DoD.nX��s���K�b3N8�z��x_hn|B=��^����!�tS��/�p�(*�F��?�.�d�G�V�G�h�M�;�OT�t�@i�C����� ��fS�b����"�j�+�����d-�ӥW�Ve�ё���^P����"%�a�ٺ���^�M�0�$"��ܓ���b���L��-��1rG��He�:w�;>te�NԤ�8`;/?��#����k��Q�Z���b����6={�	w�;l�H���4���uQL��M��vj�����|��������	3�6��\���WC،�~�5�u5Eى����+��Nm�}b��� ���E�!���e�[Hr�iB��bo4���ꈋ�,��1:�z'�ݭGca��I���n'���ZC˛uF��1q}�h�)
��ί���yi��.��YN�1��ͽ�%�^1w��G�l���s�m�����&��Y�X#����`�]��q	��q�ֻ�(�d]���%O���\�#�VPH9;<=�H���(M�S|_i4d�(�%��W�rʭ+ݬ)�{C�����s�@l�7������ꝣ�)����yF�N�71�,�����"���ط� p�;�*%����aշ�5o~�(�~��
�!�O;��Z&��:'T��e0��,Eoa��^�Z��mQ�!�8�O�k��=�`�/jRBǪ���<���?�Ϯ�V����TTX�+��r?+�j�P�	(n�z�
�y���lι�zU{��:�B2U?�ow��34Z��ؐV��;�A0�>,��4�6`�>�۬
1Q�jf(;�����#8�e�o����߾!7��-^��t\<����w3r �n�\�EQ�˘�9J�us�ϼ�# ȑ6��4���"i�Ô�ڟ|��.Y](��\��z�� S�|23��H�=3���՞��aK��ǻ�Z�256X���'�9�|��|gm+d)�h�����|,��p8���G7�6�yI�[H��2���m�PR�{�@{����l�YS�>��-Z]���:Ru��К�{Yu�b�^�\�Fk�Ȼ7�B׊�|�1\��x�jD;�h�|��u󦇀����G՚�4�>�-�3h�VR�7Ax�a���פ�V�S_�iy�el4��\�
���<Dkә{���g��]��k�t����q����H:��Ͽ��Xv�F#YS�ԙA����jv1����W>�)۫k�tK��4�t��;a)��HjZG�Z%�h��@Ck,�Hk{�D���V�et��ZY����4Ľ�J��܅�Q�(C�pY�Ƚm�ª�f��W�l$m�k�sR`��{������<�O���~�aw��a�냖0�.�QQ`��9�٦���C���X6���:׫�(�}�ڠ?i[m���W�=Gߺؾ,ø�X�P�Y���TMpM�ou/nt��K�(>��	��vJ�_8-	j*aci|BU���Q�,@\��r���N��hl��n��m(�Cq/��(�Rr܄Z���sD����x>�.��!��-�K� 尪
��v�-�j��r�L70_����~��(��A[�i��xj���4+�(z�E�x�����}��_�����B�ڒJ�+�y��*���U��򩬃��A����Y�������_�i7��c;G���t2�ʵq�q~��+J8�0�ZV��Rt�w�動�F��^U�xW�&4��a�M����=�BĪ� ��P���9=���q�0y�=�> Y�������|����VQqǦ��+1f��:5�UV�!Kf���ޡx�59�����%x�`�].7���t-Ÿ�6៸ ��@~-�ޟ3$�h�	�B����؏���u	���&�06L��j�u��ˉSy�~���gTwXU(�ABLF���������4="�����'Ϋ"IEO�_q��'��̿:d.�QH�nK<�^r9_"z���uΔ\��rv�r� �2�S	�oM	���o��ڏș��u�'���/�gHc��Ob�3p�>��!y6��m�`E��x��cٗP�4�a�=҇��0m=��U:֣7/�"oо28`�4h�C#�א"��?��
�����AWn�.X��DP���2�.p�c�5�Y�"�0�_�B��uԲX�Ɛ��0�/3��?�"]�y%A��k���Tm�bY.i���$��!���~T�z�#<2T�t�51�.쁋Z����� 3�w����T�M�n��78��*�O���	"�M��W ?o9 ��R��5���{72�^jP�ĚE�e`m.hj��=H�W��5����h��>?
f�^%����3i�Z!`���#��y��'�����Yؚ,=^ P�<b��=��񃀊|*m�LK,�vh��7Â2D��x�om�1���E�u�?���/�͘��8�SF��|��Wn�ڳ%D�o��|�#o�����PT���<�ݷd�6C���K��
�d��_��k]� MF�}=#={�Rq</V}�:@�&��<���>ɗН���7��ͣ?[,@�:o�+�܈���B��Sj�m!o�A�����~��C�u����?9�� �z� -뗦�աa� ��d��/�E�6;�^�)�\�w͐���+����BFV�V��̮��'���}c<�P��t}C�A
��U�����.�y��߷�_�)��(؈��=H�W�%�]� עb�Ў�ԡ�2YE�ʰY7	����Z��+A�ޝ��9�ʏ��`�W��5ҕ���,3	)�=rA�Ȣ3��ԣ*_���g,+�DOy�*�Ζg �y�n>RO�\�����N>����*P�n�À���4��`��@o�&
�a$���J��z
Q��Ib�R���ȞB�d��($`!�f-ܗY}�[fa�MZ��9*�ݒL��J!�W�+&��R �����CUw�sÌ�\>��E����y<��?��1�ۭ��Grp8�k�i��bLE��W���;��@�K�͵�C����DO)�Z�5�$�օ)��ޖ?,�����bc�o�/�=�n��wKV�PPSb1�+���cҀ���`��0��tc�%�(̻ȅ �X>j������["��`�	Zl��^܈�M��4��ޑk^�*�@���zN��E�;�MG�։�G�%ݕd�\�Y�:�␷S���CT���f�M�N�ʳ���T����ld*X����v)��tC�-6�����P]Yi���d	X)�����h�D����t�m��y�IQ�N2�8����M�8���\���y��T-:B(�݆+=�{enJ�y������l��e�ql�d���̓��y��pu�*��GV����;8(7nל���m.���`b��W���8��O&�gʺ���P�Y�dظ��F��ʇ�l���H@'$NAA%]i*��B��M��)4�=-��|�z�zY�B�x�����"�'؆��G�h�?`MH�$��� �dLY����b�i�������X�\�ƪ.������$�q0��A��B�)��w�HK�aW�����a�5d6�u���:��(/�u�a[������݃8a�!���5�*){L�Y=:#��{E��N#6�d"8��f���;&��D�`*��:k�d-�/8�cD���z(2���N,9I��ϵ�5�ވ5>� �f�&Ry�%�2����L
U�y�W��V�SW�k���y����d�20:d+�f�Qn꾪�T�ƛ'�!�����/��|Ճ���dk]����ݔ8��tN)G;ku0�R���o�8�i���OoE@�)�Aʡ~J�&�����,=pv�[(C���0m��<úع���