��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\���V�fnvx��ÍG_;�ȅe�~�>���9�>��Y;�0GP�5����E�57LP}T;�Qb3:�V�����M����ȃ'�5Az�	Y�-��^m&YDe�@��0N�zL�����H���;�U�~�����t_ �t��k>�D�� p�PH�!� ;-p,� � ��0��B��6IC���P�O\RBX����R8�m�Њ�V�Ѹu1�n���=���`�#�O��Y� ���G�U}�Z�ĲK�ѫ��0�-}�-)�/��ka�y��<v��O��CDm�3��"3�6vKn9��j�d#�cc�JՐh�p�Ŀ[5��<����g:̋*dF&yVf�?^�;�-�:�βҏ�����N��I��!'�G���[
3N�����0��zL���5 Mr�z��D�]�;�զn��C��O�5i�>׾ʘ�����8d�3q �*��Q�$&�Ϲ�P�e��/�~v��.뗴#�E1���>aW��$�.|�*�F���k6�
[��c�ܬ��Et �����)�d(H��*�6o�j��r�_��8�v�v4P�Q����L�(�*�Y�X¬�N��[�5J�]��,��2���*}�H"u� ������R�Ԓ�����DSn=G�c�7�N���/�ϱ�!�XE>ܺ'2,�J!��xa1Ӿ����j�VP�r��NF�>nM[�ݷ���:>���^�㭒Vho/�.+�o�ω�j^o@��o�Ack��T>P��2��+��(%���r�4�c��(e�3ܹ���T�����=���k�M=���6˫���aͣ�B-_�������~��	����7�s5n������*QMW���0(��^�U�8�v��y�DO�M�Z�~� 9����kN��2�n
N���J�u�'�K����NV2��jRl�=����kt�J'�nnOLb��j ��ryC/RFю�3�4!˜���O����3�Q�E�e�Fo��]KS㗩?'!N��l>��O�a���?��1ٱ����$I����B���?�<�-<��c��] �"�6�U���F7%.U{�txx#�z��lllO������)���}���%����+�w����l��䃷p�<=��:��z.��H���u�0�}�rw~s���K�Л�:g�]{��z��'�@o���M�$�WZ�n���)�뻣0�-֒ǁ�})b�`�mC�3���m=�!1V�����s0�U)I�j�w�bCެ��R�S)�Xؗ.<��E�Ѳ�/8��"��i�v�gLf�F")�~l��Ȼ������]�d�+��3ߑ�y�sbj�o���k�A�l�6-�H-T�}�W����j&�0hO=4ʫ�Υ᭖\G�@���5��k)%Ӹe���P�� �p�G���SEJ�y�����:E��3��kWH6c��ͿN��N�Jk>�v-�?��#>�&$<l��N6���e�n�	�G�=󴺐cG�n���V��#/[�*L��'몶M��c�\�h^P����e��u�[ꎡ �pQ������#�������4u�!/����jb&Q����_��>J�����&a�yb�J7�ou�!�#BD��e2N�_�`F�� �
��4�Hsw5��sV�&i�1�W0���9<U�0��NW�go�B�ȟ0W�T/�qGݐ��c郒PbaM�Gy�{���<���[��JvX�&T���n��~�l�}. WSD�͎��Ǻ6����J�g��Fx:Ja�ޑgV�#|��_�R���Ɛ�;0�SX~�EPq��J�X����#]��n�q���<�r����uW�g��W���N�d2�㳭�d{�JY7R�y}�`M9\<�f^������B���)d��ޒ��{���A��v6�o���r+P��:�R�C��V=@�REuf\�W�\X�{V��'Q�/�N��5���k����@��11�Ɉ)�����]�������*iw���-�ŵa8���rq~��}���<���?�Jl:.���	˄.���`Ow�Wٺ�^�z��MtGd=ߴ6�`��<9^۠�&���>�~���Y�7؆>���zsB�mjO�?���@_��L�E�}�)i�2�O��k��D��<���+�����c���f��,B��i��x�~��g���w��9q��r�2M{��~�t�"/� ��hl�7�?���x��0P;g�\l�:&+�>n��D��כt��@�e@RJ3�= Yk���4����}�B���kh@�Z��s0�(�Ӭ��ؔ7�� �������ĕTƕiq<�����?���DD(veP���e�B~���r�����\�����b-Oq� `X]^IH���(V¨�@#�\`�������3����; �Z���(a��U��\��cm��G��N�'�-�@��� w�Z��}`n���L�c�'�q�Ը�P��z����[�|�S1qK)�"tz�����!n�kJ�K@]���96\a����:X�іU��}��L_r�؜ި3�#a�R�) �}��kEӔD�e��*�՜�ߣs P~Qq���uT˃��!�g��~�b+ÉIۤ��L�M&�=����(�A��C�M�}�!���I�[@�P�g�qջY��PF*���Dz	�p�TU�"+K�g0ӽW�V�i�;�u��E�S:�s�|�g,�t�w2����e.��#|�yMk��X��80#��˿@kƘ\�^�����?b҇��[����ps�ƾ=>�-A@V�A����H��1p���=�):5b�|z]�{���cI� ��f3����A�,���,!1Z�j'�:�����?-k�Dg���7G谧��!m�����t�VO���0�QRcgB�<1��8�Ṷ�����o�������~�Q#��H;����M���
K��	�N�E*�ߎV�k|����E�����x{�z>uo	��9� �|�z�së ����rؑe=w�=ƀ_	uq�ҷ��ի'Mp8�Q���p��F��2�'kHͰ�{ �Q]������;���
T�����mk��A�p`R� �FAG�p��?׈IO�\��c���0�Ly���E�,G� f��ت��[b'~T������#���.̼F�jl2L?�GP�
�"��%su��:�H��o�-R���_��s��Ÿ������D����,������i�eGkmU�B���s�o�#.k�P>Ў�`��l$����Kj���8lKG+�W��Y5�/�x�뢹a{�x�؀��$�hg��8'&_�a�P�.�B�9���#^�sdy�M�E�������c��s��s�x{;�7�~� ��׍r[��������^� �ٰ賏��3&�k���"J��~��Bf�`H����I]�����x˖MQ�τ�2Q_���6{)v4�W���B{���KXv-�#k��C�%$J��w��ۄ�^ٌ>�y��+�UJ��t0�,�g�Y�/�[�/�"o+�Y� n�aN���2QD ;�`��xi�~]������k�"���f[N�˸I�|�����~Q����Ӯ� ��H8j��P���H�釉,��@�g� ~+L�d7�.�=ؘ-�`���|&	�oݗ� f�o��q����4?��Qe�e��9��K�Lo/S��:o��~k�8��K��צ�`S�D�W��ۇ4ǣ��=��U�W����Ѷ��E���~��Ek).��8G�a���!�v8m��ՐQ�-�H����8��L�b^ތ�֚r�It�9q�.��d�.����آ���
�L�<wQ�po����+�w�[<J��{m�V'�ķ�Uf�,#�����56��?�C�jc��ؗI@�(�Cy��ۄ{���ܼ3H��>ɧkm���\#�;��1P�4|���pq$�#���b���dF)ء��Qa}�ɸ|�(�	*�>�te���X�s���׼�n5�M�K��7��g��N�NIt�&9(�ػ=ϖ�>K6���i�hq<ʦ��K_"�lhj�&|���U��p^��6{*���vb&�'�ԍ�t[|����:���q긾�iB}�)���tG`JFl%U�u�,=tUp�#���*��g��D�if%v){��aZu?����'��J��;�%-+�cxh��U�0F|�ѱܼ_U(&|��3. ]���)*_gD,�(�l��Ľ���5WS�e6��b����c ��O�aX�Q[�І�K��G2�)jm@ΰ��Ŏ���o�~��DZ�uU�[-���*܊s�9�b�$|�K�$�؃R�-�I?]"����V�W���EC˜�~�"s�d���Ԕ/ǠK(��)���*A�"�ڔ�;p������%��R��A�d�o�%;���A�mؓ��<��ܥҘK�p^�����6�hv�Z^�[����?��g�4�ܫ�^����UDr����
Y�����n07�u�{�.�8u{{D}�*n:l��Lr�p{:����Ó� :�������n�W��ε�ц'y�0y�T���&���ȇXS�Fxm߁$��;�}�����ВOmR�a�\�Ч��`�a	�4<��_�=�Gv�,
+f�ז�X���[�@�jY�h_Q@ˮ=����ܟ<mݛ]PAJ��Ԭn�K �o3�o��l���i�8�3y���[X4�W��)J��3�X�2�b�π>�k�X}�9�`�����V#_�&�P���(��ϊ�wk�ޕ��=�n����{ɴ۝�9��C��*!���Ne򎹭z4��*����֟��� ��_�yÜݧ�6GF�}p��Ku0��zp'ϴt�>=��(H�c�&���S�'��s��JZ������e'A��N41�05��K5��T�~H��N,�c�Mp���ǆ�Ia�8q��6�Bƨ.wLq$���zy�O�V;&�{G��⑷b���M�i�P܌�O��_�\]�%=�6�e�'̴���������T���*Íez�u� ,bS֪ �U�J~1�#5�t��g�I���.ĢwZ���q��'�ŭ��ud�<K�!���j���z�׼�+�d����?��s:�jG����&��{�2�B�P���绰�&�X nzh�Ɩ�'>��6H��@2�a���W�Rf�i��M<�_<1���G�d�߯Ꙃ��T�o�q�J�Q�\[��8�� 9�d^���%�Oa��o�a"Sm0�G!�M��\Be�`���!(���B�?������{�"G�����_\�`fX/o2�qlg H�C�� �9k� ��8�8�X��4�FH�$x��B�(�ܻ6+�W?����VH,h��	�C�ޥ&��Ȣk��ͽq�T
�_�.���f�U$%vyc�r�1>�G�2z����� �U���"�L9���Œ������ƍ�����1�V��� C%�XO��=�特\�OR��IA��x���z�\/\�U]�{�=�|L�����P��p�m��^����x���٢�u�;�6�ix��ƀ����2��e�)e;�? V�}���a�,�D�W{�.�W��(����=6i�>]h���JӞ@�����Q���h��1d�&(b�y]���ۂ�;�
�U�_Ôo��P��5��U�G�q۫�ݶ':����B�
�؟�e0�s[�n3�ϕ�"RQZQ�n��.9���Ҝ]�G��L�[b��80蝿��_�>0il�z\_6��]#��|�gK��1>25�f~���4_4 +�o�\���<��<sH3� 5=g��{�oc�XU�^��a����O�{�����D2F+_��[�'sH��I4 WeI}�8��[I_�n�ަ�[��]NPh4���dfp ����$�B� ��"n.������\?[��dɟ��`��6�
�����ۥ*Zq�-c��U�!xrē�ӂgΡ�)M�wLS�	+34%�� �c�ğ������o�\�F��w���w�x�6A��TW/a|�!2l��v@�� .��o�
�X��|�/i�3����BG�]^�����L�K�cT�ʱF~�I�#$����YR��J�ɑZ"�\��)x���0E'�a�@�w�k��qYW�-�L[3-} �芘��{�NX�
{k�b<Ɔʈ��)Y��N}V�$ʖ�'lw��S5���Ua��0N\w<�N$282�a�]���R��B6(~N�F̜�utVm�eO�NK$\#����Y񯧆?��J��+�nBB����X�� ���[L9#�^`�R��<�^��E;�;��^�e���"4 ��a�c�0��A#q����f�홉#� �F���;���0��]|�;�9Թ��;���=�gdPu!���}�	�U��,���x��d�j�!��X:�6��Ȁ�V��d),)-��4�3}�������BƸT��bN,�x��H_ ��ȷ/����
#:����}ݴ?L�j"CA�6�Ġ}����x�gW����~���N^�q�G��6�!P��J�a�0N�&���A����\��qB������<6ŧ����f�0I���åV���3k�eYS�4�O�@9���G���Jd�FK9ڸ��Ts���!#xt�5�?�l<�����ח�ׁ�j�:
_��֗̂��F1���|q�h��y0 �H%�Ω�[�,�V :�R�,e>*P���|��Gt�q�j��>Q��˳�e)	�f���L�I?85�tA�����L�A|J0�iq����pCx����=`����yI�'/G�ŠůO�s�V��ǎʠsq@�M����Bh��V�`�x��2���;9��\�~��PяSh�DԄ0B�����^��	Ng��܅U=�z���ʗ��4h�p�Y���~o�Tp�5���h)�M� �d�� +l1��Y|0�}�����a����qq搱�*Q^����-�]XCB��L�K]a'iD�f�6N%R6��iP��0^=�ƭp&�+b��R<)g�����ђ13�-���qN{�8cL�<4J������$}E�ֈ�=��'ls8��)Pԯ�����>�k�cl�Ŭ
m#���r�]�<Qo��(Rb�*��Y�bH�t��LS&/_�o���-�k���*���@LR�h���ǟ$�)WTaD�o��ɑ��Ė}�� ��&�QL/���:&��H�M��;���f��rbf���HOUV���=�^}1c@���w�aK���p�h|mn��*vq�.�u��kS^�"@�=�Hm�3�/k���WunN����n1�fTj�E��B�AiR~�^�D}��kAm����@a�Z�r���漙N��A9Ds�a܀q���\
29�<e׫���şT�d�v����C�<��8�
�-�u䟴i3c�v9�
i �i�l��N&wJ�K�8d�w�0��v�Q��2�r�`�4��ဆ� ���?Z��S�8��S���ȀR�&�0�'��C+,�x��'�
c��`���&?����;'�ۛ��W9��o�l��TD�lm�~Q�$傧kƑ �Jj�����y�5����n�?� � %�&��|3$rP�~z�/!�Y��<c[4iܿ�݋�`>���+/�)Š={"�W��<���.�iӳ�g�·�-��F�~x,vC�I9��ӡx�T`��p�ע"a{����V��*ΑbY/k�q�N}������<��m����s��
��HА�����#�k��N�p��n3y���Y����C����t��{ԃ	��3	���{���a��vwA�(�e�>�00}_^�3��K�_�K�7M�����t�΀ʡ�ip�5W�2���?vX��N�1�l�]~&d�-T������� �u���������2�Z�]mn���Z���ږ_������j`:I�a�p���/#N��6��a9�喙��zk�U��q(p�R�y*��=�i'�)�=2��#�V9�����&�xeph|Hd�����������ʙ^&Ґgm}��J�a/����+b%k)��y(8���hǐ9���0�C���횁�xD@A�(�k�w���C$��N�� �X���d�M�XR�狾7-�AAmi�[�!q����(�k��b�XbuoM�KĈ��(��������e��v[���W��D{.����~)�,�_9iB�O���T]-2�p1���H+��+w z�~�� �0lB6�!����.�ɹ�i`��%����?����<�C2Q*DoW�iH�'�c2�`�<����t�0ɑx�������O�N�,���6:+�%�R�4�����5�'i����?`���A��v��dŠ�s����S�+=��k�FO ��x�Y����66��D� �	��r��E��3��~8��3�� �b�{�1�8�YԹ�%�"!�8O�P����w4���|+�@_���2�t	����j���)q�vk�4�fA�vÅ6�9��I -61�h�L�6��}P���FΫֺ��V�'Qp��=�ݵ(</L���Bm%�Y�"�X�{��X��[�1���(�<&j�o��g%]����G���漴�r�'�C���R��q����$pG����Ѻ�;|���|�+�?���\@����m�5�q�
�e(�����[%ɾ��W' ��f�:�����.�v���|A1���{���w�:���V�S*Ph�ɩ�p���c-��< �ɓ I�g�W�|"��-ea.ZA��E�/aD㽍�X�f����6��ܥh��O�Pn�<�c�Tj��F���`��'a1�u����٩3��$z'Ә����΄��Q\\j�~ r��~M~h.y��?��SQĸ�(7Q����L�<��$�4ңL�#p���<Ӡk�,n�m��D�y�����3��yÜg��a�F�4�qL\09O�ϤA=v�W����o?y	�k<u�*i}!�B>߇3�.cy+ӡ��w�=#��9c ��"R�2j`����Lo�}զ��휋:Y�.)1읰�){�� ���V����vH��ω�������⎯S��*�_���o����Za�:�D�KO����Y�n4r�������#�2/�e<�9��:3I�	5ʃ�"��k��ߞ�|��;�7C�Xq6�S�+S��+�Y�Xj��ެθ$7K���3��U|����%*��:M� ���{�S�0�������T����|yfHI�D���ǩxuA�OIs�m��K��J���9v��^H��Q�n'�q8�P���)9!����zm����ϯԋr�a����Nq���(�������A�oX����X&�/������螪��֓
D:�q�����,aVom���u��o!���|��̰g#��Hq�k��M�1�<���FkX��i�@��X`�Rz!�+�Y�(P3�m����:6pE"�pi`�CIˣ���s�z˃��q�"6����(�ģ����?a��w�q&_�j�H���]�K ���kݖwL%W�� <�x�1*�*E�e0J�'J;���~m����k���x�h�wTy3wp$�ۖ���ȅ�����#0b�H�#z�ͳ�!��T����k6]HB�|b���Nh���*�G��;W�P�#6)�s��-� J'L�u�`餸˟�)46в�@���89���`L�G �'9c3�S9R5�rk��c�����)�_�]g�� �y6�V�F!7�RҢ���(*��o���@���ZP-����yb_��\�	�pU��c�O:TH�[nN��6�]�M/���r�,3�Q$��œ�Br���j�Uo:|�G�gNvvT�ޢ�ݓH`��>����$�8�Rc�}�)v��-8�S�7�E Ke�j!5z�W��Ӱ��Z�/ω=?Aq#����E�}J�L�����xߗoKRҳ��������-=��)��I9�L�ES�C\��v?A��3���c�و����Kg9�h��a��/(�D�,�L�/�.�[���j��!BS��^7�IA�N��݊M�}���_!��jE�d�J�?�����%��cq�HϷ��97Y�!������,:wg��AkD�
����a�,�%ľ��G���g�qU߉E�D�Od���魀�34�#is��+s����e�s��Er��	��T�6j�bd}(P��K[�@F�C��m !Y��_H�e����.��Y�=V�n����A'��lNߧ��t��Cd|�ܡ��e�@z���aM��9OZN-�A��I��ȭ_��4�5	 ϊ�y)$����e��/��\�h�/^0�*��R�u�_+?~.����ES)4�#�Mu����h�6����骉��8У����b�Ǔ�'
�M8�$Ҵ����D����㙍9�b_��@,���C��f�u�J}�Q�Tp����6�;�!)z�~�Pm����q��]�Sॵ���d��<+F�S)a�̙kޕ�M�	
VW�T�[��2��d�.&����J\1T%Sjp��Ru�9(�u��,ٹUdr��sH��Od��G��z�d+�J�{F��OQ�5��Kz���_�')u�>ɂ�>�.o�g��Mj�c@L�5�{�ϫ���p����h<`��8{�๯��*��H�F|��j$P�Ii�!@A��Ptt�����<�� ��0G�ݢ0�h�U�{iӍFnD^��<(��ހ���h� h������ oÙd�^8�٣��A6�&�aJ�@�#_O\W:d㌒� � ���lE����SCﺒA��/?V�	�{��p�H�.xfԛ�B�}�e�U�4P���*�DS�=i2R���?.�Ȏ��y:̛~@pw�7jUW_��-ʇc>�i/r�	��Ppf���@q	�(�p��==��Ԓ�?	������=CS2���XM�@�dU��)	X�s��ꇢ�����.�>?$�\G�)0�d��;�/�p���=�r_Vnc�bXO#�(���uR"�],�Y��\���#�ʙ�:��Բ�����9��&
�'s�{�+���]l�7�y��%����؋H�&0�z�Ւ�J�ax��s��3���TLhG��`�D84ܧ�A��T�q�r%��r��V�	O��@0�Y�Ko���jJ��u#���Y�퉗�M�݁{��ƹ��Vld�4���@�o��`e�~ݮ)4��f�e�,q�'(�ͱ�Z�R/�y5]�Nx�*.Y�uğ9���-�Pp˭b�Ly �8��myT�]֌��b�9B�=�*?,��psycs�-N���s�5M��^�P�Ժ,�Z�{ӎ(�YU[ܛ3%S�jmN㎃,�:5����9�?�N�{��<O��,�k���6������'���������e�'���[u���T�
ݎ l^�d�\d���9z�U5��}��&�%k�Xiiv�cC���M��~Yg�B5���ws}�`����l���x/�R�Q?Y�ծB��,@,ֲ;�_J��,'�y��Tw9���Y�|��-�"��V5��)�;r�j;ڴ�Q���A��Q-"�ʕ��M<�1�(˛y!$W㹁^�Vn�]�'%��c����2A�X!�ߟ�P����z��F�u0��G�A��F/׎�]��yg�\�l2��\��r��LRi�����hq��[>WR��5�+��J�V=�N�����K DL�~��(Eh #|F<�Vw��!�����یYI����
K��WZU�<��1ԫϺNR	APb<ZFpM��XZ"Jh���~d�}�';�?rNp���@��D|�[&mG��kekf|�<�k�#]x���d�E84W�1���̛�'�d^ޭe4�@�iT�1p<�����̂Q��\�<���{QɏE7.�ӞINnV��N�!�Hs$�������1`��Q���xo�c�a��7������"1�i�7^3�k���>tL`�-A^c��b
$�.A�1����A�L�C���/2�$x�JJ��E��՝�2��cvA�a���ݥ�fmM�v�U#����m��6t�����o�A��]���c�:�������֦����K?��acoߎ��j�
�n�J�ܠ����@=)A�'�_N�[���)8h��6�6���7:����3���ē�
<`��%�X�#�cR��p���렽"�OS.��2ŋ����������~NX�r@��Ņ��ߪW�pٜ�j���p#�%+�JW�j��	gtn�˷\��.uN@��v�W���=�+������%d�!�C:)�@C˘į�RY.��h��Dy7���� ႌ+#�y��d�u����>*E�~Ç�0�4��
�֛�;�,�|�N}N���� ��lͯ�����.���{~��S�O>��{����~��沈�L^��Q���R�R�o�*m���Wm����_ Xi�ҲYO!/Re���nփ�	S�}*�\j�ʜ���	Oq�*�܆�vp��_݉�P�'Ur� �����)��be1'a1�I^����� �Q�2z���>���x�h��7��l�	S��%��Gp2��Njމ<�:�$-Q���`,��5�֜>{��W7$��ibd���#��s�lJ�{����r�l�����eQ%��+e���D�������
=j���ښ�z�S*���D�+�9�,6{j�T���=��Z6|E�/��g5T�c���H�a%*ɩW4�A^�	ó&[�(Z�������{{TX=�0I�({o?���y,�6w�UG��Μ�}.���hGV9�'�: ���j�ʬ���]�~�/ �1��I��NQ��P�%��D�{������H����zf>��)��[>��'ަ�������n�æY#)��b�N�M�tIl��G~�]8��x�mM�Ѝ��[��������Y0�"̢c��z��ŮKW����r_a�ҥ��єYF�ʟ�"�AI��3������p��X���Ds�t5��>:V�`�_6/�yUg���$A�	�+xkQq�Ddu�����5Y^��#����"��3j���'~������J}�j	��8zn�Jd?�0s�R�f2��j)��^8d5K��B"�GBs��&�d�B[����#"�~"~Qj�����@��␢���0r����E�@W0��t��4�{2K��ɶC�MGVoҞ���~�car�K��N\s���0K[�ȬC��3��b
�,��sqv|�������Jo�F	8>g'�:d8����|��|_��7��S#{�8��#M4�V#��>�98�e%���Iݝ|b���K�)D2c���c��D��9�^�4������)��}qs|�SX�6NQ��g�(ƍ�:�
�xx���W.BK�K���z;��
�T��h��ܧ�o㼭�M>�׃#�h���k�A�ʎ5��&fL�t>YI+A�mu�I�*ǭR�^9�4�M�j��_��\��ma��8ߔ�7��5�~�ӆH�p?[�3�5t3�(�"[Ȋp*{���{n`4�Ѐz����P��[�vd��Lg·�8�|! x <�D�66f���}<�����B�9x����$�¬pXf\����3Y�n��Gp� 1t�Uϙ�A�Ӵ�'=CMG�Q�s�yg�ԆѪ�I��;x�1�B��Y�;�<�
&�ۚl�=��Sj-O��K|,��ep�����?�Ux�x�ktCS\��4�������D�&[�;���ݐ#}LZ�m�ѷCQۙFTj�����rx�5�ݕ�~p��&���ԡ��P���("��,9��������.�a�����Td���)��8�)��I����)y��K��s�zρ�4L��Qk��9@a�P�m���^[O��Y;����S�E��Y�S��1e�5˭K|bè�^�Z9�fL��ff�̍^��N>cc��7�>�^�&�U�͢^�8��͓+M\P}}�k� n=·D0��E�i@ '~
�+�����?7Ħ	�|ئ*DZ�M<L}�w�ѧiL�q(�+����ï�.Ss97kD�_�[-�ɥ=L.�;!�=6_���^��ѓ����� �{f@]����z菘0�W���5S�Xl��Q�R����S_�c��7OHҠ���xo�i��a�C�$ʞ�y�z��چP��4���	i%a�\�C-W ��� ��R��>����X�/��[.&��OS�<o6gU�����ՓWD/(z���"7S�X�����_W��A���_R#�T��0w祒Lj`}@�/j!W��#H�K�XS�탱�@������V�a=�im��	��ba�1)j��E�*.�����3�N�f��s�n>[��Z��)�$�������̠+U,k�ѕ���0�3V&���x��ɤr�2��M
�h�R�B �������l�9�G�/q��c�A��f] J-��ʩ����A���6frM�B��ޱ�9�tӂ
Y=
1R�uد;�NjH��c=�3��&ˁ�e�\�����7�"���+8*@Z���Q��6c}�/���d�i1�ZE�-D�L@�Q����s� �x�������xU��1�{������D����M'a)=���',�ɾ��j��C~��G����M�Ym*�|~&ď� B"ˑn.W�_"~Ǹx�`�_�!�����[D0�o�"��!_�=�&=G5 �Q��K��_m% )%��lB4��-�Z`!�{B ���K}m��=�bH9�>�qM��V����;&��˚4�S�nA-dP������k0�L�E��qd��@>�jh�H��&�9��R�@.�>���]SoX���6�����֞��$\����P}��r�+D׷6����G�8�'4)��8u�d]�⊢�|W��I4���p��m� �����i��G���:�������|�P��C^�~���(�i^��3%g<��O�v֛�1�
q�Lt���~�l��p;�� �l��N)�cx��e�c|�o�J��c�=�̩f�
V���<h�'��J6�e�^�$u�#H�ZX��K�
9���d�d⣶��a1������HY�F�x!+5-L��FR��a��r�ϱ)��M6x���SBs�5ߍż���f��.E#14��fy��b3#�rv6�);XC��/�A5jdrf��<�o���jWR���)�[�5!���R�C��&z��m�c�B#�!##��<sp����%�ޚ�[?\h�
�<�_..��d�,�c���d���O�݃g�����g�l�+���$#�mAOD�_{kw��?���Y�m=Ʌ���n�?��Nk`0��ϝi��bc���ؗ��w�"Z������Q�O��y�ƣ���E��cV��j��]��;o�����Մ(�����Y��.��+]��0	SyZ �8gY]V=黜���T}�Dh��S�3�j�lD��������]I�D}FIkc�c%��H{�f��v��E�xQ����x[�:�n�׮�mɃn:�b��2�Šj֯�K%��cw�Bh�g$w�ӕ�¡vhiN;�N���>������@/ov�'@Gt�$ynH�.������ֹ������mS��v>�ˀ��K»���:��Q�IrBb�Mky�~�Qz���ŀ`Hg���R���$�2󿨩Żڹv]�~P4��)��j���r+��5����|��zDH���B,u�@Y�t��m�m��z��=x��R
 �~zDI� �pf�w���Rޚְ�P�;�i�'�Uד*����_m
�z ��;�����^4?F�
#]<�ӾN��U�f>�䎡y�JR<�� ��
"=��	%K��#�!	�qf������1RtnŠ,ء,]�Qv�9 �+��[��Wt�g���oQ��ߪ��5'�ܤ_�/�ֆb�YW������ԁ����W���?�k�C|g���o�Q(������Y�|��&�a�R,Z���`���&���9.��@����P��m��K������/3�Ş���Hz4\Ҟ�2��|�}A�z���%���lD�m°�j�>���ԙ �P#��X������hcSDAzj��f�)���v���N�-$xs�]���y���RT�#�c\���Ty��B4pQc��zQ"�;^��#T'���������Lr�??85�t~�B�P������I\nq:vQ�ݒ�̨�Eɿx�\^�(��#K>	���"��8��ք1�W�-S�u.�_�mj��c�҇\>9ƄW��tp-D]�Sj&��X
�Ok+��ٌz��>?�s$�=q����$�{�p<۝��(!����/��&u�Ca���!:�/E��%'��G��TF��7��:������)&���}]����	�:���2�� �O�w��T$$?���a1�,��􈍁u·"�z�Z����8x	�`�k��c����̋3�7Z�ap�@���㐲�d��h��-3X��Y�/`�\���w���[���n	�7c��r��XD�N騯#�cB�!$�6��@C�CZ?ov����@�~�uyt~�P����Kԏ'L�)�(�@��V�20҉��֑��|�}�~��$3UC�X��O{4��83����8��tз���% ��N���r�t����|��|��t_ /�5%�n�(����Xp�����qZK��pC�X���j�4R��C�acA�}���Y?骨<0B^��>��~M�IID�կʲ�:$��yRr~Ĩ.�qU�a9i8̋r(?�DUw��jAr���u�	;�p�~���+�o^��W/s���<M�Ŵ�k��)�;��[�[c��-�H��L�i4|AEqx�������@]�>�BAt��$ɯ��?�`O��g�+=a���(Q�@�4�iWp ���K���GJ������3R���wz�򨻚��U���%���7�@k�;��s߆#?�3�Ug�S�$d�tG]u�7���z��_����͋�X�f����x�Z��>�ZL��Q�kƺ� ��,�8	�]='(G�~���Lv�p�s f&r��1��,���`�F��p�����-q>7]�Fr���i���ܣ��I��՚�1q�x�[x�m�75�f�,י�,�>�w���q�E�ksɔ��Y+�	ȁ����=9Dҥ9�`����B�U��j�8��C�B?$���Q x������[Ŕ�ĩ`��z��*��\ٚ��5���������TNFI�<^�B���J�l����I9�5���",�����h�+��-9�S�ZOxw�?���P=7*XԾ"��R�Jj(�-4!��"��'�,V]4�A۱�V��a����p��.ԧ� X�s(��������o��+�yL�gv�Z�h8)�^��^�D���N&��ys��J����Y�^�io�XQ�<S
0�\�#��G�%=,��o�1�⒓Bv��\��X�0R�E��%��#��Ԅ��:��纫փ38��g_��FENd�Lr����
J��H`*���f��z�R�;�I)ɣ����\	��)�LK�>���$��!���B_O������i�Qen!�q�9։��s0��Q~��0�!���BAUwk_�0�%���tW���|����t�o��s���~�S�a���ɔ"#�ݔ,_�3��L@,1�ߝ[�?D��^�u�Ҟ4t�+���ҟ���o�_c�V�'B�DPFB��P�����hI,#WYC2h�f�����*��de�3{d��~�Ӎ�4dJ!&s/[R�C�Ǳ!�e�.	�!9O���tq�!�IX604r��2:=ȓ�?�Sү����Ӳ�:0�\�v�E�@>�
���y#$R�6?�I�Q"�Ɗ,8~���+�"�8�5���Y�A�9����AC<�U�نs���-6��iV����!S(B?cA?G(j_���r��ۮ]{�Һq��" 2C]|�}	bpV��|܏����^�Y�d��r(`M�*�������¹�3,zX� s�"j����܅������Bv�&��hU-�`Yb�]D�@"�T�4N;>X��,K!zO��6rI���M�>���������^�V�������y���:+�x��J��B�"�Ц�%�/�T6�+F�:����@�����S��d`Q�A�9E<&��燷�l68�	���&K�v���0���.W�����K�Xk!i�7���Er��klUө1SǞ.p3ax�U3�D����SQ'�P��6��:kt#�i��W���d�]>5~�|�:�1ɉ����!��U�(K��Z���-�����Ҩ����L�Bv�'�gh��d��N�!Z������|�ﲧ<Y���E)�vońo�7e��\���b�O���+��h�h�I�)�
җQ�=�����5�4Z�Lc�~8���FKH
Z�V��]ch%�&Ԕ��>�tV���ć{{�<L��@} <�#���:�=cv�bJ��L$}�օ�����p���h���Cn$��@Hv8S��-��S�J{o��9{���W˵%���e;��(xH�U%z|� �Əa76:����^�5.�F��u��v=�/����3�.��Rqi�f$ �q4V�� �q>Ж���9�_�z�����o�C2�7m�aU�d���v-L����˭9��e�Uq��k����W��U��݌�?���j7Px�닆����B�g����S�q%�:j1�䏱��/��s���bO��Ƈ�}���@�0>ͩB�i�[��y�P��=¿�a��,�(o}���O�Z�P����)���-g@�R��������0L��E��pNBz
oH�J�<�g�ճ����@4h�+Z5�FB���h.�Y%�#5���Ca��ph��6�\�q�Zk��Z�Ͷ�[c�D`�>���S�D1<)���]�/
�4ظ/�+|l���t�"�-�����N���}�ǒ�H�'��дw����d1g�x�=���7�{?�����k��Z��S�&M\��>X�},4΁�����]�B0�i��o�WI���.�/�d�#�2貗vXW�PF����>\S�����Mq?z�	Z�){e����B?�[�Ǆ��T}�fܬ�TK�[��d
��ՙ�Λ��������Μ6��K�nۈ�����R6U�1
��E��v�G⹉.I��J{U���3+�@O�=��ñ.t��70�{�&llj?�6�����d�r���OI�q]߷l�]kKrV� s%t\h�oV�����)���M{�0�&� �恐Р���V".޵�<��<y4�/̼�=��Fym�P�����G6H =��+�����2�5���&�R�v|�)dh��!W��-��Ic��FV< �8 �$�ZJD�e<��$x>mRb0�S�����`'W̟��;��<�q
�4Sɨ�nE&&���
��=gK�GG�R�����b��dޱ7S��yby�����<�ň�QW�G� �⛊���ʭ�GJ��2�oR6Q R�$�D�om�����= .�(l~��r7�J�Ƒ�	����iE��O9�W��KN6 H�
�1.jL������WqF%j@0�v��FBA�����nv�K����1�WX�ӃA��LP͑�����.���T��)r6J?7�!����z�]���A���^)�&���|p�E�B@[ڄiXԴ����1��	�b^����Qs�w
-��ڌ�c�E��@2-`	�OK��@��TS8�\(d�h_HM����KI����YcE��L������/ Q��rk!���񍉋	0�ֵn$*#%���< �Ղ��B�.�}����������^��x�̻��H5*���*Ǥ�\��Y��9g_i�\���6�y��M��z�7�rDw���f�tcB���c�!M��z��&�d�3�PQxV{��e�3?G����/.��X���ۘL�quL�a�O�P�Vw$(�<R1�5c ���^���f��v���$������]��S�f��i��N��YƩi�`�29��^�B!c=���pzPR:PL�H��I�tK类�=^��%���:���!�w+�$��Q��4VLX��`�6V`����??�\��r�?��P��~�[&�H�׮L�~����I�_-E����u���ƈ�(ai���:뾕���\R��kۡ��6�u�"�����5Ǎ��ƣO,Vt�n�jJ��j\���������B����A͋�W��r��	��� ���)�礟@��֮^�G݆�)���a�����묱x����ˣ�ٟ�L��P��.�v=BG�D��S>�&��_�FU[͕Q~��t���8U$t�n���0;~�V�^��y�yMe�X\�V�ZJG���tqwfώA?��/�_�����MX�����Ի�� \-�]7�T2����M$ixx����4M�C���c�y��zIgLu]��x)�����ٓ��R�w�тݤ�R�4�Z����>U�m��\��)�7�B|�����,K=� d��L�h��Il�g%�T�K��-�W��V (�F��V V��{k�����:vN]&��J�Q�x���g�(/������6q�� bQ�"
��� MN��VZ��%�-g�E\k3�8�f韁s"�{��}��LAY[�x�����dJI�F�<`eXgĥ�4~֕����@�x`�񜬽�k}m�_�G2��7p�m�l:�w�U���Ғr�n�ӿG}n�*,�x�]�Hq.R���_y���b؆�8�L^����T�>���`���O=�m��M�ע�	/w��O���k�4�ѻ��l���2�ï~K��[�Vg���o#<ô��ެ�]-9Wco��)A_Y�;Vf�,�.�	�Q d���~��#{����9.�~.���53FZ�Il��K%�Jh[erc��lrTR�;A:�Ҙ� �\�J�V:���#O�jZ��k8�#�?ú�$�9��s>��gO�����%2�[��!z2Ny�����=;�v۰\���3ބ]�<P������Q8����u �skP�Az�)��j�!�y�_RX8֝�u�������؇�G���i	�0h\��=�L�!C6�.?��zJ���
@�,�9?5����M����S.F*
Mى�	޳E#�R�󽓀��$2l���Px}p�57D�6c��Րw��
�nS�	�L�w��x� -�B��֞��gq�On�#z���d��@Y4�a��1��9�뱞9�l�7�4j���أV-/��F$������`�l&�5� �y6���8���i��8�b�z�# q˟C���Md�K/?�|��]}���w��{_ߘ
Hw��Hr��w�i�+��/tS�U��acG=���qʙ��.+�	�?��!���P�X�d��Q�HW�UD��9�b�����
I��/F�Ӵ� ��0?�"�2��G�Q�5��uD���B��y1�q�g�3{�k�e�K,B���9�e��pʷ�V6��a�~��bç$�W$�Y���k�(��#L�����ueJnq%W��^�c+��B	�a�H�WM���sR��pW~*��]��4�H(���T����ց��e���.ٖ�	��\/F^C�ve�i,<������O�A�/#D�%;-k��h���Ǿ_��$�q-7S!���%J�fs5�SCϘ}KL��63aIף��hp��c<@�$��ˡ��f��=�µ���Qg�
 �1f��h�pqB�W7�Yzn�/
��e�~�Il�c��ap1H��0����y��hc����L��n_"=u��E2��Uӏ=E1Ŧ���������v��ё�����J��nYh�K�lv��c���9��(F��7_������F�TH~M8lc�(�����!~�T�z�<"O��L���է�
�0F�Gr�F�әXC�GѲ��4���O�nά��+������VFk�C.XM̥>6����ͭ��"KvG�(H��'P
0�{.�8
\��G����;�S}+�|&�V�B��)j�jUr^p\)��ޞ��@N�9}d��G���4�[�[W�Y�y��\�+���]vg,ƞ��e� �kc�귫���Uo[_ύ��l�A)F>�����8�[��1o�1�6� �񋩲��n_�mo���D�4L������� F��u�H�|�~[���Q��U��j��t9VQ��\�3ubEk�OA��Q��\K���3�4$�O���Ɋ%��Z�(n��Rְ������M���h���'!�a�?ƹӴ��¶$���5�2Y��K]BXZ�������� yIT<:"�͸&<<�
���Kv�GTę�op�4����<�jXVi�~�%A7)�q���³ɁE`�,	nrr,.T�^6o��Z��5��מ�V�H��+�uKb����ɋJ2(��{���Pu&�P_��+�){�nV=�Yj�����H+�u*��T@B~�h0HĦTUoޡ���(
�Sh��g|�QgO�c�xYZ��	���8ŔP̟���U�����#��9��p��X/8!�<iw<����_�.�&5/�E�B�&!;�ƾ���]K�6��E�F�h����c6/Ã��������|E�7.�-^�^g�� �@ ,^�z
�p��1a��3���Z��qx0i��;?�y��{�Tzr\.+@
7�2�,�M?/��|5ؚ���_U���_�x'�'����B�9�lI|�-&��j�f+��!���$��PI���'�K�v�Y!���s�MVȖ�5P�(���.�D\N�C���1�rG���1�b��� fz��ja�h� fR�y��B��́I4��6�[ac\�gɑ��!2P�Y8�uM��1}aq�S# ���gSyt:�/'�!�X_0���^����]�RoI�x,�n̳��QVXq�͈1I���)�l��M����aL^�hC�>2:w>� Dm]�9G��ǵ�F���vXH��h���Ut�w�AO$��.rǡ}R
�\�
L⹂e���}@���/�h�fdMD�?s�8�Dղ)kx��jZ�s�8�\E����	#�f׍mȠ��4н)�8���ݦ�dQd��G�Ҽ��-mC�$d;���̄�* 5��=.����p��;����ʪ�X0��Q�VhZ��Z��Ep�����s���j�����)k�0�.��V�!p_�30���^�GTsz�{*��,I���}U�:���9b8��E����ע��&�;�p�#�8}��~���l���[�Kqt�hKVcTJ���`q��L�q��80T������7�9:��CˢgW"*��Ao������y$>�j��9����}f����Q�%���8��b�i��Tm��j0{4�Y��y �����I�RԘ��!7���[+�{�}K��U������b��p��8����l @9�׎9�f~�`R����h[.h\pM�s�/@<�'�M���'��+���+s7�з�/�Q'(����>��F!>�<�Zߙd4	��'$�G6�l��*<eˁ�=�16v%<	#p�VF�}F�Ką�#M�0�m�+���Jfr숿�"Y�v3	�*�1e�2}��[Ǳ����1�DW�p۸	Hs��mcR�������ⱋ�G���=�,h/)eSs偣聢�j����R�&�k��vq���_�E�S�@0�g���$����"��Ҽ@�Ĳ�q��yn]F���G����;��-v&n�}��!s5���O�#��]෌��H-~C@���H*B���E����C7&
���ŧp�*����	裸�t��[M̑�ۢ���Y
A�f�Љ��A��&��މ	 V�^������.ܾ�ҿK���Rw�mM��в�ZE�1ʌҾ�쐅�`��49s�����Lu ��{e)�c��8��<0Ѧ�	t~#~��~r�â�u�Z�l9���JR?�� �֙97	�(j��f��`'��W��K!oU
��(�ōA4���a%��(�Ey�#1���0)Ig�MF��RM*q</80��m�	�oTϜ�����8Y�H}q���G?ۻ�;�;a<8'��N�1�<�hx-x���.�6ۨ��vd^�:M�DG4`���\e{ŧp��В�W@Z�P�yc���C�il���	G)�TN[�9L/����[�d�0W鱢�9�G{8�i5�)�b�TF!��<~���Pk�C�920�w�g��A���\�>�(���
a��q�6�`(dt��v�1V'������X���E�knbE�#��'���=r�J�H\�謻������3H�~j"�Ɓ�!-����tR�S/@]��f��J)oI�%/�v�ӻez��)�*K��5�U��!l��х?<�����Q�'Ŋ��WK4�v3���A�.V�b�L�<��k�*5�cwݱ�*G�y�\�[�(]���� F�)QU�O�o�?>�25<�e�\�b���k�	�H�k\��w_yʠ�':�x :c��X��@�v]���^38mt
d��P>��L���?.@��%!��;;B�)�Q5� 8�h��뭈�,z��������!�Ɗ� �Ҥw�-�3�
D�
?���Kyx�2���VwL�J*)�wc���+���#LBXaU��������Kv��~b��G���
+�g!��d��}iHx>G����U"�adc��7��vl+ηt����X�EVe0E������b�E㓛��g�↼{|tY-�S���L�^�C����N�Xf�0���e��
$�7JD\㠗�8`��WGC�Hd�6˘I�)ϙ���B���h(z}F~��!J�B�OU�z�.y���x������ȟ�Fԕ�c�@�Th�E���T!�s��]Yp�@���r���{$<Ч��9��o����@�-��=�oNl}z�l��o�l2���v��ؤ�����VTz��\�br_E���L��گ�Y䔋�1�c3%��s-��
ѩ«��穟P�A�^0-��?A�R��h�3�!����m�p�v�t�-j�\���=�a��՟��r?�Ѫ��!܄�~�gIY�R����	\�A	��1�!yZ-GUn�E]�.BT_�Ci�*ps	�.��'q{�Y��̶F��eN�޶Y�1��MJG,(���S��B�Ȩ��k����	��sC"n_,�?�>j���7�5�R"�{�Y�#9��|a�"��S���Uu*���HEܖ�e�53%��fͻ�����i�����/�q]xD�6�:b�U��Vȼ�^_Eh-�;��z_3�$=��>��e~f;����3�]�)2��5���]f��&�_�-�*�R�5` �kj�F#ȃhUB�X�	f�Ϗ~��
!��9!��,����h�{���+�~�Q��r�`?�nP���h6N���6�'C�l�%7��1!��u*�'
�ḛ���x�����SL�5�����1FHp�3�<D�Y���]�ђ��� �pW��v�������|P�3�6�CkS��(�?������	'�Z�\��m�蔒W���J�,�!� a���ѐ:�$Ƿ}���uY����
+
��J�\ �%�d�)"E08����	�\��UX�!��a�y��L}^1T͈�u�9:Ez������t53 r�c#�_�W���id+��ޓJ�B��=``��C��ӣ��^������,Dų|0�#�Y��%Ao���ǂ^#���Ej�s8��`��S�o\��;琄�E�Ǝ"�%7�2�o����٤������t�چFV�ǁ�*���_i��_�X�y�i�?^�a���Fϕ�
�+�-z�l4wd>�j"�&����׮	&����H�D�j�i�v��kX��c�n5�5�lq�~?W�QD��~���\S��!z��1����+�l�%x���Lԗ�'~3/�ְ�//"z۸���7!�IF��/�L���t;�����o��oQ?%7�Zn�Şz���9Wu&D�	SS|K�=�O���$�Um�Ņ�Q�!D԰�&�b���l��뢯��� h���?P?�!��1?N7h�5�G�ZAw2�f�-U>�B�{���!è���i>���y�]M��=3+��kj�9���y(��q@�k�_8������S
���8N#෫#B&<���-@ڇ��8���bjZLX��#����Fo����� ��KN���%`�y�3��k�YN����c���r�����O$�����>@�����R�@�z9�yM90.G�����<1������'��I�(�����s\�{�s��'`<����I����I�������?���}
W�H�;��e8M���|�����ĩ�	���ӈT�������ӵ2���Qa�qP�;/�aJ��X/m/��mT�?X@�2wa�^כ�s��L��7�3Qpt+��j&|�j�GE
;D&����)��$�Z����8"���U;�*��0���Ol<�k(��)E�#�.`shi-��Pϖ 1L	F�nA�w+�JY7��p4���|"B�R{�j��S�g�����Rw۝È�a��5�P��6R*鏏$C�M�>���"�4y�8�����胸�f�N��5�������|i�o�Q��"��B��Pd-�<����Z(��%j/H�����h���^fn7j��&��3;�D��=a�]p<������?J�v(�UV�Ý�����=�[h��nI0��V��W;�>���u�@%��2��:ځ�bi�oR��됞�5v�4��w��(�	��4���OE/���U��"5�
�g��*@͵�󏫠�
Y�1��,&��O����
�5W.��h��x�G��4�u[�����ZrG Q�Eo筳H̀dӳD;f�Z��o�z�hTPcwϵoH��Ӆ��;��螙������zl��!\*��s�ᡗ�U�����2[ԔZ$X���A���&c sف���&����r��D��x��3��R>��{V]��`*`HJ/�G.^��M��\����?�dq�-gc��x�ᑽOl!Z���`��f��{���B�J�7����������k4fJ��w%/xn��l�t����1�rA��T�Ԟ��_��{S���y;��,:��(��2QO!��p�@9�s��c�#����*��."���� h�$�_ ����R�g�K]�r��3+�P�:���b��lN�T-���<����Q@@� ��v�k]BP%��FX�K��"�V��K�����lsg�k���_�'85�F:�]�@�d�2'�<�
�Y��Oo��xo:..�����!��|��"[�)��9�c�é�6��ߏ������ћ�F��)�^�qd9e�f����9R��0:@*�g_6��V��Lh��*T��K!��!��M��8��~?	�6�����I��D
t�wU�@��TP{Sb�'"��x��/�������Z��!�~g��s���dі���[��!cD  ���;�!�~D&9.�r����9w�S@m�-���[��Q��I��o����R�
9����?���:qΝ��(k���t�
Y���,��}��������h̖�W��3Y��#<&)yu&��B��I�R�oo��E�ZU�[�|O���O��U�QJ���ᨡ-�@����I�[H�_d��-����:h���-���&�������̸��{����ED3_��3L�"W�^j��|�.ǎa�M�b�* V~�1�����7�E=&� ]�џqplz��/�"�kl>��7�$!��>#�~�^>_���w<3"���{�f��)�:-l.7�g�Z�x
4�:
,ߑs,�t��\� R &Lto�]�jj��zY��p�ND���۲ht�ȚE�m4���ӨJ<�"pG��\