��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\���V�fnvx��ÍG_;�ȅe�~�>���9�>��Y;�0GT��}��E�I9�L���DZ�2ޙ_��
[՝X��^jE������V�����qL��ౠJf<���]��]Ƶc�yK��j%k�zZ����_�q$�@���↹c���g��cy)Zy?~�OB�ፀ��k�ӓF_x�Q����7j���DF�Fr�\�a�z���>��^��{_�?3xz-�j�d�ʸ�i�[���Z5sn7���Q���Z�Ej�qhT���zXf6�1���7�4��1��K.��ۓM��--���yp줕�i�G�օ{U�d�ܻ�i����B6.�	7ב��d��k��9�R��=W���GZ�J�e�*�:n=�kja)p���}��8����l*�[�,TY��s�vC�B� Of�o�3��o����kB%�Ihv^��$V7��]�����O��B2����!V@�#JV�ݎ^@M��	����}A/�k������]���Z0� Y���`$?��~�(Fod�%�eb�T5<%g=6q�j�<�|�Dp�6�\P��b�>�{���}�,�,Hn�
*1��KʴU!��8���CZ��i���V�\�����C��?��&��؃06.��
g`Ǒ���(-$�V��,�7�f�I�	�;}��5�s�z��b�z����$@
�$��#��xo׌2�8�-�)��j��7��K��,� Hx��Ji+�C+O��VG�:*�Q��;��:��'�C�*�\O�qǰ���vڽk�������]kU:��CO1S_�g�~[^�X�d�6ͪ\Y)�l�xڝ�7M<0����0��R� 1��Pi
t,@FX�-�[y��=�����=y��kU?��#A�b�tR�J�ԭ�"�$J�����1�=��j-�<�S�J����bb@]k(��+�h�O�°L*��������g��@��� �f�'���z�ē�:�Mav�_𖆜F��`;�.$�#3���W�~2|,`�$�+�-�T��62Ht�������C�X\�xO���^v���3ץ=4�����BW��Z����bh�����|z\2Ts�J�F���V����߳���V���QY�-�h�T�&_��C\��t?�|���x�#I٭��tE�h�YJ��5��#�J\`X%|�� ۺ�ݮ�ڤ*�P��G(,4�x���>��.�7 ��/�� I�A�Mj�F��r���h���b1sʿ�qDڷC�R��W��~��%;�7=�]��7qx)�6��ǾU�RI�AP�����׺$`#aH�ԦΡ��y��.����.�C� �_������
x�l�y�:���쎄\wM"!��{f�.���kp�����%f���/F`�9k��G1���Pr���=�@5�v�bI�q2�=���_�E�?��)�h�e�0�u��Li�e�lE-��7Qu.���[�o�w��@%�:1�N(�����+�D"���g/��tM{	��'ⶄ��S��Sw8�{���c��߶u�4:uǓ�Tl|ڹۯ�"�ϸhc+ɪ�p�;���?lia�5*��4u��*z�_��a��|���w��:��獗��8ed�Wln2���}��Xa�|��S}��;d����)��Ė��5��8 ��/��Dn�ԨCp5IV���@��].��t�8	�\�$���o��g�	߉�%N�<�.�!r'�'�8�P.�h��q g(�}2B�Y���@����Ev}��Y��<�	���3��CŜq�o�[E�z�'r�|�����M=�:�7 =����K7"���2��ޝ��=�瘰gn>z�"�{@��P%�q�G;t�ݳ��s�� c�&�Ãڗ�@	���9�N�|���4$�<�g��݃����OY���B�Zd��@��GN�P�Q��~��q�XB#{�G�f�}��*��`�$ԟ��N�띇g�/ª+�]�a�x��l��!>D�	f�*ev� (@� �4Zs����Z���Mʯ���
�H5t<h�>F�1�d6���sm�WDf�p�.���egjʈ�r�u�FT��)�r�T�����eJ!�˙DI�D/��{�*�!��_!��6`I��c�7���[!���y�sz;�pM��V�nA��R����&���J�"����is��8ge�*D
�d�CY{Y��t<�ʩP+W]u��"���E�g�B���#Ū���ܱ8���]J�E������ #�%kX��<�,�4j�e5� #������_0��<w"�_P���z�E��Ŋ<)
�_I�^�
]���ƿ�:��U �3\�ݧ� f�B׶[�ϵD1B���ev���xT�A�o�7n>��%�gy~_���SXv�HH;�.�vQ��ŦН�$$��I�vo����!�H&�k�H��^0���Ju{�NU�~����+�`��Z������Ч{h`]/�{N=BTzEm�v]�ܴh ޽��#�;l6��T#2���f�ME(m�,B��#љ�c�G���z&BbI�fu�7�w'�/����E���fO���z�"�P��*���<�2���P���T�PC뚲�����ˌ�L��E!�L�G�OO�@'>η;�@UV�Y';�~+�y�ɛ�u��L������+�i��'�!�@a�pŠ�
ihPp�&�|s�q�� ~����'��Xsa[&㹂X�#�\�mKŒ�spL�2��?տ���(��N\~�*���%n�+4h@����6�~��%�w&�f���!�ٍØ�a��'���f�|H�іq�^�g��,աr����U�G��ҽ;��_@Sݎ��;�R��\ �-dW9���G bŕ�q��#��,uy��-���x%��`��B$n��6��y�NwY=
u�;� 5�#T,�� ��Ebh�{����Jm�)|V����u��X���އ˶�J���B�K����9�,���n�"��T�B��뭏���ʶ��8�O�όm�Y��_Z�`yA�������'�	��۟�)�';����,2�É#jg��Lr�V�8�:xH�����Z%���ER�MėW��HR��*�@���� v�[J*1=�h���	ob`�J��T4�ʊ������ ������=fƧ=@��.�b3�<��1r�
��*j55Il��)��_Vk�#�}�-����"Mns���hR�a࢝�/W���}C���Vv�f�k>ܸC'�(�U�%ڎ�8�{#����UN1�ͱ�|x�1�Zω�=�(���\�l�P&䦛����-K[P� r(�.:<&�&�]��ۥ����n���q��3KXO�azQ,=�2��.�r18��!������K̑Y��1v�ٛn_5{N*K�}+���H�4�d�_4mnM?��P���1��WB�e�c=�j�
�Z$��z�.���/vPQek�Zon}�rv-��E��@GO��u�!CǤv����,���s�m<(b٠(U���\j8O����^:y�"se�+��&/�Q�T�T�v���Þ���⊙<��3�'x���G��ӾU�l��xu��T�5�@��_��(��UbqG��(�d9/�ԋ�M��u?���r���;栐R�O6�pd����x�|*��(�2O��-�n��I���X�lT^t4a�|j�]�avw7��.�U��)�`��B&u:-+�R�<�ϯ�%}KPP���cUҤ��T��%xt��7�� ���(X����[z~=+���:w������o���Um�ޔV�x���P)����L�!�!���ު��4�»#N��܉|�t���F�/��l�x�,�=\�?/�-Iit��o�(~�Kތ �5>��:qT6/�K?O��=ؽ�B��IL�&g�3J���3n-�͚����Ļ�����8R���^�`��wouFIĹ���v�����ZG�/_�n5h�7�I_�E�!-��κ��6;���ߴ=t)�hNK7�4�_UW�������1 b�Ę�v'ؚr�O �|-T���
�K�$$��͑X�ʙ4l�(���^|�� =�u(ŏY���:��ic�aC��~��E������WZ�r�F)�F��R^C�M���%������R$[�|�ƃ�r����j��a������E�r�;�2 8���^�����^���\��<ϊ�S̊�OR݆�ʦ��n�8�{J�I�+��7.��޶C�FĊ�o�0��[�_Vsj���- ;LLΧȯ�y��p���F/����j[Qo�A3�Xr.�=�3os���$����.����m�_�̟�â{��� �ݛ��qYC�0���8~c��n�]"�7��-�������O�߉���/�Ć"����l����H}�-�bS>1Բ?}�|������:��H�o�6Z�ΈN���-JF�k��=�T��k�0N�63�&��ɴB��[�	���:\}��K�:ɧyݯ��q,]EL�íB'�� TAx�B�FK���v,����@|A���J�'p_�����1w����0�'..�Ʋw&N�����L�m��f�Lˬ۽�������E}��P��Êsu".Q��.HN������4�2���*E�Y]_.�R���2��d���`0��Y8%N�N�8*.���8��pea�Z�W�a,	���cN�n�����X�!s@��v�c�i=�Ʀș q��Dt�%���ϭ&��� e�����몧�;/6�$7l^O��(La�'��$��٤*;௶^�rĂh���Ts�?�p�ʮZ��{-���.<G��'a������^�7�����1g�ͺ���2ӝ�d�'��}��Ǖ��[�-��`mE{�8��f��(���Ӫ�P@��E��}ɿ�	~�Q��;�Oxp��%L���_��'N�A��&V�~��
s���|�ȱ}��S��m�Z��ےL��}�1'wF�B�K'2n��
pM��T�%�:^x�\qV���I`:L���T��Ք��R���z����O!����C*�52���TN�Ε��I�{��_QC�촺1tZ�9�p��Y�K��ɪ�h��J�A�s?۽t��*���6�dgFkd��t�7O3����LP�jj0�L�؂$�B�R_yȼ��nu�^Oqr���=�ʭ�:A_��/a]$h_�-&@)�4���-���gv�S�Q������&Ƿn.��l�b��5���,�ca�d5js7k�$]�\62�a��[�J}��y��E�!�y����bS���}�]�x�r�-�w��{N���|��m����] 9�����f�AiU��ͪ�8,r������5�D4Hut)3:&�WY��ۘ�^�Q�>	Q6�t��q�����gq�S��2�~��,����dB�٩/;Iux3�k���_�O�^�a\+o�B,���VOM��J*�����&��#�p|��f��²�W1P龕���K���������C)��:| �l��&(�|��弾�,LZ�C�3�F�x֛�-�#ť�z�7?:4�����S��5qh�������Z�T��!�ǬBQGm�7*�>�-xSV����C�?�i�5M�F�g���N���V�}<֕
	��io�jq͍rU������c��!~�{̣��y>+���a>��ʮ[�&��>�*�)�'�G°{.��ZV{;5�<܄g=��;�G�w28�yOj�ꑾ�ٵQ�n�`==���#p��郞b�r?�7Iǻ��%<?���y�3N�ȴZ��B��5�`�
5�g���VQ�9�:����!ɣ\M�7�_�q���w������Ax?lP�3�MD2\J���7���~���`��ChNܸz�m��ͣ�߰19��S�eV�]ۅq}.]TT�j��/g��?wq�7<K�#6���k�<�]b�@���IDB�&�Wd��D��6�G���{�f�J�[�p�d�#��K�&h0�ޭ��܍�O�����|orM�B���t�w H��®?3��ƨq%��u�\�=�"�.E��6\�S�:~CC�\ �P6ee�m����_��G<!�H^iL��Q?�vիu+��p�C�
�wg\�h�����J��CB�oI���)
���;���AE�(y񬇬;�
�U<y�ٽi��31 ��Rq/�I�=~O�'�pW�ib`J��k��>k,Ey�hR �ϲ�O��ZH�^���I�,��wdp�9�-= ���*��-KX�T��7Dk���� "7�[k���MՈl�=x��L�ە���2"wi��r=E ����p/��_X��>���F	��&�Wa�j�w��yŰIRWD;���`��SaC�Q	R�+��q�Ex��%?�Cm����HEP|N����qK〻ޜ-^k��h�5ü���͹�KnD�#:���K�TqAi�W�&FH�>,�?8	���!$c�1QAIu$u~�3��-+��źr��X!�� �u����PW�I��I��٨=�c����e�o\�Rv^�������_8�2L����Lo�
W?�iY��I�8y�@0ՙNv�d��!���a��Џ�}z�Gƚ�hl^Zθ��E���Un�K�1�Н|�A3H�M��?3Jo����uɐ'�c�)��=�k��U���;%D��Y��{#a\�"e�ѹ���|+1uI��=�?� �W#Xa,yow!�(�\�@��k�\����D��iڪ��X\�z"�������n�J��*���Y�ۭ�)��e�rY��:	���A4	K�� N�6��o�`L�r��:�Fݯ�U~̌sZi;c��]M�q'	dY�jw&`�6y�Di��'Mf�Y"R��w�+��vk�Q�T �Hk�貴=��h��C�t�e�s����Ψ�[P������,�a}:�g�|�/s;-#H�#e�>���I��	)4�3��t
?�V�8Ж�&��]���q�mk��6S���CQ��2��u�y��j�������?>|���%~K��\�Oƾ�}�I��4�ڌעeQ.թ���m�Z��l̋gTu�%�)��75<Ug�\�ֽS��I/^;cq�x���.N6<��L,m��;!lC�!d��1!?qH�=����{�P��ʲ V4V]�߿9�т�]~_��S>�.>%!�0��ߒIU�.*��[6���$[���3jy�q�;�CK�/��Cz�C�f��K��kO�j��PK-���Y���R��� ~�9��1�k�I�=�s�D����6�½�����Ke�2�,�i��ȰUc_�{XW~|,�w%��M�f���Mx���3lo�OO�θ ��m_P@�sM��v_��ʍ�DX�%�s�ho�@Q��?�`�J�h}��P'�U�#���@x���O#��v�����?�>p�[�[�V����G��Y�U�Ru'A2�ҌX4���v��
����J�����gJB_$ uͲE�%�[��4k����q#�"u��ْ��	�7O}ZÒ��9�c��9�%˜�g��H���|��а0�B� =L�Vqۉ�������]��.5vn��f	�HT�Iˋ��f7�NT�6�ߟ��n.����
L`��vHǸ��B�+�Z3���K��݅� _l�ՠ��O����v��>bPr����4����T��=�?�<Z�6�H����~x��8tHf��*-_�(�G�+pC.Jb'1*���-�����3�&-^=.x�b$�_��q�x��c�����^���[��:�6���PN�D�	�d��
]�#|�C�F#��и��5�{� �T*R���$�kcsC��9C��F����Atʜ��!=��ZK���3����?`i�M���f��?�#�J��5��@G�=O��i�lh����-f9�D�s[z��]�4�s�e���ky'��_(����I���V�:)~��-��Nr��N(�:��/�3�KL��6gb�_��/s�Ԥ�X���0/0��J�,e7� \�G�-0�E��|�%po��b���ꕿK%�.j���U�x�rMZ�ļ��<�q:iW{�fO����:�欅%�&���͔��~K�rW�~#!�E�6�@�����\��)qi1+�.`w��śwg�c�_��3~��������åh8E�Ju��	�gSBb|�bH��U_�يʭ�@�2s֪�?' l�����Z)�@��FM2�����"�f���3�d���	GZ���7Ǟ��S� IR���v���(���9��Q*���G�1�)��.XL|t�A�+��33��h���PuM���
Ԫ��0��C�����&1d�(���_v#PM�ܺK��)5m��dE?�SXx�N�3�L�Pb���[�P�xc:��=?�+t
!P��pZ��F�}sb|]AA�5�*�qV�1�~\[���?��͡=�/
�����Y1��:j#K �E\E�n�(w���ȤW���n��0�t�Q�����?��BT"��
x���a26��i#j�'���E'.����	�M��t��	|f�sí�-;���m
퉶�tƚ ��<I0����*�0.�Կ�8���A~����"� ��w��=���w�X�7`&2>�-u�*/��.�C��}��H�HZ�H�4Y�J���Lu�	Wn̶�|iT����C77�x5��%\߷�� �(��.�ʇ�U&wM}�n֚��䍮v<���&��Q0h����N��<��?�&�}6}~�qDe1)�z�)x�ƒ/�c<�iަT'����c��[�$�i|�"G�䯄�h�{�H��ڇ�������0$�����Y�˛;��ccoc��	�3W~��3��[�/�/v)��t�]g�	?C�&2�騧ȝ���zjupؕf���T�c�h)�H�o@�S0:jB^��q����M�R�YF�ܼ�E�