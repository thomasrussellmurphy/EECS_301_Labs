��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\���V�fnvx��ÍG_;�ȅe�~�>���9�>��Y;�0G�Q�Z}.ed�n�n�HP$Y���r:�ɡȺ�i�:%'��������㤉��-"�{S%Ů�$B�Öb��i?�����U4g	+©��v�&�������Ԛ�1��o�vA]����5��6��Xx��=f�lbF��>ɜ-��B,��?�T��F��%AGM������y�H#�T5j���2H��z�8�9j4@�\��B�x�`�Z�j��_!N.;C��lP!��-�Hx\�k��w���y[��My WF�Ӄ�ē�Bsg��ﳈl6�NB��LI@7�����
������
Ϧ_ˬ��=�g�E!GMC�`�b�(��$��Z��6���Ӳ�ҹ�*��
'�
xq�*<Wݟ�D�������.��N�G�i }��KV;7F��Fi���I&a���1����<�2��E���'Y�|%a^��� ��^�}�.�+����+U�_�wE�j��Q�'�A�⋭ڭ�GeՊqs)n�j�j��٬����� �!d�Dm��������Hv5�#EFN�exDߥs&+5��o��Q��,���3v9 �ˋ(�9k���q�*?�7S�LV�ӷ�'z�����X�qa�8#����۰c<�g��ڢ��v������>���ġ�%��6���'�0z�A�+����������3=?2-���ȝ�g��_qߣRH���4$�1��+T�sw�&&��KCSH�^�����-/��� �HCK���;����+`V��de}ߐ�u+��砂_hb+
�)�lU{�!q�y;-�,����}6�~to�Kp��Flb\PM7��G�Z6M�M�C�i=k�V���`n�=���{�e��r�e��SF�(R�׏���)�pg�UKȧ�7�-���@�C;k���t07<����OV�9�l#�fZ�լ(�-�8��K29�腵�$�� nQ$h��'�7E`F��d��Ѕ*��$3��\�5�J����*f"D�eff��ep̨� �!���fF�
�[��K���>hW��&�ܔ�K`�C�Ô�D�7j
���e<}�p�Y�U5��/��B��P�+�yV&n���.��&ԝ��=L��)�)d�ѷ@�r���(��h��=F��9�l�$C߹Ka8�ϋ�%w����D��I�-em��Y#���� �H�C�+1���i'��B��x�_�L��5�CpViy��9 H���G��1E��������F#ɤ�y^vm�A@;	 �շ�~��\t�����@jE�M����"��!SA��%9P�hHo��Ų"�ёW:`�K�'6Q�V歈,nT�B�jC��ĥ%���Ѡϒ��!p�Lܟ]ڋ�&m�Liڙ�^F����gn�4_^�,�
�L����7�vЦ�;����~�nAo�t��L�;ǎR�T�׀�#g�a�����i�~�|�����8�G>N�	���4�a�1\y,��UEX6H"���,pX�<�"M!�y���S�{n �Jk[�in�}�c@��;H��ֳ~}d��o��k�n���������B�0�c�{�,c��0q9S���Љ���HA����6%gB�Z�d�����Z4@��=��sD�4�}z��WD��=�^�X�GT��i��ѱ�@�mcb�":�)i�8ュ �-��z}H��aS\�nNΘ~�-�,#�~ðeL�yя9���;��Kq-���$B���g����ez��U�+��Pio�QM��`��#w�8=p��D�w��R4M��1E� �����BA�<�H�X��.�g�<w��
�[T�M��f�"���c#6��XN�>.5l^\2廵�S�=�1a�3vxvJP �5�T%�T�1����b$@��D#���R��!V�'��=5R2�E\��- �t$�SA��Ș�'	��f���,�C�Y��A��Mm�2�{��2n��kq�XϦ�����b���>}`�<��!�D�B&;�,uu�刃>q�8�yYk�f�h?�����ż��Hv���@��1ԗ�ȱ��i��³�p d�r��tʑ�~�?7$���s^�8.�%�>��p���#݋��Aoy#Q;៊��a{���e*<�ņ��E
g�2U�SZ�K�c]P�.;��
ɤp��S
t�M�?��Gx�)�iz=b��V��~W-y�|��A`a�	wH!xR���� c�Sf��ڲ��lkm-��zB_W�6�#;8�ggb��'�c�Ĉ�}�;{|�Ѳ�r�M��l6���U�,��7,��|�d#����-f[y.�,l����b�D��[��p���5ۨ��$�0�^x�n����l�veE���c��|����f-�YХ_+�Tt=���P'~c�5�a
=�d8���"Y䲚`�>ǕZ�ӔT|H�7�Hh���L+N�*$�~,G�kG���U�%�7�
\[Cm�֙"ϭ�ʥ|�wt����e���a|�����J�gujx�)���D| \9�E����$�%m%�%���9���w"����
]�X��^G�J�HY���m�41{*�?��ٳ_��|�7�Xk�l�Jt�.M��):��C�?<;���Uxs�H�z�#E�_��9�ԕ"�/ퟯjGH�a�d��j�I�O�kE���.�\S�d7��\]��-V�d�n���9�����`�\�t�fQ��mQb��.�Rqv�1%I�9�?P�[>/��N�iR��$�)_���b�2ƥ`�Ӈr�	��E��Y_W`���ܞ�`p�P����F��OUci���+.n�=�d�h���䨍�:�8��z��?��ѶH@֍^���CGK�.g� E�AB�doTN�>+���~}���
`����h5&�W��C{�Э}�����z ��e%�)�ٰ�`tҶ=(��r-���0���	#�ԃ?��>�446:�O��khrݥa��&l�6�@�uDl?�HZ�Z��9D��o���G���G�vV�t�*\�G�â��G��I�N�^���r3�^9�J�I/,���#��{�(�(��}�A�}�iXMPP���|�x�@rp1Y���4�j����L�:F���QA�7��Y���|�2ڢ ����S��Zr!5���^T�2R�p���d��9	�#��d�O�]��+]��I�	��U<z����R�`k#�~B�Z�C�h���Q�+��ǇT�F���(�5*���W)��\F����[��7<캣<<�	��KV���^O�U{����C�E����F����'o|�G�ƹ$TU�7�L����1��`;6]D� q1��|�i���|A���ݸ�&b�SJ�]���C|�FME���(T�|$�������{5%�ʇ�T�A�n|����{א�2t�����7x� w�8֫J�tB��衙�;`�V��
=J��F浟ip�7�22uǦ4L%��4`�?�`��<��d�5�Ψ��꺆��63~�-%���C��1Q��� 
�	���"-� �r/o�P'&�S��_�E�c�Pjut���?�N��%��2���g�K.#��X�Q����b�x	��;�����F����8��5��Y0We���O�;21�tR.Ñ3�B��]w���e��?�� �'h�7�0T�� ��yU���W�<{��i�����(���"�E;��-�����	kd6�"^ {πfk�f�HAM�^D4g���Da˙���\K�l~����p���-���,ƹ���Rd���Ɉ��TN�W/^�A�#Ծ_,�j�D�d<ƴrq�I�)�]>�|pC�7z_˼-yl�����!ݵW����=��y��[$\k;4�	΍�$3W�o��Co1�Z�&�35���U�w������c�!��F��!������?~��7+�H��Rs.��0�w����e�֐�]O3�l���y��ͺ���ެ�� ����M¤��*AX0j��K+�{� �a��|3DIA����豭�GDr�߶��mv�#j�\��p�G/jF\L�T���No̖�*�x�x���C�͎h�i{��FڵZ����%��xV���q�G��|3l��>&r�3���p�#7�D�{^�b*$r� 7A���SA\���F�Jp_XwK��:�_TP���l}�/W�dm�}���ex���=հ�I	�q��H��F��^;��������m��Ayв��DQ���96i�7�17��ڄ���Ì�]C���:7r�+���)��z$����� ����K����UPa��?�]
�W�z
`&@������/0�0}R�Fz݊��< bq�K�.������!u���<骇��V+�#.Z�gI�o0߳��]�l�;0��8;<�@��J�d���ê��9�q-��
4��SŹd10�5��: ���X}���숫�3�Ui�jUY�<P�����(�~�JM���b.���&��m�,�����7O�Ӿ{ri-5tj1�w`�F���Y�)���,�R���N�F��,z��	SDNY��wɉ��t�`E�I�m�
��k�W���fCy��A֙��A��l��G���zD�D���i]b�0�[yF/��1*I8��#,k��������*%�x�˖�]w-�A���ƀ�mݛf ^h�.��pw����'�1�V%��e���O�y�>�?���~��];�H5�l{[�DI`�S��7ELj�4�.Y��yR��:��X!�Q1���W��@́�����A��U��/.+kP�O��p�&v����c���[��4^��������O��^�ROT�3�^+����0z[rΨ�����3�a_�jbi��5��%ϴl�o��A�MEQ*"3�:�w�5{���!Ѻ��68|�=s�'�E��{,��k�=R�+����	nN�]|�ܬǇCl�P��s��/�؊�k��� �w�VW���􁓊�=��al���2��SԹ�NkCo��IP����<���@hn) {�'i�c>"�2��F��bmaR�c}�KX"W�c��P��M�)�!�'��'��:n̝6c�L�rj��X�3懎�����������+�<FC�e�c$�8)E_S�`���%���-������W�7�*�QL%���jS# %Jv��v��\��[D`�tY��(6����*�E��kze+̼�%��Q����>gB�=t�n�-�gt��������C旫��y�_��P8���6��$&E��[���x��'
uRU�ڕ�I��m�����-���I���j�)�M{d@3�؂�g:�[Z�$F֐�3ٰ� $j�Wʷ.�'D��ʨ��j�f��	�t(V[t���p�dWL=O��3�L܅'zT��w��N�"��o��ג.jr��sŖ��I=?Ս��[��7���! V3��HA���C�C��G�׷{2��@���6����K>�>+��x���|!�o�"�~W������*�<�q�4��
�,�V�P�J�RT����P��)'V�r'�#�!wX~�7^R�9�m�`|�8emm�C+f�Ʊ�S��#�X˓ӄ}�E<ӭޓ��޵��v�)8d!�t�=x����ֽ�ԅ��R¿��@K���l�'l����Z�����'�����;}�~�A1=��i�;�[B�g�.�QB�{���d�*�2O�\�o���@U�'eٌ�-��Xc!��z��Y��z1��xM��aî�ǐE����jU����@R?�,S�P���0r��Kp��^��:Gc>�W�p�rಹ	ʛE���<(��t��� -����⛓g��+	�\��wlb��Z�����qF~S�̣!�1�s����D@���3�@z�k+*x���+Lst���i��9 �~ao��E~�������ˉ��&
(&����Y7H��`bh&.<��E'"���M��k��
m\�X��z���Uv��;/4(6o�hE��Ķ�exy�=N���{Fcݚ7����P�Дľ%���kL���<�i���8�v������.�+w��xr�'?���~m3ʅ%�r�緢/��"t
h�w�Ճ�t�V�'
;���YR��̤���` lE���p�}�������?��F���0fw�C�D�,2���C���yڠ�p��m�Zdh�C�����Lҫ"c�&׬�ǭ�܅�b�X$�?�E�0S/T(`���*(�Z(�J����3xD�"+�K����J�A��Dn���]��{x%��5mm��X�-��aQ;�k@�WƷ�,��,��J���i��.om�m� _(ѦV���u?�O9P�'1�|YEM��b�|�A�N���G��U��0�� ��Sr�^3G�Dr�P�`A��0K���W�`�������K�"WG���J��I��-�؋bK��������'e��yw�A0O��+0J�;Q�Ǽ$>��oa��s���q��i�� ��G���Q�yWQ�R��jg��I���'%���^rB�}���JD������3���=�
�_�u�D�B@_���Xe	�S�{���W�x8.�B��|�+s]�"�Y^�q���y<���s�8G���jt�;����"��y��N6��+⛣�K~.����t�|WWJ�1�1S(�c��4�c�
i/�������t'h�z�ADɱ���}tj����3��V�|N��IUp*�I�l�����0{a�&U��G] |����z1�8�{�Phw��eI�"��4��ղ%.Lȋ��6K��Ĳ���o4�a�[�\j�?%��0��Z�����F�gNE��,�G�Q�b'�[�ֹu�<Z�'D��y��c�Ou���0�����ͪ]�gr�%|�
�$�3��2d�d��	W%H�R�k �LL:p F�4�O!�+|bz�t�(J��N]ʣV^:NB/q���$��t@��2s�`G�@�n���������Ә2���Z��IzP^?���B�g���L��堨�:�Rni��*��s�`�"��qk�M؜gU�+-���Xi�\C����^�X&����֋�w�}�k�$��z%�2l*�M�+@l����\�Ke� �A��~�� ��6tk�p���9�+�[p(�7�U��ۆ2\�WKA�>�x�THY�u&�����\<��!"����s���@W��K;DU'�c�� D&���]C�8hЭ[���i=���uŉ���O�PcV6^��o�$�S�r)~z/}u_�wEd���$�w�r���m�C�,
2H�ك���������6�Vi���q�@;>����'�e��V2����"�ۻ{5fRs�j�Q����\�2Az����ܣIR���W��f���p�X��Sng� *3G�։����B��G�=��\'1L�a���7(^��8'��|�Q��com��nЀ���.X�o���*aYDq
Σ+t��؂�P]��=��mn��$b���5|��|��cnHz�� W)llM�d����E����b�1�JV?q�@��<=n;kUU�ⲺT>���8����
L�{dL�deU�B���*�fi���El���!n[�OV���"��e�~�;��ȆbH�\�-ȱ<�U�!o7��f[�M��a%��e04=\�u�5~�j��"a��޼�W0ཇ� �1��Eq�A9ꘁ���I,��M�D�8����i�<|<y����?�Co���0g��&k�y��2L<�!�>~(����wؑ��b1����]�O��D9�iU��P�!ɩ����U��w
ލl��"��E�ٖ����D7�L|-�Š�ǔ�_��2AS�d��چu��Nћg��M�P��f����O0���+�?��v��^Gժ�x>:?T����e��Z�o����&���[UTl�u��v��}��}�9B\��ڗ�~$^\a�w@�D[E *���O��԰��T�lǪ<�B$����X*@�C&T-��e	����=����kN#��ݪ�����3�\~�2���2��c[z�W��=�	r�L� ��r7�"s���^���tj(̪������&�N7�;�^b��ī�`���������է�.<A��N���/�����K�5��(a���������/��D�/=9t)w�$�{UJ!:.���rg����佣,��d{�UKN�?�� �Y|�!Plu�i��n!A�)j��ds���Il�5~��U @��v�rH�`F��;��i|�8�<Z��?��}Ɍg��?}�O��23���U�/ \yF��5��+Bo:(�z��!Xw����&��q�V?�[o<m������	���oN�1����B�a_E�6ο/݀`�±E�c��˾JE���ҭ�Izu��TdAxo������B?�Ĝ}�֑�K8s�锞f�V�^�/�����#5~�Mo�`]��]@���%��u��U?�Ħ�q������ݤy�q==������i�����B��M�e.�q�*�*�u���EP�2-.c���u9�J����D�8���#��H��,��+� �{���y.b���^��i�1�[���X���s1dK�z�F+���j� o�ڝ��v)��ݯ6D޻�9H�a��.
*v��6Z/�4��ϭ6>qo��*;��Q@�*�_�� JWيC�-Z���O��Ǉ�R��{��U���n�&] �M�	y�g�:b����#�*�]�|͑r)B�����Z�}5��5���04\>��r�����`��fmmE�@^'�O����̊�E�+�D,�C��V�(9�C)˩iΎ�~���&�v�l�Ÿ����zgM�J�R�#��,�� ��7�
�22@o��*�2W�4�݂w��~ ϨZ\�[��?J�A�>%���Ű���z�)E�3u1��#+3��\��_x��sZ���.���M�����7���4T����L�g�v�88��jb�l���DO�lj�����;��n*�#��hI���� ��,D��H'Xk�P�sB3��j�*�#�,���%v���L?��3��Ik����r _Vf4ؒz��3l��.���׏�+�H��̮�38h��������N%�	ɩ^P��DL���H穔!G{]�mH��NEf����1xY!���5iƏ��F=�>؟�)��j�ϻ[|�2�sB	Y��(1�O���܄��v)�m	��n�A����	�p
Ǯ� ��KowH_�?0�/Ɠ�=a�Ԏ�PH����G�_�ng��M�c�14r���2�UN	*n믰+֨�Cg��k��d;�u�<LVe���#��D=]Ɂ[�����Z+Ez�Kw�ϓ�Q!�op�������r�>�]�3f�0��v<�o����JY����M�0a�>0�m�k1�k�_#���$�Y��f��%��e+%`Crn�O
0G�n�ҭ��9]� M�a�FR�?�6��$���q����˖�ξ~�ū�BSN�*>v�q�[P|8�*w��MTZ�Iz���s�j�*M�]�ٮlq�-�r��j�K� ����gѮ	�zcU~Vpԥ�s�;�<6�2�ü� M:F���o} �Z������zw�gכc�|욹�r:����G�uP��yh츽��I91���T��'xH']9Jߊ��v��%�?�t�8����2�)h\9,58�ljh�ɯȏ��ͅb��U'�s�$P���lt/���4V&�֑ٷ|����u�4�� ��N<����˷��F���sZ������g63:���:-m���"�'ƸR�� ��	�Mfd����L$���1@`�O���[�ޅm�gG�g���	��8���4|l��M��xz��A�W�j�N����HB1��2�#���;���s�a��?��X�9����#~ sn79�9R�z������}2:I:iq���)�{�s��l���S1��hN!��zL�=���*!;v@����l/$7��ֆ�Y�0Y�"��@�Zyz���f����Ҟ�.�:�{��gϵ��N�\$�[>e�2�Xub��xe �g3��/fe����h&F�����I�Sv+:��
�Yڈ�@�Fϱ�V��m$��c���z�-�+��[��/�2���n�u�l���imk	��x>�.�#�ڦ[5�_�ܴIo,�PS��Xm��a�im`f��?E� Lv`�K���9������p:yQ��{�;z�_e���r��2�I�)�?�o=�+_{����J�+ҥQ��&��?�����W��@!�F���^�k�H+˕��$h��s���_Þ遍�F3�%"�is���&Z��,)on��U/����IJ��'k�K�RX�j!B�Q����@����l�t,8���2i���R�����"^�֑6����)��DL���~㗪ɭ�[�4�=P�x��O;3�<+�`��}��-�b���&D�w7��Z�� m<�����Z�p�l��C�
\��Wi��6�����v�IU&ٮ�(20pv��CQ�.��u�"��ȷy<�����f�h��W���a�17�I$��\e��x��iӽ��Y�]�jpt�O� =Xd8�F���6�� ��9�%�`�ceM�)8E�<��u�2]�Xڠ��\�k�~J4E݈ۢI`k9Lէ��dD�&�.dc!�F�~ó�S�E�KzE��fN�Kؿ�x��_P>fkY�~8^���s"}��
��u�V
D�6��؀��B)Y�$�ָ�JǣSJN�\ ����MH[�u��3����7�mʻ��J�/��Ё϶:(�鑌&3��m�5,\F3�����z4x�I��WK���0Zq刅)4��0����b��{�i���}Nu>��E��bt�ǟDG���~	Z����[>U����{�Z���q��-п����W�'�:�?�%H���UW��,�6�����.h�� v�@�dgʈ$h�Ѕ{!�@x��������\�~�����c%tH���K��vL7:(H���U7s?����z=��`$�a-�9��^9��$/��qh�!җPU��4J�bϘbW��z {������h��̑@���qP�L6�˩��Gf�C����0��8`�n��y7�)��+�&dƊ4��V>���ao�9���쏈F��s=4]�XZ�{���O��j�bFF�WJ�o<5�����5�<u)�B�'M��Ś�Vх]�jL����?�+�W�]2IY3
�� ��l��3a��U�rA[u"��-X�a�Q�"��)K��t`�.�!�{�Xi6_��C�ѱ�-��o���{~-{c�xQ�R� ��4m�}�W|�f�M�hj��0��ϰ�>�5��ݘ\6�����>��bl
����Y�c�X������x�Z-"xg�w�/M������GlJd��k��#\F��9�!b�xKs�y��������<c���xy�J��:�м�ڡ�4����#rƐ�!�^ʧ�r����/�Ud�U�l����d?"�cTRG�*�j:z�5~�����Ma[�\Q�O�)v��'L�;c���ւ��˔�{��~f�������|.0��/1VH*T�V�8�g]���p��Ze�MY�8���Oɩf��`�Hɱ(�)?uEy�-^ȗ�$��LL˵h��T(-�+��2�n[ >;�+�/G��=B*�U�N�zKx�LK=#��K�UK�kpM��M�N"���'6B?���H?x�4����,ȺN��� Ͳ���·�xsX<����i��ւ?���d���+�j_]�!���'?!��uz�]%��?��:$b5�������NM�z���5`��I��ƌ�_H��r=�-]�z�p���9��aN����%C�������$��"FVRX����F�[�J �0��� ��ʚ��ם�� N�LlKh�+�޿]��t��+"I��N��z���z_~*2*����5���svz�z�ut�9Q�h#^`d������ȉx�s mTA���d�SX�k��~!9Q��(O��K�4�Z o�-�<C}F��|�۔^�0�gwQ�?a��5���&q4MvqI$�\���f�Lبt[O��v��penX�̮�Ϊ��0�&�F���	by����\#���
��0�5�xX��Z1wd�n;k{�%�ϡ���<h�NN1:�jT�?f$� ��H��!$m���X�[��K�/i|}c�c$�%�\��G#�?d�K�1Ph'̂�6�����P���z+r��"�\�d0�k��׎�"p�J���i'=�.�<�<c{@
@�O+І��ޣV����װ�Z��\�L9�����q���([qEC�wĈ0v����^�buL*:K���&\U� փ5�c>�����-M��0z���� ��Ý�
ނDC;X�"�=��� ��U6��t����6F�~x@�z��AZ�������� �ڲ�l��Y�&�k]7���{w!i�@�+�����J���6]ni�V�9u��38��f������ZL��������O���]8�7��7x(\0�ͬ�v:Ǘ�Kc���W�lD���1������ӞV3�&���0�:���F����������,��>��%vܝ2���H͉�
�T�W�E�W�	���U�n���Ay�Nss�M��=������P�-�>8������ѷ�4k�j�d�e1C����yۀa`	f�ƃ�k<M�D����5��#�7���
��л7�7:W����˝k5�T��o�tD��]	p�]��U�L�����/Lp��*���>��~��X�g���E�d���r�����z($��$�˹̸̯)'�ӽ��*���1�n����zY�ϛaz30�Up�O��e�Yk��T&JϾ@.�y*/X�H�VZH���(�8���@B���+a�h��`P���E��.�(螋�(�#�pp��|is�n���(y�����L�q�>j;0�v+�-��� u�)�3|-���
�n{�s�l��S@"P����\Ū?q�հ�;�[`s��	���񥿬�a6�-�]����"g�>�b�֥�N��a�r�q�h|��64p���!|�6������~���v#�`�����i�^I��d�t�"��ʶ��C1p�v"��D�dN��  �.b*q&Rn;Rv���g���i�r�ś����}���@p)�sp=�y���\Q	���Hl\�&m�Z�u�|���;�y���̔��Y;�8d�{��:u���dz�ĒO��Z�'k��g U	_��)5�K�����A��g\�{�&�z���F����J�]>��p��ZL��^BlJ����~���7\�)����')��$�RO�`����=�U�w��]\�$$����zJ�
��r�ٙ[��֍;�$w֐S�${p���2�hXb��H
����R��)׀K(�;����ȄW�`��U�h"�tij�V6j����&�.r�q��n�JI '�X�N8���-5�Efv߫I��:��ʏ�Bm�rD��L#�33�]�a�N��J�v	'{D�u�{{u�-�+�ܠ�)޳�v[ �Z�{�b��E�����w�ڱt�����eJ�Kz�&�<0��Of ���6��'�y�}��#D�Ze���c��H�tB�ad}�?W��8�?�;��J��I!�����xvw�Qtdjl��v3 GPTʍ�ڙCeNw7vU'���,I���T ��cP����"�N~U�ˀ��i�@�ʮ2����+�Z ���K���W��@������,�[�w�5����ʲY������@*}�Q\
$1''M�M�~��1����o��"?%ڌ�[K�O��+D:9�I�b#<�ݣ������J7�:w�"iSj�R�-���=բ@<215|1��9��K�kf�'�Yb�m]/�s!߁ݗ�@ٶx��e$^9�_�������+0qٲ^�p�3�X�\��F��(y/����'�E�hl���7Ѕ������ZI�^7Ҭ�199ʼ+�z g��!�w����>s�⡎9�U�#��9kQ�1��3��-4�.`�95c+ߥ0ρ/ 6�{��6�	�!�ݺ�r)I�t��Y�OanņR���9��v��b����l�hL�G�B�*Ea�����j<<���ݭQrU(R�Z�z˅���~.�-���C�m-���n\2z%��շ�
Űh��o.]����Ox����ϏH``��񎑚[p�.T�8y����ùJPH�&�Ëc�=a�#9�Ζ�
F�!vo4�a0���U'�y�d�q�g�wC}�x�Xsky�@O��`�ٱ5�M"|�s�گ}�y>�yT�ڜ��I"��x4����_��MM��O���$��vd]��N�\�Iw�#@\�Wa迶S:���V^�Fx^���-��
�|q�$L/t�]
�=�[iitf��D���|ʝRZ�/ZTFp����/������#�����U���jb@<�T�ƌ�g�Vtz�&��ŧ�^�+�v<�bFs.$T�`��#K�8ҟ�+ ��>J�[������P�#h�#j���((`��������L�"���&�C'�և��2n�m���[�Ce��A	OK��y��'L��n��a8Qɀ��`J�ꅌ��~3��80�G��*o4i��D��j�����	]s��W듅|ǫ4g�/^��z��EY6F�zX�Dj�d�&:lدͶȎoxp��C�q�	���1EV��h�k������{�^�F.;]a���~T�ȑc�D���ʓ+9��z�m�'@�q{G����7mga���m��44ޑ�51��
MY�G����{�<�@���