��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��/��Q�w���a5P��B�~�/�'̙���S{���^�qѝz��'�hřD~dVr�F�!5�=��[�\�bYzy��d�(5���*������j M����J����Cw&�u����Dg��>_�,��o��3�9=]�sn��5���A<�-��Y�,���AU�G���̻N�	�Ϩ�g�ϵ�w�Ω�k���R�9HO�o�u�(v�W�T�yVL �q^�Q�0/�����)1�cڵ�E
�W�D�t/�Ș���~x��R�X7�]0|��?ͭ�m׭��e��%\rN���H�i��8A(_�P��0];�ű
�0y�����
�F�(�}�����6�o
\�Tf�,d���b�3��-���y�)%$#�mU�Z�%pS,̓<|�hֿQ��iҺԱZ�ͯ� ���DP��̺�
��I^x�t����ؿ�H�i��4��ڸJ[�����[�4!=!���O�F#z�S�։NJUm#�~R��'�Z����HA�.߯h���"<�I=�1���w]�G+s|���|�X�����*�� �R3+�(g�4��Ҧ��	-A3�.j�=(]ŞJd�p��%��{`0y甆dok�Pڤ��EUt�ȃ�NG����,��&dڎ��0���a�of�H��q1Ո�NG�?]G;>��|��*�͊�B���E1|��F|0G'�p���tk}iS����j�i���G�>G�I���� ���f8�����&�	�5Y��Yh������A� ��x��,'��� �r�І͐Ef�z�����Q�0�Weaν�����K�|����+�%��h�i�x-�2��r$0�G7�	x뒢ʀ����Y��x�\�|$#E��������ےĈ8�[��TEc�]2����-�܋_U(K������UB��"4�%��%� ��p:���yv@�����Γˈ�)��c�3s��t��b�K�σ(ׅ���ኳg��a�8&Q�����C��c�H	�Gi��:گ��%:�^�(b���E����\
��X��$~�߈Z�.#7��A�z3/#Su�{m�Pc50���H/�~�u�P��b�gKJ33�+AS���e T���~)������<� ��C�h�t���i��؞�����s|_m�p�6�o޾T��_�N�ls�0AHK�h��ۜ��1��!��yn�Pg�
�:���mD�Xz5���i��A_��Ǭ��⿯VZxzalO�"�S'�� ���@���$�7�
Ck7s��k�B�;Ɉ1k��<�Z��*�c�F*�ץ�m`�A����2�l�@��ɼ�a���E���G����jD=�Yo��=P�W)�@=�1t����VEET<�l� ���$
'ʚ�����b��r�i�)�k�I�zE�&e¹�x%=�)oĻ��3�	.�F��K)VB�e�1���3�!����}?mi� m�QP�EƷ�ᵾ,�D�)f����B�����uء.�����3-�UvLjr8lӤ�d�:���z��C�����kL�Z|?z�>��>ވ����U�Db?uuP)j�D����=v#`��O�3�۶?|g��4�"FVI����9WaF?��1H�
,_�p����5��NJ3/��(�h�Q���Y`rM���`��������@ۦ���ɬ��i���%̳T$<�A�E��囈=c��@&/��%��A�٣�˧�07�0v��D�G��kk���"�j�Y�3��|��sA�G�֫׮c�&�m���]��_�ߋ{Ky ~�9:4"�R��9�����t��B���2G�ddɑL<�Q�L�Լ�*�������K�4�VG�P��i�ЎM�DdI0�2i���Ʒ���a��{g������p/�A{M7�k¤�<�eͤ���V'� (u�d�7��i��Jg���WC�!�����N ��J.�N}c~�YU�1�m���,�[�Oa��j�E�N���
E1�u�'� �>r|h��$�Kd9�l=�a5z�1o��<�b��Ͽ�-�]g@sKC���,���l�+
#�S������K���3B��FB�;�\����d��5�  �J�o��}Ii���� �������̋{�M�2�&)�V�9M&d������8���9���$��Qa���]�^ 4����*9:G	@vxu޷%d��U���� �.�g�;K2C��s7�Z ��ƕ���D���NTb�o����ƕ���� �TL8h!e�QZb4��bdv?�Ȱ�an�3���'(����ա}����{���2W�uD��8K[�/ kV�Q`�?�݆|I��w����)U���&)�g��0{ݕ��^7{V�DM�%Yޑ�2G�v��	b��fg�� �l��H��`�� �����q������!GId�ٱU�^�����w��J���	0$ƚWp&*�����_�"���F���Y/G-�Y���i8c��U����;�oS*�f����X5	�������� �j|u�m�;�ޥ1qn����z-�)�k�X!�,2�����B}�����
i
�{zW�Ӆ�f9MI'G����E��� ���,xb�V?\�%ll�! O7(` �h$�jgjJ�
�V[Ή/�9�������4`��L������\�=�G�&=�����/�ݷ�\捖��¬�װ�&��2�,������
ͅ����@9;�;1$ufp \d�%�����I��H��S��[��(m��!ߖ ?BĹ����Ŝ�\��!�D�>���
7��Ğ�����,����*� j���$���0r��O2�z��#b&	��"��x7RZt�o,/o([Hk<�[��ю��*�����>u��[
���"�����$&<�6�5#{�XJ�����o4�MO����Q��Z;&J�ƞ��8'>C�5\8[U��}]̞��=S"���ۤ�1����'��3��۟����0X�l:@��<#�!�%�_�y�n�/�r���U���SJã;=�Pg�*em�E �^��~�-�B?�1�%�����tÉ�R�p�+_�7���0-�1gp��Qv3�����,��J �~i"[<.B�j��w3����-���[�]�љ�v˭�@_��&P�+`c�沑1'��D��P��CM�NI=;+*Y��cV���TVD��j� u�z�7�/���_Q-D&5�����K�V}퐊���o}RCc�vHr�DJ�cM��+��@��CU!Lm�Z���i6���@Ɯ�7���f����T����������FF��i+�*����*QL�����^�}Le����q���>���Q�L��Ö��dL�Og*�"��D~tp0�0���oT�I���oI�"au�sQ��b��(��]Uߜ���MhW*�rAI�$V./+�P�Ǆ��3o����k��\��o���5��Y0����C/s��SJ�N=g���D�[��/�e ��m�"T�nc�2�Q^<<]�Psa'P������,�h�R+�QK�zU��Ml�v��b� �g�!��W���? �5
9�{����y#+�HZ�K�ZvӝMP�V�u�oB�#
� ·6�d����n��ֿ}{��cD⁫�_����זg�� l� N�F�av�A�8�9���|V�Pt��T��OR�� ��.Q��3?HG1>��/A�-�����rXr,�@��{j�a�p�i�)Ic?�=s�1&b2�A�P�w{Ü"�')�ﰅgjM�Q��f(���[���J�YO�������#��3ia�5���m<Ϥ5��ϏC�h�ME�07rȆ�F��;�����L�]�T�x���X��O֑�
��j�&UR�R�7!F�0�z�V���b9wD�pz}>��Xp����R���w�����d��ʿ��.r�r>�������^�6�*#'5g��V����8����6��W������='7N5;´?$L�m4�:'�t7�nOfds�CuB��#�� ��*�Tݒ��?�k�gq��iD#&C�u�ɡ��^��nB��;�r���QiQ��Z��;.aD��F�4f��4���ޛ�A�!V���X e7`r���������%=�t�����2^���m��N���Q� ��.[-�|��Y0����h�꘢b9�u�ɼ�К����Ǔy�²!5v�G
�������>�i���?,C^�q���la�Ӷ6�	s ��y�����zӑME{�'���;��5uW�� �&�$7aW���В[�e�Y,jr��ķh��A�?=���څ����������	[˧u �	�L��s��]{��ό}1�#��o�<g��$�>�1_�'m��1gJ��\�%�5����.��[C�K2�Д}�����p�3o�ڠI�^~�/ϣ����v�U��Z~h��Ś��:��3��/=�{f���*F�/<�&dj4��Y�X��aF�*�����ոϯ��c�����^k��*��X;U+{�V' \*�`����n�K�fs�%w�!��K�����]�����o ֭z���pi��1�(Cj�+�n�ms@(��\(����R�̟���N���i���dT� �O���+*�L��h��p�c�Ω5�p�]�ͣ�^AG�̊81��,F�O^/2���K�l��K���L����B~ǔ S�ӌ��<^1��8��z�׏!%�e���V)��������Z��,(�<���q�D�>
T��-Ԍ�h�)upC����?)�����<��*nC�'?H{r`Lȫ�b�B�r��,j�l�M�C�����a~oF�f��}��}�����HL�1 5��1TP��L�|r�1Y�	��8y�^ڥo6�>`���K0:J����ĳ���C�2��4!kdѣ���ұ�41���%�n�e0ٶ�<�����|��>鶚ԇ^�{ّ\K ��'�cԆ����xT���@� >Z-��2i�@Z��9��n�G��3}�pC�X�Zj$�EId����T��zUg��C�Ie��F�IԚ��E.6��7��S�w���u��1#��3=�72k͸_�h��ocW^�7���hyc�o���DdLքLK����
�T|�������8��q݄I�GSϩbؙ�p��mlJ���j��8*�.d��]���7�F�A+��-�2�|�v?���/��(��E��K�� 9���{�$��1 �}����Mf�u��8�^�s���k	��7��\�9$⋫���A�LU-��ط�������-���l��~��ZB���aI �5N���(>m�O?�odԳ-mu��۞3/
�R!Mc���tGZ�'�.�$��j?�@���0�Tp������m��܂�/C��7���2T>�Y�����0lQ%HX����e}��?���n��b���>dL8:����;�@p�
�H�|
1��iw�V�BN�f�o��=�)s8f~��4r̴碗�.6�+TH2$࿃IEe_C��)��������2Q�P��+G��L��J\���rY����a�����w!�*��z ,i0%�h���b�g�O�KhA���Q,�(oH�M�t���0ׄ\�#6uw����νa�9�t�d4W�%
I	�H�c,�i���Y��� \F���B��Ln>)?�11���D&����>n��G����Q�h��]�ѳ�Z ��l-x�������%jZ�h]�"���YΩY(D8�V���FCM��_�W���ĭ� �g�8%9I���q�5���1��a�N�!�q��T�x��T�j]*I[���r ڗ��M��Q�0`�}�����*Sy�4Z���t9���L	tz_DkJ|�R1��)V�m(��b/��s&��r�ܸ7�4$egl�^�K��%�E�������b{~�-:�/��u�7�"e�MNr����w��p_����] ǂ)� ���'̚⪽vJo	A������N,b���)�qj�Vt<�0E��jb_�tƽ���-�9������P�6��)�IԌ8��;B����vUN�~֎rC�����$[��h+ܵ@7 y��^�����O��1L���^0�m�pF	�9���	(���Yc�#�Ћ�aA�ѳ��*�.�&h��0zT{};[��}D�x��m�5E�z-�c����a���>������!$�X��w�`V�B���x����'D�h��,R���z<�m0�.�7�����\j�d�+�JI?��'$H�.�G��z�	��x'��=r�<B�a�����S(�/���b�N4���l�"?��vb�j��������9�ߥk��V�_ A����HY�����"�n�k�q�WQv�D)�Jw�0��2ϳ�^-���v�t�P�j�/ʰ.7g[["��Q�CdW����ҙ�D���:����Ԧ��nx,���3�s�j�3���MR�4��F�|���4�Q�(���,!At�o~�څs��;��|��^+��*�@���E`�	�My�x����BU��݆M�����B4������ju�k�Ǫ�w�/����L��#����U��o�o�u+E[\1���d�Tm���qŌ��%7^K!���*��H_��n����3%!�	_V�,0���\��w�$�\��d��,�Aψ]����#�I��LYT�X���B_�w䈏JxW}�
����`�S��_Q};� �Ւ#1����ۯZ�%%H��W���G)ܗ�֔��G�/�$��p�VM����,�w��k�{�2�o���CXGlh�,���TD�N�%f�[����n��.)��X�O
Ԁh��Ť��Ѿimn�S'��M��9UC�+��Q�|G��#�0�v�����sA)�Kk��X#!�D�u�O��,���f�tl�+
A���oRJ�{��᫃c���^�����{�`�~��G�Q0�������_�����@��w�D�M9J&�|�e�f��[WT�'��|�Q\�e��?��O��Q�ug���!y���%qķ�l�j��术8�h�]9w�h
��T�u�� s�k[���Nڍ���h�B��EC�Jv�=����
���R��w����\���KM���r�i��H�#
��d�[��(9 ���W&&�@��XC0?s��J�? �m�*�ܾ-)s�����2�bA�JwgJ��غ^8"s�/+h<�>� ow>��g�l�G���g���0A�
�H�6�:��6VT�t2��+zH�C2]ld�5���t���w#E�ؕnt�7*�Ck�����0N����nm������3]@�@�.�pBޙi[{H�<����xJ�S��ɢ&�}u���N1x��d�k��Ƃ	0���w��'�ƪl�L`|�'���K9���u�5W�<'�c6�g�F�q�4
+��/<z�0��Ob�_Z���U���Zt�ſ�*��;��]�L|�j���A_o���2]�,�)?3TOЭ�g���e�\�Z%��TL^T*`D����T�)��|-T�^\,���3���n�Ĩ����=�4�0鮊X�+V�L��r�����3�6��� Y����;[R�k�kr��f6����� ��J��l퟼�:�h���׵JJF�W��$?�qG��������xK��5��xslq,�jv� r�B��1��+���؎qeԲ�����<tj� 7]���8���y���,�:��-hh��^)2��яEÊ�ƅ,��'b�n�/���+���U�1GI
n�	���[�0�ؔs�$����;�S�tM�0A�|I*���'[/I��C� N�c�ks���xx�#m���мOR�6�������0���7#�ǝp��1��k6��8�M�@T�xh+��j+�T+��)�fHT���V������6�⒒�M�9u�Nd؀؋c��Vl���� ��WЋ�j��EX�7 Ҩ�]Ho����?16p�;d���wL��K��LD��	>��dG���a.^kي��S ��
�����.��jo�c�+�xY���&���3���n��X(�ۋs̡%��~�!����H�	�c�����d�
_�A�bK�I��2�~��zpgcKj