��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�i��a
Α1S%� �uj?�L�3��TLei-3^5]E�$�ԓ��_�d�탴�,���yN(��"]�@ % T��U{��"�[.c5�\���J$C�f�4c	'J\c8�a)B�M�:H��g��TW���B*�_���Ƭ;��@ƨ]G!������9��J���a����f�R����I�Lw!:Y��#!C�����   ���\�8�J*�O�ϬpP�KoWY�x#��9׹W�"����K̇si)_��aΛ��m?�q�
y��װ�w�.�/R���!à�m����ˆ���>&�z��=�	��=bӥ��J (AkF�����%���T�	pΫ�\I�Q;Ӌ��ف�\��Tْr�@� ��z��Ep���/����|���qJ�Xl��/8�P�}7w���AAh\���
������.��<�#�yTAP޴^� �x��\aDn�.<M �7��
�"̤P�!Z��ti ���u�Tẗ́�j�/� �q��GlmK���P��PO�3t^���������Py�i�����Ԧ㡡�=uG�Z����Wd�h��|0�7#�7xzŪULfH�?$�H �f��Y;0��e��DZ4�V��� !ߔ�/�-�G�}M�X���	�ɿf�\�bet��y L�� %�1xG���{�nZ͐M�+Æ�i�dE"��b3��F��~D�;������d�����'�]���s���o�ȩ�V� �O��s;���y�:�L�p,!l��K����7�K lN�؈�|��X�R?��e����(>	2W�d(0l�2Z��"x�)��)���"0���QK��!����/�.����陁����1O+��a�{t�H��_�P�eYc�(>z%Z&	�'R����CL��1�
۽!����V��|�cg���g�_h_	QO��]�]YH@��t
<��Cd�D��=򛜧k5 ��J�A�a����^��㤆�$?��p���*G9W�OK�oB���\朅����0�מ8l3/��P���:����y��Ś@�VöcA��pR�]��Ǡm�:����Ok�jy�>��2i����b ��[�����r�+�� ����o�k�V�"�Y�����wT�@�����Tv�6���l\�K�S�.4���kug;-�	�ָc؋Pj���F]�3��sAe���3-��J�:! iw3	��a��%���<��9wH�~��_�;h�۫�`N1.M�}uG�j�5q�=�\�W��^߳�j{$��^�aU���d]W�����v_���V�zx脄�[�Bԗ�x$�2��(��Hz?~��1u���j���C��O�2<E!���75����*}�p�2g���U~��p��q�=���Ѧ|���3���G��n�xm-���!S�ೂ���?��->��Z=���loi��Ĝ9z+ؗUi�g�\�z����;5K�p���U�(�}�Ub���{QEA�j-o4W����1����2ĆxO�|�� �r[���.7w�J�_ &l�6�������ő����u��S�6���=�\B? IU�>>��@RѶ��Gx'��Y�w�/�tQ����x����h1�Ń���'����ռB�Ä~���ie��h-��R��~����Ⱦh
:��F:�Ҧ�C�q���MJ�����|ݰ3�b¨����A�V�}�� $Ʈ>v�J3�p�a�Y��*���'B���~�^������!$���Ia�����8�V6����Xx��W-p�y~����7���b*���,��S�������&DT�I��B�)��Q��;W�����ņ��fFv<�Y�����[��t0d.$jz��i[z�.k�����&N���'a��(~t�����;V%n�2w,C2�ޯ����?v�.$�W��(N����c�� nV�L�#YgoN3�[�xTy#����0ܔm`��G1�����KϷt*���@V���<1��SOXJ
�9;b�w���j�m�DѬ��#}��"�>��-�:k�Nl>Nt��"m�;
U�z���N�4>ѣ��'�:�<X�S�1	���f�1��&~6.#̺���!8��C�=�=\@G�w��������s�w��}֤,��DiLW��T�R�^O�ؖh�ς����*Lz)�^��ZW���Ш}�^�)��Ad�2iӕ����00fi>+Z��O歛HCŴ�(��ۜ]�Z�bT�)M������bz�m���]��1��$�2qz��}����7u�� 8�T,$ݞ�%Ώ��&��vG�`>��16�"C�����Ya�>��x�}���$!�*Z��t=�A�cn�!�D��
pcA���Zk��k�,��"FP��}�{��G;��taz��a������w��f��f�|S�6v�qk�W�x�K�s�\Ɂ0a���c�����%�'��+���^Y�rV1�y��`w]	8����<��p=t����q�d�$ew�>���<�E��{]Qix��&�nY�I����rt���W�����Y�'�hX|���؛�W������v7G�#)����bPg��p]��JѮ��*���K)C`֧0�H
ͫ�l/������D5�����_KzN�-���1�xf�0�^�A�}J�4mT����q!�+�"�P��Ռ��el���V����D�lT���u�f�GQ��"IT��㤀zM'X@Y\����`4JD�+��O��k���o�z=$c���[ʚ�����s,|�J@j�{��r�Q��+���3?��L���� _�fd}	�Y�pN�)��{��yG�*"�6�i�n�VM����ջ�x�h44���R1%L�`�l�41M��s+�G��;*��~�4Wq��*|�y.�^:��m&{\��SK
4��a;���V���*��?՞|;DdPP
�*�s��`'�
�F����Ʋ���b8bFz�Xh����U�_"�V#��հ����G�d����߿���db�M|;al�8�t�IS�"nMo���-u���$�%��g9�|:��.﮶����!<؂���Ս�J3	�����J�D-M�ƟN�I�0�������KwK�9�5/������OC�ٟj�`��/�X����!�S`�7V6������R�Hm���X)7�1��1�Dg�	dU��Ǉ��[��%�9{ۊ[��IL����Q����sKM�N��?�����{����,���TN�H�Ts\kW',��~�U�R��af���~Ҽ]�Zl�]�.�����fQ���_�5�V�Q�rzBDՙ���ژb"/�����DҋԎ�`�<��e�fN-˱ő���u4ϋ�B�%O�k
&�	�|�*?�ZJ�ڷ~�K��!"��hI�Z�ۑv�f��վ�o��(�g��?�b��f��F|��A�* c5_r������]���lڐ�  މ%����;��u�Wi��PYQΐ*i���`�u&⋿4( �ͼ�*��U����F��d|.t��z�r��i�(���$DJl�$h�O*��(q;���7��/�Z,�y�uĢ�����1+7�R���(���Dj��6"�d���U������	�5�G���Ba9�#������W���Ж� �(&Z �H�B�m�N'�8��GǷoq���&ː7���`�eR�u���(�*`���N���O9����!*��6K�;�0���\��aJ��$�rt�F���x^�o �S�8�U��;�i{W�qNG<��@�u�nDl� �2no�?]�����V
�dy�0��q���=A�Ӯ��ŗ!5+єo���@_�pB�|�i�w)�V���F��D5(F/��B�{�>��y��d0!KK����qpN>ju,I�lIl�J���Xl(}�܋N/���vMg��ؕ�)�:'X��V�'v�..C����@���a��>�k���I_B�2����]��̛���ZpFJ��yU�)��D�M��S�н����$Ɛ�$�F��	�l'j��4�a�JyO���״������!�~�����T���y�oI~����K�
�Ͳ�D���k��0
��#�4�~Z��	��9���=�7}n��b�/�
+���O>�7ƥ�dv^i_"ф�Z|{��4�6G���֐�l�p��K|�{�`��*�A�Jxrvum�Dh��i�Y�g=h{9�Z��F�L��2�$�I�|�8�?!-|H�#��=Zm�n],�<�6k^����͵iz1[�UN�a���L�W�R/1��X!�p��m���sA��ވ��s�yV��r��V/�;���c�j��������^=,}:��إ��H�B�=���
_�eⷤhtA�_�(�
�� 9[�3L��f����K���R��=��&�)}�ǚVk!��D�H�C馁9��k���O�i��+�u�&,q�T�|��K�o�<g�ɧ��is�����ꯠ2e.X.i��`��u�g��e�"��d�e=\�0�qڢ�R�~����n;�Z���|�擣����gpm;�kh��6�;%ՙ�:�=E=����$�b��$�{p|^���8#m\"�ws�E�'�>DE���%L�B�Q������`�S�``����1�/��k7k)Kh�V��*���c���I�M����❆��	�f��o�$� �� L,�VqF�	����K3<eN˔o�B���R��n%ڞtjYzޥab]C�.�|;�c��-T;��؈*�����؎(�W�0'�\O1*D�j%,Ye�ȳS�g�TY4��.N"B~�aOZ#���1��A�����)��R�Z1[[P�RɴWpA�n<`�H ��f�gw�K� A�;�bD��{�rxN�b�q-�����,q�vl}�v_���(]��D����j�YK��X�Mac@3��Ƕ�r�p����Z �sD����FX'�I����)�����0�M�p���^�^�K`�x4ib����#+Mʮ����oM���n�n{�ܾD{��b� os�@
��+g��V7(R_���}(6�$�_��,�441��|1�x=t6�Kv��0�>S=_���p��R#S��L����Ϗ�Z�sL����t�u�k_h'�B�ĉ�I,O�`�/���9��~�ak�_W�`�))U֞��� I
��zm�IX��V$�OGT�W���cS��uG d/���)��ƣ�Dơ����3N.���e0��d�M�p�	h�雉�Њ��~���h��Hi�#g��"�{K��`�OrK�;���m��S{#�o�W���喿k��Ģàc6��' r�Uf��3����
�ҡ�#U�1�����U�&�N,��:g����L�$��11���){+e�޵"U2
�ذ(�$+�Tl5G]�qٹ[��i�m�!cZȷ�F#{�4�:�Ҝ^�2].E�����︦�-�8�%���P�� ����&q�U�q�I�c�$�8�D����
{�7��D&)���i�|2:>�1��ptT�K�y�����¿�֎z� l���%�I88$H��m�d���7�D��mO�y��:��l������#���t�+c��˳��b��!~ٔ���~��T���˟÷Дj(Y<��@Β�x>:fx�bF�?�O|��{b�rm�/��V�S�-�����EJ�	��Qu�+�Q4J���.K�\�Z�^�C����J��)o�As�+<ll�42�^R�j�'�C�ݝ�<�2��b�]�6�Q�+�	w~��?e7�U��0L�Л엺���N� �; ⿣����¨�c3��h!Mk���X���\xiu)�7�=��b~w���\��b3������c)Ux���P<�.KeZ�~�S c�ֺtW�Ŵ���Ot�w�<��Q����Q:m�2a��ɽ�JL��,|�qB)2���V7N^R5t�a���{-�h	������ЄO�7�ЗQf߭��a�e�2VEf!�Rg�Er�����vr�08�7�h�3D'zG�s�X�Ϲ����|{3��.&�^Z��\@V򞬬k�XH6�#�Q?�crI5?Z��/?Iʲ^N�	ȭ�v����3G�ɲ!����^�����h��G� T}��t%l��j��\+a zs��B6� ���sJkv�/�h9�e��J4�����kzj=���_�['�	*u�~E{��!�;E��ȸ��r�i>}�0��O/��k����-Ne���|?YpB VN�F�����ƀ�OXU���kc�����|�-��n �O�B%E/�(�J��l%A�{�t^`t�L#PGxq�=����,��h#-���W)괽g0���V튊b�W�*��@���  � _�їp��ޯ�	�n��:}���V�,n\��r�́ڙ߯?u0�o���/H�S�u�hPZ(�dߨ��l%A�Xguz�pX���ދ���]wl��mi�`iu��jV9���j�'�A�7YD�vw�U�4��2�#�6iZQ�M<Eܺeu���v���z $�j�nEœ��=��F��V�1��e��ܻ8l�C��3Rc�=�ċ��!r�n���S6\v���g�j���k���վ�}��C�)�{��C�ǳ|��S�d�L6�aH`m���3HȂX>��v���*-<�;xE��n��nCl���N��F<����6�F���u<�٘�κ0cjy���������{-x[j��[l��~���
���M,B�~��,<������~\����h�	$����Iv�2�+.�]�o��k������z�щx4eMny���u��ʳ����[p]��5$Ѿ�k��m�X��0LD,}�������O,'�X�G��0�.C���.3�ڨU!�$;y�V<N�+ی�����a9��tv�a~��E?��fl)�ò����]�;�,�괿�
��![����:��\k���Pq�j\��t` �҄�\��
�H(tOC�$ynuS��!1C7޶69�	H���sg��~���ۡ�&�p�ۅ6_�  	�!}��;�������T������p�-⸸�b�5���d~
��-�p^Ǫ�ȁ7gcȏ8[A���|�?s�p�����L�+P�c�In��N�ؠ�3�ȭ����I�9��Qp��o�G�R-���3�_z0a�02��ahc�?��`U��{�/v��Q������ �F�߸��o�K@V����`����r^�{�B�lU�J�BW��5h޳�~hå�>QnL�.P�������a�~P��\�݉i�*6��Q<��{�����o0�s�x3f���Z����9+�����T'<�W�O�w9l᱂kS�E���M��#�������n���̿�d�����բdX6���!	���Ϳ�I�v���G����]*B��MS|��!���89��M��#�W"�k3ۘ5�S�"������g�M3?6S����Y��oG�)a���A�V�#e�y�E>w��Y�^4�ô�h��i7t%<K�Tk��y��{�#J�7;���}�u��Җ�P0<ɒ|��v�5%c�0)�Fy?�4?a����Z�x�&88�u'��9KͲ�a�)� �����f�~�w4��o2<��Caʭ�t[�ϒ�˒A�p;�I&��L �� Ӂ�u��Z�@G��Ņ�h1�k�k!}�L�"�lϭ�r"K��B)ӫ�%�DR!xY�{8IUF��hշ�XM��e����w�C��w�D�y� �����FN�F�d�!�	X�%k����o���/A���_��I�G�|�<$\S��a��'^�BK4��t�($�jK��du�=i��{ހ+�G��9�
L�2��<�>P�ܠ>�k��T��cEO�r�tF�*q�~u5�	��Uq�uF-MCK�ϗ�=����RY��.bN_�q[=Q�@��P�������?�t����u�*��~�wNa�ƒ���mA�멾��*�������M����q8w�	��8��6���m�¢���i��`�|�63oi�*I���ǋ�ՠ�g?;A�r���j��n1���JE�Пӎ~A��jOÎ8��r#&�V]W�J� G�U��H_��X5D@����4(����7K���|D\>��k%����V�*��:(0ڈ��1ȭ`L��淐a_�X:����@3��?�4D���U�TYd	���2f���L�@L ��_�~���u[�=��2���9=�3-VG<%�9p|�Po�0�����z%��S�lv`k�`0�I���(�R%����cÌ'$H��{�U&.�����1����Ҫڋ(2O#L�,�[�rW+��Q��0���rG��g\;s���+,]6��Cȶ�F���Q���V���;�|U}��҈�"q	�Hh��&�]�.ė�X�D���-��v��8D��|^�a�2í���'MY�ue%�G/L�CՉN�է�/zKPf���O�z��Yh��UH��ృ�y���Qj�Y�VN)SQy{ieE�i�q���U�o�}1�9A�T��`* ���mg�5��'��M����(,Y܊@t6��3�*!ҝ�4sF�Z�,8�����I�ZI��?,ۏ�}���G��?�F�~��]����a7��*����HL��@�r�?�_]�Ɨ"���GV)?q���]��{'�+�(�R��H$�y��t�wK4t��B�+���J���|�2�i���X+\�r�gH���-�=r�ۨM(��,��5	W��Iz�KP�	�q�d�l}��&�ަUaԦL��3h�����[�v"�sy'�el
���6��
��I���ӌ�B���Pc:�0d'w�b��J\�"R�zP͈��A���Fr*G��ZFa�n�4�5}��"�i��+J� �����V�]����,��TҞ��,�����X0v�X�	��ٻ��b�1�޲l�W��.o�f&eu$��Q=�+=�Ӧ� ��B"K<1'eL�8��w�w\rzduv�)�����f�
>x�2�ޥ-�g�!˕����(G�D���ňj�M��,C��Dj@�s�kRB��U�u	���'�l�?j�V���}�7�KW�@�𐒳Q䣍�eA�IFmi��;N��W�K��O[�cC._�l�}9�:d�a���K� ^�D�=Nm3�D�&U5������JK�*��]��YÚ���U��@�88ad13^��J󧉓�����)���v�
�e�4),\�1eUL%��/�d�3��igx�]�<�p�ї���"�5sn@�Җ�G#."��D@�L2�C��:wT ���#���3�5>]ę�h��f�O������dYF�wA:J\ŉ�<���'�<��,^�.��es>���\�"�w��$��f���'w�_����8I�5�cK�@�$�5�{�C�(�Tԙ���k��Q���)	�d�]�F��ȃ�P��4O��"�^�9� �\[����_���'ݲ�-��0��2����}k���_ȇ"�Lm����|�����Tg�I�F-c�Ff�ݬ��59�~��C�~�]�!	{��Cw�e���]L3��N��Rb��◯����hF�c����?��m�(i���g������
���\�x��&���S\cC^�hX}:��c��n8�ͅ�I�k�><��F���&��'_�S{��U��~��. al�m#�i�&�GI[UJ�����jmm���B�7�@:L0H�D?���`�B��x��u[�����g��])�N�8��k�FP�p��*�g�_��o��v�iM���1��P$�f�ޚf�S�󣪗S�����,�$$i��"IܵM��uƪ�5�CpuA��
�z̴yq6U�^;3�h�>�0k�c*%p�H����E�ưy`��5e?��k7��<EC�.ʛ�L�j�&9_�'����'<A�#n�Ҝ�,fC�t�}gh��>��Ȁ��mP�C��d���D��}�����u1J���R�;�B�}.��D�����E��Xyx��a
D� ^z.�!��ޚà�a��.��	��E�ҙ��R�x=n��g���#M,e�!��xm�ٗ���*�G��g�`�u��v46�����(k�o�l�/���V�{��	W-�E���1�g����-@�$�q�ωԄ8,��r����L�c��i{3Ř������ۘ+���޴K�e+
�d$�WǢ+aGm�7FI$?����fb�E��RW��Y�`�с4�/�Z�)�nB�M^*��]f�E��.��3����9 iD+َ/�K]D�uA�Ս���
��MS� CE;���*�~���Ԝy�r����M��Hl�~L����Z���v-c��rLt9�FR%UvI��8�ZF=�'{"/���m��zϾ�_8|�R��O]������j]�$�Q���!3柲)Q^`�g7���r� ���Rp�K��V��<-Ѯ$2�:��๱D�t6o�4��~�.!�\"��
�}����U�S��0�k��s��C�(�Mk�Y�<��K���i-�ns�\U�ν��:�z�>Sw�6+c�s|>#��ӡ~l��7�_�[<���� bE�no�!6W�F�Q�ź/޳7���� ��m����<�������$v�>����T��u�	�qu��A��5���T�'G�lC3�ං���L��ܦ�
������!�:ͨM^�D��e%�[��Ӑ��l��3�ᡦSn@"u��*g���e�o�5��/�]6�:c�����bd��@L�%��a�
�kw_R����9��"�?��L�t#���{� M��8�g�Z�W�I8}��)��X6w�:D�.�}:LS�`)\���܉ܖ��~Z�i��a��g�\_��$��IAQ5����B\��$��Z;�0j�>V����m]v�J���W���qGMP��&�Q8�n^��2�s��!'�>+; QyP%�2��5���0qq�+�2>�m	��GY�O���kg]FF�K�r����gY� '�(���˛�S��h�@�_���<)��`��o:��.K�5�U1n�#S>��{���Wϑ��qT/������+Fg�d�*^>�y��k�н�07Y�{�Ó_|�#7J'n��\gY�0���<6�?���bK�����F�QI�aT-	��;� $X���>�mI�T�zK�3uG�{�5k�yzf3[�����:�P�l�Sk��m��C� ���1Q���CyJ�6N
�ꭆ|�B���R\#9�	�_�[U]u�1����/�וw^K�T������8�������&��'¢�T:�X��ʗ���t
I�F����#PEx���%Д�\��ͬC	J#�_Pl*�+2&�[.��M_B�n��-y*���Do���R� D�?��§9�2�[i݃�=ybMTQ�L�������MVcON$φ\�`ó��O�H��cc���z?&��U�'�ɄA	�-k_SJ4B�vi���1�沛�:�'#p������T���c0U�k�s���f�9�:g��E�_��?]�v�VR�~�Ѳ�֐��1�n`!����%�:_;ۘ�����L��_�v�m�m˩@*L�r���P�a����-s:)�1�;�¼g�xABk�<zOK/�該�Kr��D������dQ�{��)������ď��#	������1r=��KHeH�S@�$�@�s�rʀQ�G62�R�M��_������q�;�+�K�����Ys@��(�)A۷�ȡ�eK���3��|4orz�����C�V�e�n9`�a�e�b��:�i`��O��e5�&=9dy�	˳�ih8�t��fSwَ�C�h����-:�V�*����#6�����ޗE���?0�Z&gO	�ź�E� ����E�Csd��N�v�]W%�{.D��!%]�LD?xo&*��� �R���Y�t� G��	cGU�k��7<�*]ĵ�c�2����-(Mz����}qL�r夜ʖ9�\�����o=�uƄ����$Y�5��D���t3��O�����]�*��`<��0:z������AyI��Ǐ6��l)2���^ՒH�PP�nAK����2�����>���&_�;��Sb��QOO"MaR�<�nDi:XJ��k�����O3���7�Id���b8t]���:y�*q+��ґ���~�KJ�0�ʙ?�DXas�iQ����K�R�/�]ە#6�"��1s�\���]�^*$�V�pO���Bz�U�4��5�S� q�0%{r��f�
�#����x@U�F�j�����ߠQ{L##������m/&z�\���圵b�p7 �,}$J'Ԁ�Պ�P�0������_K�����}�9����M��]�� ����l�G��<b���ƅ"L��S�Ej{�|�9
/�8��'��u�u4���H}6����&#ԙ�잾�����rc��{
"������e!Qe�k���u�vyka=�z��pѥ��y�}.�X2��}��uw�BgXv �e4`E�5��@z�z���I�6�-h�A�������G�]T�)5���`+Q�A�2I)n7� �`|���~�]*?��X.��U^;��l$1F_-�	t��?x�9���l����Ō��wP3jE����TE޺5���%�+
Ȫ5��5w(��]�����/�㲐q'���6���	X�<�=���j�2���?܁�t\�O_+��߯��7�S����	.��}����'asz�����(� ��5kw�.��Z��Qx�Z��p^�/�߃TVͰ李���W�d�o[?���k[{����<�rSQ^nI5��������
�i�i��Ţ�M#�����V?�K74��� A]�4S�c��jE�S8�!��\�wN���Q��ŗ6a�Y9��=D��t�w��-���gf!��{X�=��XGޫx�����Z�$�<=3��F�b-�B��J��[[��r����t��rM��F�}����x����e��Ym] ��7�'�4�D2�e��.I^~���o�d����ւ�:Y��8�e:�щ�ߥ�|򭠰�|��/�s?c�@Ɂ:���"#���U7"k�a�067R�7���B�W�H4h�͒S�}K�iX+ۊ6Ǥ�Z9[L�bi�ľU��W���L��m���U� i?�Lt��#⪣�"&aT]�Щ��9M�e�_��u6�L[���fS�_��v��vi���Q�k�%�w�>����Ŝ��<��7P#�:ڛ-O����Q,rV|Q���F�p��R@���#��3�2k��j�X�������,��1N3M`
�Y�7�����*��k�s��vl�F.��5׷?��L�ϩ�R0�����ioJ�yR�	� �a]�۸������c\?�oY���s����f&d"�U#�_6]��4+�S@�
U���J��c��|�)#���'�C�=��G�Ib��D���p�ݳ�^�̕��L#�k�~䀐�.I��3Zr+0�B��^�⯛�J���jʼU��N61�b��ם�}�`DPY&���9NC������Is]�8u�I��$�[�R�g:6����Ǿ%�̟0�f�_��s	f��.'Lg7��2�R�`ׯ���%��u�訯`�	��֩���������14^�,&��Yٿ�,g��k�c_�͂������$ծ+*/��~ێ�d��X�, ��}�@	ӣ��9
Z��p����,A�T��/��$� ku��b
��Z���ъ�����;���|i��.���z6$��`x��|߯�Q��8����E)4�P�{�E����s�R�TS1h��?������qqy�0������?g��>�䋠�Ɵxͩ�4��;�������C/7���K��G�� ��+̻���I��7��]�6?s=�b� Sp������5!Y�ZY�H�eU��2��.JbC%BSͥi�QR2����/��Z�՚�Q��:@�d���[��� �q�����5n�#"�3�%�Ӝ?�9�i��K�Ԏ�� �w۔�q�: ���5���n ���>�$1��W�^T��}g��z6�q�^���EA
P�Md�^�"��f锎�Q��f��2�:�,֖�k�e��W��b i�R����:�l��L�S'�I���%�8H"0�����R�8�p��Rta<��!�)уCXQږ7�A�r�J�'����T��&�ₒ֏��"��Fa@�'�Z�2��>R�=�aٻX�$����z��u�z߬(o�ټ�|X��44N�	/���ƃL:���3��$$�����+�*�ڎ�x˯�QDs��R�B��%P}�����G��\2W$�uftI���c�"�ţ�J� ֛�G��ʷ��A�c{��R�Y��岲DkV@Ss�k�� �z��&i��MmM�D��\����bҙd��qp��v��\m|6�h?ej;@��-�mH'`M�3��<��|�i9����T-4�}uǢ7`�g)��Ip��)����lq��.ٮ_�4g���h��\_��u���.7,�s�Wf���Sk����p�t����S��c/��$�h8ޙ��z�.(F�)]��&=��r�l�ҟ���_n?A��?K��������Wt����Րl������h�/�ɚ��<���<����8S���W��Ø��K-'#�B��J��̴�ď��=�b�!U#A��r��w��n��FZ�\BB����s&7At�!�1G�,"dgHz�p����X���I�8)��h�]�~ڙ��Nq�yV�+��WS�G���
e����".nwb#��t�b���S����~�.�N���_��3�Vg߃�C@d�N���P�]o��.,S~˖� ��Z��
<����N; ���*L�e�|t��]C4쳧(X�]g�!Pʽ��V�7��^��]>�M�L� Sl`�6�ޑ&A����[�qx�`� b5����Z���U��H���L j�u��9�]��C���Q��������"��'Č]Ko�ގ~�q�ڐ��>��ˁ��w�p�Xm!�)۶>���z~��R߉�a/��L܍ԖUU?����iWJ�kW7�.�H�)�JE՛�6�>��Dw��!�(� ��d����������b�������/n�$����}�� -��[��Ygtt��юS�^!ql��Q�6�[3���1ώ�_\�����A����.0�6_ߗ�d'��ҩ<a��ў1�d����Q(XV�;LCmp�R����q*�_Ѭ��Ǯk}"�Tƺ���K�:O�H��k�ۋ�B�/M��_�:�V0�Jg�̙���L�'��Z�,�#P�Z�=�Rև�k�lX�1d�vc�^�KAEH�S:�k���顭Se�-�p5g�w������NP�Ȇ�T��P]�� ?�9���tڲ3���%­xx��v��v����B�K\0�N�]�-'GW��?��4�'�h{�AJWG�ʼ���j�Q����N A,!) ����a�=1��%u^H�:��87���_OWz��zS�w�c���exAIh���q�%�~=^<D"&Yܦg�*�~��=d��%����u�G��#O����Fl�cU�U����R'�q�6oa�ɟ��P5�Ih����V���%���ePGc[�s��.���)"��D
i|��
�6�߳|�^$�c]�ڼ��aѓ�/S�&1�x�liY�4c�`o���+��I��}>��.��q�T��oߏ=�ыj���m�.�}���$�[��p���w�t,ln0����֭�P
��g��(՝kI��� r�wJ���s-i�r�� ݅G ���ߥ�Xn ��1a�^ih��H�Ni��{��z�`�h`�~h�f�6x5Ũ�T�9-�%Vֳq|ז�1hـjc���͘ڤJ�����4I�X3�?�)|�KqN�C�'P?w��G�_b�Z k��b��-J��8oT˄�ٵ��/{��oY�_�HO'
ep�?N�~񴜬:��{X̯w�X�&��a*���-��xQ���Q����n�ae�^����)$��F̡3#V`��%�7e�׻����WBUZ���
OΖձ�q+thOf���ux����K4T+%�ax�ׂ�ӑD�4 ��� �dA����q�&������G�fXkJR+>Y+pYP:v O� ���6��t��)�]�D��ot�[>d?:�~���Ub�(���~BL͝��ǅ�1Y5Fe��z���J��.�T�� �g���WgB���&���L���j'ܙEũLK�����.;<=��h��*�MjT{E�'�[��>�?\�+��rؑG'[QX��<+$��:{�n��{�����T pǩw��� <Z#D��I���&�=�%�xd~y�M�㓴�6��aJy[�/����bR&�VgH�B�\4KĦ�ݗ�Cb&<�]a��eb@���ۥ�f����B��k]L��FZhٖW�#Q�{n8�����:����oyZ���+�
��a`XD�
!��Wd]��$��|��.��w2�c\��v L���/� |��B�b�v�P�k�s�¼ޘr����;&�J��r]���ֵ���$�)y���l�KZxe�-`��J[]����+D���%���G���ք~�/vP��@�|:��n{���f)�YY���&=/%�K	G�xƍ�gw�*q��Av-^kHw���H��=�Z�"�Mm�ű����(c�� ��i�b�!`����"g��+ �~��ym�T/1E�o�]K=;�ζ�xi�c�;ꝺ,�\VC+y^��<k��Pr�n��Le��~�BUd�	8�����%rG�@�㓳NtR
o�}�䆴�����<�R�sF��RDo;J�?(}]ܵ,�x,��H�:�{�oZ;���RK8̊Z�q�y��N����݊&k�0q��'���
��*Q�/I�h�&�"���1����t��5���/Q*>ɣ�zX��K��G�O�Xϭ���J����a�<L�dV�ͨk|���f!c��P8���8��8h�G��۟+x�j��Y�����3������" �D���b8��h��s�^�4fs�>�Kј��l2tWB5<�����}��r�7}��I�#o�M<�s��\�M� ��h<J�Ł4�?�"��-\�6q���>ו��ٙ���BR��k�9\Pk�]�˚S��� h١�s�)�>U�e�h��b�M�)b���]���|�}��̷���x�.���]/��<���tbV�{"��h��Ur��$���(^�R2���C1�ߑ�K��)��l�?�8vـV�<7��ﯸ1�/�QЇm&����?��&��	���D0b�<�bU�w*�W혪���zm9� ��3�/���>�|l���p���=�ɘ9�I鶶�rAu��J0qUJf����F��,6�^.�M�~�%_���<�UMZ������T�
�C2�ё7B�;[�� N���7*�ƺ�_�;�:��LA:,처�ǆ0�ȅ�9�u��K��H�~��>�W���-}�O�)6%i @��pB鿤"�1���	'��$��dδA[m>��<���Ă�pͬ��w�#�4I�\FY�Rv�F�3i=�ce�v��5Z-�5����9M���p�0"�-`��>���b��G:��4��'�3����%Is����!���E�<A�ߚE�+ݍY�w��d����'�І�:�4���G-1�U� h�����(ޓ���?Ӻ��N��b��h~{���n7hJE+�3�s�g]D�h_��nB]��K��?����x�+����~k�y2�l���v�ɻ_j[���}Y����)PN��CC;I�Fu�U�=���l�7L� ��N��O��MZ�É}ƻ���Ѝ��t�x�mਂLu�~��n(������xT�����X���#�c<����Ŗ:`ZGe5pcD��M'�>������~�2>=2�\&?QVU>�����pl,�� z/�}��1���I�'q$a�Ev9��wUװ�%�d*sU���2�8��e��_ �r���8<>\<��<G܌{�,~{I�sPK8a��/�;q>����g�i�l����D��IT߷��]_L���O���Z�'Gy�ՙ�n�{���V���ߢ�=�J�Y\Ņ�LԺ8R,*�(��M��)F�;|�'�-�Y4���0�j�k틛�zs���s ��R==8��J"N�d;N����cR�xm,�����i�.��e��~iY����ơQ���q�4���-<�&B��.`�y^:�E10����G�T�Z���m�����s!��@�<�x����F�oi�q�Xq�Zβ�%o�;�E��W��n0=|�*�2/W�eSk�u��N�l�9$m����&�Yq1�1���y�K����g+s*U�cx�ë�u���P`c6�"�����0E��j��u�������*^�<ϳ����ba����(T���R��I�,Մ ���u#��5��L�/.������c���TLZܻ�R'F`��%�E�Cc����е����H7/jk�L8aT�˵E���F�����!"jݥ�qf�2��EG��r��e���vlSr��^|�veg���%�%>}4J1��d�#� ��$���	��.���n��6�u�D0\�f۳�I�C|�K��.�y\�ٟ���XF��ceg] ]Zk�����<r��9�8]>�|Ԁ�۬@Xɑ�%�����4{xTh?�\���G���mz�o8s,�6��#dB�mT��@gǵ��g�Kk�Y�m��4m?�������,�)h-*q���3�К��Qu~���� �V���
�fl��� �ʟ0'`�W�%��9�!��L��A��&�ۑ'"��N_�f�$�@����GdT�/���&m�˽bq^�y3^�Ċy��d�e@3Y�C���^����#��C+mM���6(W�R�:0�s����Q�z�D��$�W-&y�%�,��n{�ґ �'^�k��U�,�ߗ�GP��e�,�2���;�E����[I.)���݋�.�����s�&#u�����t?D����l�� �
	D��x�;�qCH2:�]ݐ����b6b*%���p�Uﳲ��t~�X�B�ܻ��LT�>�� i�M'�L.�¤���<Nu��,���nu���e�1ǽ����A~a�IPRM#�,��T�d�gM{;co����w�Z{��W�fLL4�ܘQ����8^*��$�6�|��t>��� ���n�>$:Ί<6�c(K/H$���".� �:5hk���n�>�$n}@�_��%���gR���ң�E�k��i����!S��ZC�y��q#�]�_����������}-�d=Z�/'g�8����y�W� N���I�1yM�����a���2j�[w�b��փK��]��c�:�0�U+q���+�W
���>kԦ^3t�A�T�f3�}��;���Z/.�N:�Q���궙��|�9���Ҍ�m+gv����)��^�A�]�dё0��.\�mn�x�L��g�����u���-���9;r���������.�.�����)��,�� �'
R��"�A�5�?G�)6�9JX��"�?�ℇ��ѵ����AV�β*ZO�Xe�,�H!&=~�U\���@ W�������?Ϩ��0��Ȗ��1����7b�a%��j*=,���Ѭ�d��d|k�w_7�o�V{mn)s0t��Bc8�5��t�=?���0J0�x�J��P�����*���4P��'ސn�x2��Z  �ī�S��Ղ��`d9�<i����U]X'=����կ�N3��xQ�K���}oM�;:+9�P�hJQV�k��pZ�@���U���³���=�NT���o!cŇ����U;��^��w2���!�_�ܓ�"���qXhS~��������*��Pϭ�����p��_ˊM`@ ���A�Y44�	��+4��ua$xy�)È��w��pK��2��{�{k��B�z1cB����i8|�0��������|��m�|ܻ�b2Ķ�3�?:�<�ҷsl����<i�Krk�ejR��ƪ��3j��~T��@��g�`����@�\l0��0�����m� !x	� �&<+�9�;��m3Eso_W�4Z�S�kl/�'Oe�uu�>"�檅ڔQ�"a�e]�	�g�m/@4���$�N�}�z}<#�uM�*º:�t1���i��
㶩V,��F������沮V3ϲ$oP+>S���/zJ��e5iPC5_��et*��6�%���T����F��3� ���9�[�j4���K?v��M��S�c?�a����e*&��}�urKg^� �{�b�����ݺ�֕)�򴭆�w�Q'eq��\��(㰰���o����L��l��_�e�ՓK���Z�eHR�qPOy�������j�a�%�[�*����u��bi�G�͘nh^mۋ� j&����24���;�zI՝⢴qU�X.`�[~"�Yi T�]�AX�
tY�aM��j450*�ȹ�L'!�i��F�L�9jE�D-)Є^���������X�y=�Z��F�Un�������ƽV=��=jV҆^|Q� �N��x��vyӜ���IC���I[Ʒ+�զ�/�_I�RX)|P񗡷� }��������˹���p���a{J��� ��G�c�z�V�F�6Uֻ��uHRyiJ(qT�e=
� /sjc�T&���@��"쯉��L-(�Y��F�����6Ҽ�����@
uf�*z �]%�m+@g�J����>`p���zx�Ā�h��§Ooq��X-fO����4�9�T����@����2�bx�ia6R�ᩧڶio�Dg�B��b��Y���	mk�7�/�<�_�Px���6�LT�h��K/��\ �beP*��<�ճ�P a��F ���Iѽ�
�Ro��HQ.v������}�pu������]`&�,�	�����a���~:��&cS��<�ɏP�����n�u�N�-
�1�Lh��䳗z�p��&b��պk�O�FN������;�w=��khx�;ʳя�#��Dw���djJV� `�,��Kyn�tW�uz��>���Ա��\���?T����#�g ��7��C{x�1��x�8XCP�zgCW;Mq�t�P�PϚ�5P�6��n\$���@����Y_j,Xte���|p���@����8O���y8O2,���p;fK�y�Z�r§W�H�I��+���������6t؃� �P^�n`���M,Ԇ`$z,���&��/�0�*�.ʾ#�`V-;<�Wf:�������	%�`��o�Ds����)Fw�KG���NMS����M��L�kU{|��A�9�G]�U�ޭPg �R򰀝�����j~��?��E7zח��Ra����=SY�����fLdUX��L�o��8��wI\��K���eÿ3}���MF��/�0Y��p)�C�������c��� �=��F��!~���.�U��l^%�I��F�zpP�8WΙTɂ�7��b�K���/��D�T���z������t�H�@��6�@}p@��*	�a]�s��#�;^���}���w� (
���Z�t��fGh�"�����^����r���r+<��Drq���]$" u���m���<���9�3���@��Ȁ����"�U3
{��)�����j�wT[�&9Ț���PPDT0Z�G� �fH&g0`@��Hu��EG.��p�� 7y��5�(�w�ܙ�N�O �,_�(����O�n��5�5�0��E������� �H��gh���v�F�����5찖���q������%�ϋHQ��p��X��Jz���E��6��«�l���x4�Z��<�*w��阾,��Σ��>�3H�|_TX��rL����棟�euo^��#-{��x���I(�Cw�����m�)����p��5�WySJ�v�,�5��~�)}e��ֱ�@�j.���?XE�MM����������^���k�1<#k���2A�<��i[�Sӈ;M��Գ"&	��Y��~(��]̕'���J}�p9�3��Q"�6�X*�!V�����fi����%��P�` ݟ\��Ӕ�g�ּ98<�qc䴁ħ�xxI�AAx�dKN���y38�×�D���(��)G20��s{�vy5��8O?;+�ޕͦ�s��� 1G���3��ף�B���:����x6�or�	�� $7n#������Oƒs���n�{h�ͣ��  ��6��YP*�n�V
�.�b�XJ�پ̨��ޫ��kG�	� m!ĉ=3'У�ʰ��A<CP���3��n�՜3Tn�1��0�5����X�¸)�mqKtBn�$��Ѵ]� z�P{�=�[�:96�K�_;H�|�?���橽ĽY8��7Q"�]v�������n���us�öo9c�;�䗾��Vdа�wh偼���{�"i�|)�Je����Heqg,��}[�����8�5Z�+^b.��wJ�y��>Hw=?WZ�Q-?/!	�Q���*�	t$WX����{�i#1���#����VC�����TPz� �M�� :���e�<O.�Њ�]�pSnX��8ƘZ��a�k.��:�/���ӭ����w�����P��ز���w^�Ky���p�0kɔkLX��ݪT6A!�1��!�t��G��α��-�:�]1�xN+e��
���2�;��a�N���~��z�m���n�CE��m�	�I�]�Nh��F�1N���yi$�0�#/HM3C�!n2"Y��8�+����(�G���GK2�� �O�@�����A6#�HNR�t��x!��)
��1*�e�8k(J��?vY'~.����jO�2�PA��f_󌗺���#���t��	A�O[m��є:p�"E��5U4�-���kc7/��M.��=�1@��P�������&ˌ3J���7=u��.
JS�zQ�qk�5!O[m!F�X�Y�̩���
�!J�FJr=���M���ʻ�/�jV�Q�e��
��\Z������i�V�7��)e4�&�8W�O�S�<l����͇�"��d��R8+��}F���ˁ�/9щ"�{O}�Zگ}�U�f:F�\�Xc�.@���f7F���|˞K��kٻ����_˩[�:�I�T��H�w`��;K+W��@�̥����ZH������Pt~GA����m��1��{\L&I��;ct�Q�����Bx���$����,o��͒T%"jAr�+V��NV���N3�N��-�@OO��6`V��7Y떘N=�Ы���0 2�}B?��Q�rbų�+\�#��D#��K��J)�� ��7"�M�6����bh�̆ej�-tr1��*��i��O��UP�y|�q
���d�S@�]F�<�2�m�����0��Xg�W�T�w��.W(�
�E{M���<���@[��l5�&�8�MHkE������֓�ņ®�{���|�cЃ�!Q�y�:����5��*��k��@�dBR�dBz�"�Y�EΌfms��q1s:��d�d�Y����r��72�?_|z�᥵�a��n�f=�����Z�p�Ē��^����>+��I^�>u�6��!�D8��2��^S2�x�0�7�����R{���/�4V���T��Y+�����K|'Ƽ;��ypc�#'�;U ޝkSl�l�Kc���
�šK}�
�ʒ�� �~��� �+S.�B|�������DT���$*4V@P�,{^@6<�Mrl6tF�'UL7�9�%��D���CӍYg_�A���ۥ,mKx��3� |l,$��3:U^1��f
���w��@�t��p�!w����qe�9
o���(M�o̐a�囉W��҄(K�TƸ���c;�EzC�� �u<��ȶ&R������N�;�"[�t#E[z�=B��C��v��쏺r1@��hIl�w�wUM�:.�WT�Ԣ��FĹ�&��T�+�y�4V�]�6����#%��>���"�~���ר�1����$�ʮ����"�/�ކ����t�H�q�t�@4.0�ܰ�B�T�<2��	��}+�d�K�Vq�i�U��L2®f!�49A]g��[(�d[�G!0f~�����k�}�b���Rx6�SZp���Is�p
�#�P��<������Ń�_a���Uo�"|�����e�J�%c�k���<���#��>�S�����/�ک{^Ԃ�l�y�D��n�w��9�"�m:@����Y�%ܨ_쁗B���C����N4�&�����x���?N�lJ!3�K"
���6����͒i�_��VFd��6�v��
� �S8���Ɗ��-��2Y5�)���c���U�7�
,=Q�@��p��j��U�:��$Q��I�L�;6u�Z`*�M��sQ���&�|�^�������
�B~�Qط�6�uqB"0��[8m䳢��/�k��k�� ͛�î�g�;����l�d]��N��n�Ƿ	?J�,�,�筵�����	z�1Wm�b�>H�.8�TZ��/�گ��������̊~�\�Q �_�Ԝ��Lu�b�d�e��6���g�Hn�|h�Lꀽ:җ���y�tjb�N&�Һx�D,�VDan|�%��R qp��A#�P�Iϡ������v���,��gsg7�ʄT�F�"s��PP�	Q�"!���$9�G��DD8T*���	2�nֻ��>�V� ф*��$���;N7DSj���������>+�Fg���Xfܢ�W���(�$�>ʆ�s�d����#��8���IE��X\g��_ޜ)s��r����{�B�ҹ$����>��z�RMC�r��T�����PE�;8���)����p"�WiVO(E籯- �n�I�!+�}�ܷ��ʠX�;��c1ry�s��Mbt�f���c��>�a�Y�?�?��5'��#}`7�Gp���D�qr"�8wb���>��o#�r|�7�t��B�'6��TX.|�Ī���ߖF��Imߣ Ɂ����]�<�ik����?��=X�4bP}���u�[%Ěŕ���y}�_�������0r �Ӳ����c�쁽��e�.��[�\��CF#,)X���� �}_*�xZC��^�܎l"����돁Jγq�A��k�dn_r����"�>)9$b��Ng��yw����sx`��%s��?z���b|����%�QK����;�7tV�e#G|T$@`��dQ4j�����4��,����u��^��䃖$���֛)��t)�'��C�M��"I-�w��W�2���y����1�m��Q6d��:��s2'�Qe�(����t�!K������۽Ņ�&�%B8`�SI�s�_r���B�:�e�kRut����Niqw��K�e�JJ�Y��1�Ӡ}l���tr�� �T���a�5�a�co�F��(__��>�ơ	����/nfձ����Q��G���VK���.�,U��7�T�<��~��.¨͊��p��$�͟e�Z�7��x�10��|��+!������=��=�>�|4���#TK7��t�{;�8�[Ȼ�V4��BA���F��
� �iϬ����(,���]CYG�B�z�ӢĜ�8�X?R��j��^j���,��]Hھz��ܐɷ���ԏ��=f���	�����IF�@[��*B?�[��z��7o��{~���v�a�\�VF⟶8m0��*��e�߳��{�Ik�����]�iY�o]N���N���Lsu�f��o� ��J�	w3W1����Ca�^D��8�v7��%�c@ّ�@+�%�#+
��11��D��:�P�n~�0�v>�b�`���D��.?a���9Z��熯�MC�~8n2�D}�ܲsGv=f#�٨P��/3d~�{{|1����ߎ���v����8ރ��Zs�!��.�;/�/�.�-I�.kN�X��%�bK	C����i[��H �a�N���,kX���?�$H�t�}Q�a��p��g��4�<$FSu_=7ϔTkd��N`�A;Ȳ�E�c�==*``�1�l�Ї銲�?�.�p��BgK��	�p��Ԛ��5W��D7�j�D�H=��������#��shr�>s�}U���L��B��^[�1G��Rp�!5CK���j,��j���^$�n/�s����e�vU���c�/�Ez?��u�4��U��E��_����ڹ+����������UN�yl^�A�-ǟ�v����J��M����n.��fџ����=�Κ�g�����|��3��"{�~J�;����UhE��n|�P���b5=8��tF�]V�l�����D:N�� (�}���Chz4{��y�$� $I��O�`�g����[I�,��I��:p"u�p�?S̶qr��q�£�tK�ͫc����ĠwX����p���,0�5���R()Ͳ��l��/������y���j�y��E'O.��u}7ۯ�|�i�������^�����Rt0�3�̍�# '��Ъ�c}H9�>���9\����� ��V���+eoW7�=ri��nk̰�!!� ��ͻسt-/0"A�窰҇���
Q�M�U���� ���
{|���f���ɂ�0�R�I��}*=}ܞ�y2����Tv1��K^[��[:�>`�9J����LR�K��t��S_Ob��#pe���_͙��� �TS��b*�,j�:2��1��s���eČ�Ьʱ:���k$EG�D��5���c��~Ϙ�� �cO�&<bQ���B<�[��6W:E�ͅ���762�@A>7X'��_Đ�eT�zG
ǆH}�Ҏ���7��XS��m�]؀�Bσ�X3 3�U74��[L�q�������{��qI�s�uN
p�%��Y��Q�S�.���z�"(C(?��b�$�4v)a�Ä���D6�R� ���9�ǧk�^�1w ������0���0�x��*�����XM����s%�G����.�����?U��I��Xq��h�+��0ԁv�"ǝ:rG0[��c�v{��>K���S_��a�`���m���ʹe4^�Z'�g���wi��z�h��^@��/�~�^{��Q`NR�G(VMFO,f�!:Zc�,H]e��=r�4ͅ�;���-d!��0.���N�/S�t.5���~>���Ç��c�BsUS��9��Ȕ�v�!���\"��v҄�'v���fyW6���]��Y�T��.쫺6��zEh���ٙ���$���XB'`�19�����=Eer�k'�	�!@����V�r��gd�+58�Evq���l����e��v��ν���쑮�n{�+��{@�<Q$0��>oa.��6G��ᴱ��I��6o��kY������*�����E�]ݍ��k/DQy�ȥ����3 ƅ�>�<�у�NT@����9����&-�FY$���\1�mk���λE�W�q���h�B�@�`Y�L�D[Z&({��=�(���lF�G@*4�p{`�������E+�"�G�h��N�u��q�R��r7)���c��S�@m��P�FX�zu�l6^k�2-nW��|ء� O2�6�ea��\oo	�>��)��/�c����K�����ie3!�q�u�Y.����t�j�_ aIp��x���-��g����Ml-�=n⏗�y~ C��n��N:��y[��[.����C����g��>��π��"(5?��>���p�弯��QG �*id
�G��1�����	�P D���XK~�]� 1�~���S�����?��)8����D�t�r����f����=��°"r|������Z�?��_�����gp�䧴�����i5c�'�.�u�AG8iǨ�2�@�P��U��j�����u΂u&��?arʉ�����3���� d͊�JV=
�?�r����a�u���YC��;��{�p2�TX�J�C�'#d�{���:��.��9�4L��炐�_ٷ�؍��1q	d�����s�r�g;k���hu�.��D�2[� ��"ķ�eg?�=Qث��]� �s"a�ɉ�g��Ǆn�t��t���:�33��Tf��o�m+f�6X��;H��)a�����ڑ�r�H�n�b�Y����ݕk]({�,��T�wq����H�)3�����̾0���7:�E�P�@��g3�WJ��vA����M�S��������{8�TۋP7Vrkv�ͫ[�\��U�� ; � < +�X��{:�d��@k�C��g�N��~2��.�q�iF�,��)�ï`f�z��+�ɼR�<��ȶ3�H)��"�Pii�>��x��N��c�#�ѓ��ge;�`Q=��ǰ�U5�����Ym���{�u��`��!-�k3��[;�xU���J"��G{�0�����*E�,p�|R���t1g�����(���_4͍����}jY?�l]��tB�n�4#_��#ˊdQ��_.k�H�X#Q��ƭ�LZXO�<�A�o�{M9��e����:���������xZ	[Ԥ�P��CK��1�vV�r\�8X8��ck��GN�ݑ�tgfj&����� y��S��P�YUX ���b��~�h�/=2V����5s�(ә��A����%�����id~yy�
p6�.ќ��V��P%�;ϔ����iU��G���C�	���渿��\U�u����Wp&�9��_[�.3�� Ş�l��@c�*��$�1�~�Sߏ,�58L�=�݁�K�jS��M6	����;er���9�QT�1��D��4�|���.9��C3�>}�RX�ꄥCUa���*,�gҤ1C��ގ�jm	����\�^V�ˋ��s?5L,�3�IT�������w,�6��������`�~�K�;v�~=V���7�OeO��>�X�D������,��U�'S�bF��a~�.�iUH�~B9o���n������.T��>�-��2<���RHG�k��d������lj�9b�'��ӛ�O)���>��Z�����iF�j�?��s�e�DF�bSSh{z� �1���)rż;Zۄ���QܱF^�P��-�A�
2�p]z/�/��bv��A�9�|N5@+%m&���)���%�4���
�����;m��w������>ّ�C��2�!�47��ԣ^�����>s6iP����mdbmcrd@�Ms%W�?��^Y#�nL�V
7Q��j� �N��X�0惭=��E���Z���(�����Վ�s(	�Q�:��=��L+.�����d���2�o9\�@��;ϭ�_�sy��`�Moق�-��f�[�h<�<P�=Θ2֖������P�:0X�SI�Bd�OSy�qqز��k�$������Qrd�=�WĘ����K���Is?��U�x{����6ۺP�K\�� �A/�s��
�d�2�G�p�(���0fqf�a_����g*!�6�B@��S�p�O_{3�1�b��*в��2$��"���.���g��,Ũ�8YP�7����	�J#!��b�/|}G6ֶڿ���������Mr*.��T4��*�+_��.��FhI�R2���4���Ϛ���D[b-Z62Gt��G����q��n��S	82l�B�1	�U��E9�i��W
�����3��.M���#�i�Ⱦ��B\��If� E��%��ѿ�2@��&.�I�<�mp�oÂ��zz��,V�4�V�8.Gko��j0u�����06wGI�`�< ��˹?�1�^�,	˫<`|�Ջ�w����<��������8L
���X��gV|w]��Ͼ��@`��(�
,%'8ڹ�ʆ����rmrDm)�:)�����6NE�j��7����������UW��K�A�a� �ޮ|:[M_���Tm���B����6d ⡶����a@'t�Ը/�\�_�*Q������l�3BU�o�9����;�g��l�0�L�`q�.��������BCX���T1ޥ��+���,����!3�ePRi��������ӏ)��0�K�)E�G4�Оbe$��T��``�c�*����J�?�<�鱲��=OG�<���U�I�D�ϘG����z\�5j@&3>�%
%Y|}�N�H0�_���$���`'�h_�.zt(�xLX�z}�����i������J��������<R�N�*"ӫ��LO��%������#Y�Kv�	Ij��aM�¨�y��e��3	&��V����*@a2C��C&��-^.t]v����36�8�9>!���O7�DL��x�#���iO�5���������B�o�����$�7�o����^uʻs}�?��B-�I{� �u4:T~��WA���L�G�� ��q��<�A���2��4�9L�r����(0�5����zC��Ō�����eg�&�4�Q��25���9_HEP�����J���rEK�������v`��(6�Ëp�hg��?��'Y'�ݫ��fXN����I�AܺJ7Is�ɛ蚘L�B�/��G�i��eRk�"�{�s�\�Q��ic���1��3��0���>� ��R�3�� ��/���t��R�l�w�� G-_,0�!�4*'E.��^Y|��`��%��A8pu��+ϟ���=��*	xԴ���	Z�W>�m��0�t
���n��z� �y����?kQ���1�N���IU�Tu���7mΪ�ҙ�:�^޾����6��5�y�<��	k��ߪS�$2o{�.W.h�� 	��`cwrw��>���v�o��D�'g���'3��B�ޭ��̈́�r����v���>�E�ȬN#��T��}�W��zTHf:��2�h�,:�}��)������@B����ַl뵵=��e"����^[Ǡ��;�iQ�8�X��{Xo�^�����1C��GakLV�cQ�U�zR�_�4K��5��>�;��Q� ��{
NQ,l�7C�~�����kC27w��N���`�&C4��*�p/Cd�a��6K�����*U�7z���%����ςj�'A��m2MF��zp��ܭ�O�8.�hs�B�W�K!Tp����Ȱ�����T�xc��b�I6at+�ةo���qk���f�d+��k:8�t��ϙx���PL0L�@�Xd[ѼuER�w\W����얊���u�/E��E�(U���D�;��x�7�%~atu7��Ӿ,K$�e���Tn"�O#ŜݞX����pz�s����6H�*r�r�Kzl�c�Lͅ	W,]�Y���"z>���_f��m�+�g�����6�z��FN��%c�a"�n������ӧ%H�l��#��k��gȈ���գ�� K���1�����h���؊Y�,r�R}�P	������M1�4e���O��6����MM����k��e�W�Do��� g�[~���qs�}�o��9�!��n���>����FU�uF��K���$��}jy��6 w��j�\*ppH�`�����$�X��7��� 4z�
G޵���٤𧓔��^�D�.P�T��,�F�X�cX�/�0 ���@�iִ~\�!z��,TWw��zS�ǯ�n���IYo�d���~+����Լ�wd���Bʄ�`����8��HJ��|�0��+ݕ���wV�Mȓi���A���t1AE5���y-�2#չ7i�֜�x�V��>b�������L��7��1OEt[�\��lv��=���]��}���;a�<����nUYp�((c���3#�`E�Ks�x�X(����]��>WG~$SF���.pS��ͼ�eg��N�8Phso�����m]fX!3|"�r���%�Y�$���q��h�#~XH����e�?�514�{wҼ��}�n��7��1Pj��t��ݧ�1��VQMb&xy�*г��(O�Ԗ�T�lM2�����Cx�U"c�gw��B*��=�%5d��"����Px�T�m7���$��'��#�߁,S�A�I�B�)%�j�utI�S��"�Χ@8x&��~�LO�Z*E�ƿ �r�*]�M�?
�JW�?:��q���J��oYl��� ����VG$j�Q���1x"��'�^�Z����R�]�Ht�6����Ć�;�L�B!1C��0��| �ı�sm�̈j��"f�� ��8���uk�rY	(ʚ<4�)�R�V�[��K�����/����>��v�r��M�AI����tBS��NX���tn'a�]�vU���Z�q�J�ۨL��3n��)jytO�� S��Z����,��5SL�Ǻ��n�j��&����)�&B��O0k8YĲ��8����	�!:e~������C�r��k%���Tҁ�^aL���P5�v��?��-�@���N4��8�mN�߭�S�2�j��~���d�m��@�Y�{���d�2@aNץRk�� [(G�q�V~>Mi:
�GD�o�#+��Ѱ�����z`����+��~�o���H[��x՟Q�n?.����9�4_2����\7�jĔ��=E�����Y(��sRuu�m�*�G
~�澆����L[؋�3�~�h���/X��?]7a�[_ă8Me�g����r=��Q�n;H����b�s:����Ejw�|�]��4fG����W�������cÏ�E�� p{�\�#��|��r�@y�|6ސ=�6[�|O�t�cW�P��@A��8u����z�j�\Ǩb�D��!��|�tg���ei��'㿟~e~F~-P��u,��5�qx��[�\��1�A8�,���Ʌ3�@¡����W� �u-�&`O(��9������e�Rh]�o5�g��T�I/���V_r/��E3��j���lN��2%��x\��P!cI���]�7�Ha }��d� �ߴj�����҃�P�P�@lO}�#��A��6��J6UŉH���zEV�$�jL�?�k�ܒ����S�(���9y������H=��,#c�N�%����-{�JL�#�V]5���F�wm,���.=��W�A^�&/� �Kԡ������Vq ��=L%���SЮ��o̫����������N?f*�'2��҂|�ּ�?+�d��*��+�����;+]�ǩ2��S)vr�*d���|{m�z.uT�[��h�#�`YJAE���d���e����Q]K�-+�X�?T�ZkH˳^ֶxo������qf6vٌ�\G4I��vU�@ɼ�f��U΃f���Wș�a�!�`mK0��� !\�������?���x[h	.;/c�͕�7�?1Ox2@�
�m��yg���Wߋ}^��b���f��,��L����*	Gv�`�})�=���p�
�������{>�E\So�h�''��� ��(+�v?�-#����S��<�z�C�\_B�j�"u���Wy�a�.��@����/����?���u���F�xʖQ:�U�u�s^��S������E�gδ���ݴ'NVĝ��Z�d��S�K�2�D��si8����诹	�k���8��T�uyB/���җ8r&�
B��_c��@���(�>�Q������đ-��g��cU���Ń[���2��}H��A4�9ʟ/��=�,����j��!ۉ� 8�g��(��$�;���㬜&�J"QzS�լt;�OI1�p��l�k�j��yG���H��.������K�ūFk%���*>U�f�:�����T���cn�@k��蓋hR��,{��aN����:���p�_aH�$TO��R�n�H������(}q�p!��N!2����y��eʒk���M��գ9D�]rr�(A�lJuM���8�d~�����o ��>W\��賮�R�
�>����:f?�E�E���(���B`�5�oզlL=TdQ�)�],�g��o1*�F��(�졏�Q֋?�-B�/t�w��yQ!$5�f�@����������]1i��&��g�	�Ԉ\�'�0��̲�<����s=��((Y�,�X��Ё���tJ.��i��L��rw�s�qk⟡��i���
���M������/�\"B��`�� @�ڝ�K�*tF$q\�pV6sZDq�d�?ڬ�|�����`7��
��ɋ5"
Ż�[2U- �#J�_��&%�Sܡ�n��A"�Q�!nߣ��=#�K`�ˉ�p2<j���D>@Y�p4Ծw��f������渲�9O>��C���
�@��ݬ]�;�&��?�����9.�{5V�/ ��͔9��:�Q���9�Z��0n*�ϑf2�3�?��B4�@�Vƕ�7U>�i�f{����
\��㢟3�I��|�-۞Q5���R���,'���F�*O�Ym���GB���;�A#���h.����$ܙ/t���
�e����ss�߂i�.����tؠ�����f/�u��o�~	cΓ����k��R���F�)�?_�!ަ�t����>�1�u9繨^H}��jg��D<��F�7�?�R��mYp�D��ϋ�u,�|��0E@ܕ%a�����o��yt�b�����?�}/^w�\�"�L®��(��Wߖ��}!��#^��U�71ڪd��(�݇[Z��E;LNp3k���n��s3��-x��#�~!@���:�L�遤�뫣�łĭ{e;�4SϗF�ճ�t+f�F^
)�P���&2�Jq:<	��J>�WۣW(��S~���v�S�ŨOj\U�E8�0s]��3T�}���0�~Ol�5�>J��y��y�����~+vV��x�K��g\��@��W%�e�ىco����}:�/��q_C��]#���5ݕ���aF!���s!�b���~�$Ģ5�^*�c�����UH��1����8��gY��g#}�5�}�5�
=
ː*��%�`��h�v��{�%�@f��d���ҷ(*S-��o�!����2>N���b�od�*Q���-��_)�P��k4�[@��n��:� (�|*�-:�1�"��A�(�L^/�E���t꽪gahC��D��~�[�Ӱ{���a$��OY�]�A�%ε9DG�_�x�J�=>A,�:ٕJ^U3��|h2�����L���v$���M�T>=r&�������*���d��a�v�`8����!ޢ�E��ƞA�Qtm�~�������L��t%�I�%�E��ɒ��z�%��i����S�$N@�i����C}��Q��^-J{�$N�4n���`�<ߣuFb	�_��ڃ��G�8�ӡؔ3��m\��u<�sS�B�H�Q���|��6:D�O��p�ba�t������e����G{́�Q�*�W����P���~��ӓ��9�ά���}�VA�B��<}�[=g>��,�<��Zn��4H��3�Y��ɴ���ĥ#U�`��&F��2{4�6o�{���uC>�s��u���/2�Jz�\>Au�.����/bC�+��MՒ�̄�HA�n+IV��tb2���B2�8}�� �(�J�`(�d��S�%Ko����F2�"լH�
X���J�^-l��ޡm)3�̊R�\LN8g~��I�y��'X��+l�dޟ`S��|� bJ�=���3�i3��^_�F^Ә?��D�@�UTY�����ح�9���TSb�1��Q��
].zݬ;��2�%����/>m��Vӑ
قώ1�6����qO�����T�q�/�r�4hR+nK�X��c���X�'٬r� z�ä����P]hi���]�$�0���#+���~,��A������GpG�	�ب�n�<F�z���t��]�j���0I�y>}nH�9��Ik��=�'a�Hg�DI��m���������5���<�%�x�t��t��Fg���	d�Y�O��gu�-
�|Gh�nf��M:!�T��l���@�`U�Q��p�����t\����l�TI�i6��������&����7x�x��m���@�
�őy����߭�w�/���x��>��b�Ǵ�#=�W��"�Y{'�۶	$z���/:h6�fT���(�{ʫ@�41��R�ZS6ӌ������%RX��+��_��9��O7�F������S��|08��	�K�^�l�>|�B?-:8��{��O[`�	�{�� 6y}��׌m<$�p�ո�n?�^S���:�����V��$������R����YH����ru��Mv�Z]XO���w�o�a�����U˳�����x\��D!z5ׂ�ɶg��D�H�"�<�2Nk�M����M��G	`1V�[��IR���ڟ��}�?P�=��Ԑ�v�V���:e�T�
~�L��]���g͆�T`��Ϯ�����݆�Tm/�*̱��Nr���*$����w��o�l�P�����˜�	�kv�}1�%��y��!������m�{^�R�5�4A�w����X�k�p�����N��O���6>|�mr03~�G.oQF�V|��U�MXz�_B��'u�;����;ª =(b�h�.�%��A�9��r<�����w�?V����ڥ��ܿz@���.��3C���Ԁ��������G����kTS�M�4�70���9�NYS�S(ɰ[�
�W�j2N������1�����|$��(>ƈ�m�z=����d�fV��
��X9���$�&Zԡ&�hI���0��Pb�g�2��o
6Yr�>�.�gK_y���҄ 㮼�8粤5a'�0m|r��-v��ZƧ)�[�1��).���#L��,�Ġ���P��`�p>�C�H���O~F�LXpbg�����,���x�cgd��,åk�N2ُͯ����A�b�+�䡦,䲘m����H� ����^a�G�����K��p��ca0r���Kb�`�-v1�b��7)c��>�)�E0�E�Y��V������[�=D���/���|��`WH���c���n�����r��?{�D��E�\3v%<������]ԷnnRt�
�q8�#S*��{�,8w���8ѱ$��{��>�m�;��&U2!E��F�ϱ	7oN����B�)������Ǉ]�v�U�/��
����`�w��`6��{�_"^�c���o݆��u8�W#�P��,n���<�f3��;V��]��������@�z?;a"���2[������"+p++p9Ã�	��!o���l��L���$�b�6��2�,	TW�K���$pmv�V�x��ks$T�H����I3�w?cd���]�T�n%�5p�ЌK���*mħ�zf�|b��3-h����YRR�?SC����+22�v�Ή�hKP�vŞ7+$7�N^k�A�ؽ�e�F�B4�D��L�����A��.�ڛW������EѸ)�tfO�Y5����z�>����k����X�eL�ɝ������jߗ��U��MX+�����6����{l�0�	J;��'�%��r�r�������L��Tċe��B�~�X��=Z��ry4����Ʈ��&M���(Ç�+�P\;�?��M���`>4�#�m�},>�����&�-#�d=��68�V "���z�y��D�X�(�Y�Էv��7c������C��YA�ǘ^ݤ�9O�ȵrr�>�N�{
��ȣ��y�*"���ɝ���ҡ(�(�����<�b�9�����c����"��������}F�wd�G����آ՛A��8]�5�-<ˍbج;{4R������s?l�ˤ2��
�`�V?��F$��[*���j,����6� ݆R��9^�Io6l�C
��EC��o	��5��U���{+�"�/N�+(Т�+O��P�h-L���Dz&mYں�9f<��_��7����x)h�������OZ �Z���9z�q�3%f}�a����-�i|��R�u��w}���Փ���p7��z�ڝ�]Ԣ�̆B�v�]H���;p�n��Pmx���Jpr������l6�{��:��%�ц�a�����o7�q|�M������~#�9�������3�f�o��nDk�9��|�6eO���^�	�>�G�-�ᔔ�~�i-�K�`�0Z"��J�&�.�l����*��]Z>/�!$���"wr�a���9Չe�.���w��h�#,�e�c���]�^i8���5��{i�c������n�.�X�O\l�x� ����Uٸ�wq�Q�P��*//� wE�D�YWF���f��c>՚��Ǩ��i5)��F�t$�.���bdD����K��H�yH�=1�[�2�,�V�;�׼e�(�D��;��k�j|��)���HS�3ڒ��;_dxԽG���Ɩ
>ߟY�%?	v�`��<퀇�b���ݷ�lC����p�"�+Z����)��^7�!�@����!���&}% �����Ϥvm(U��<���r}_���������>�W��A ZB=�}�ڈ���a�j��h��ӹv}	�U���� �K�V�6� �`�]��\y�Z�"w]lo�!uG�lOp�t?�C�����0+�4A8X�8���O<���{�F���������$p����(s��r����Ϝ�����Z��$lWy�X��hn�?��t�G�������v���|.��`�G���ݷ��gahe0��/l����Hb������BƔeo��;�L����7�g~���m&���{��oJEd�p��G�7��_�&���Y
P���*�z��G	,��MR����n��ꐇ�l�(9��~�HTa���2���{�UH
�8�N�0���>}��R�(����m�.�ÆЖ�k^��d��yG� �uH���k�!�m���6+�1�8���/�DO��h;{��j]C,33`������ϐ��
���o�V[�՗��
>j^��*Mب����ٖ/�V�t��\R�c\̞|}��2�A=�JJAjh���a����F��'zx�Π&���#Z�o��P�~
����(A��V�������1G���?���p
�>��y�̯۹@=?��4Vi�!���9۽)ōZ���.�Ö�V��}�i���<��s�\�jaȑ��*�Q�����Z�_�B��w�!��p"܁���Z�A��"m&)�W��٨��<��$��(��̝5���VAm�$�$�Pi$W�����q����,��xS�=s 3ϸ�ҥ�=�8��A%���3�� �= \�sQ���9J��e���H[˳���pg��`Ƴ�v�t!�|/���E+��'�@�+j��Z�j
�����%��!k�:�#�	�Īӳ|ވ�:EyIuYa�g=m�t�;WK�0���-��L�(\��e
'_�r�%�J�-�Fe<�l�Jj������a$~`��Ȼ#A�{E�������^���̥�vS���5K
����W�ƛ�o{��4�b�Py��Hbc�H^��^c��93?5�^D:I���s��s��h�:���eY�حtam��x��\ȏsH�T6eZ�j�ª��M6�2;5_����_�ѥ韤�^��/���v�������`G3�������鞀�����h'�HF9�:�a�����'��M���:2mS���2��ٟ*�5�>�2Lq�UL��y��g������z�1��!q��@q���:��Ԡq�bm���3����^ƿ�z�������LUMKp�����V֋I T�]��E_pdx3���nLF��d0�G�	�Cc���ם��;)�ˮ3�9,��&���a�,<LZ>O,�=oE���
���H�3�����U�%��	�M�ہ��)��b"�a��@NB��D�zh`�k�a�$�1��­ů�h�\�C(�dM�����"#�/:˨�o�ޖJ/�y��c2�V��0��B׋NrA����/�ir�y�?A�S_�{�ܢ��ϩ�=���2��F�Z��q i;��6L�k@�P�f�.u�r(�(<����,~�1SW���S��Nݻ�)5C��ۛ�U[&��I�bt���z�)s?�09��Ŵ�Cx���ge�jY��7=ʣ+�ҝV�G�nz�Y�,|:fsjf�Q�~ԗ`�Ę�cKj���I1yRa�<ܗ�נ;W1��������{2K�{ ���NA^e��S�����h��|� ��%�B=M܎�j��d�N�3΃��6�|�w�L��.I/��M�gչ}뷣<�cȎ3�Se-�2#z��6���,y(3[���qG&� �|��L���d�a�!C���{?�!y;`z#��JpG���b���t���{t�kh��5�ؘ�aJ�I������Ϳ=U&P���w#�?�������?P�&���z��:����Lr�%�|"D2�����M��7����%���@|-��j0
~я0��H���%�#�u��C-��	i{b;�@k�|�zZӘ��O)}ES�k��L��.{�v�fb8��C�"�`�lU�O���t�p*�.=u���$��
��Y���o7���iX�c�}���BI"�]�8���8�9��s3���kx�1���ᑍ��m���21}8L���0��Ҏ�*�>����I�co,���	��h��Y��$^Lz?Wii&M	����n e-������N�#$�1�x����T�h�2��a�[7�L��e��H�S��q�>I�6uA�'lB�yB��[�$�
:\�Δ*.��܍�����em�G�=�5����G`����ȿ�q��v��;g���C���8��W��BW��Է��u6fe��#�:�`i�ǋ��������q���V'��1��j^�dM��='ۚ.>\t�ǱuN����B�Y+��p��y�O����"x�њ!��|c]$������Y�n9ш ��2��D�?��n d�V9	bJ�wkZIb�:��OM�%�R��������҅�+t`#�1|���vID�9���42�,1�� �y*W� B��!.Jn �� �'C�]`gd��.Ң��EO�ǞDr�A�m�2�N\����V���%!+)�⾴�u�:��:��c�,I�"��!���(8�IaR����cu;1 �\������?&��uϽ�2�C��t@ ����n4���l_�0oc����Y�� ���fD�e��H��0�����y)�� t���Jg(�Cɳ*P���X��!E�v��� ��x�Ƿ�9����t�f��-����h�a�^6��oU�Ԇ��T�?�h�9���yʚ�a������4B��'UgPd���nd:L�7��a�=+��P�ঢ়�	
V��b���rψmt��|d����L�303��ʙ.GUw7f'y�=쑿�׎�1��A�NmY���ш���r4ff� (��!�l�j��C`��#ӛ \�1j��N�A���?��׽,
����3h����{zԘg��� E�߻
c��B�N��B����m�a�nG)���G���Jw��9�}%n��I����O�'��O�����M��gX0�ú��&����z�����������V��l�Щ��
�x���b���o�2�5E���G��e}b��H6x�<����Jӳ�Y���$�M;�@[�0Z�[9O��cc��ɘE�/ٞ����T���Ė�e,�������KI�������Ć�I��#<�sZ��_��,`����h��[;Q3^)0���o�����k���J.��-l��JZJ�E�\�uI�]�7`K�
�G'�C�'{�7m7��t��[(��)_���4�Q�j�,��8d����/Yr�hލ�E��Ӣ�F��$��-1U���0���<��(��%�ܼB����ՑC�2ꖬuΝ?�F�Nu�|�_�o]�b��2��h"�W�����rl�sj`V��4$� Դ�f�On���C���JK��g�3�io�T�E�ܓ���ȝ���[�{��7-�;�����!QBg��)J�4���'��6�x���j
.`Ȕh��9�z�;�r��V*��C���EzAwVHt~΍��#��� ��|��X!k�d.%K:	�8v��iG�?����r<����oE��n"�ؒ�eR0����dTF�s
T�>�|_��,x����JKB~�u��$�H��=epH�`Ҿ��Xr'E�z�@��W q�P|�`o#'b���)�oGm�����u�;w���6�����`r�(�g����cmb��¸�g��2ZFl~#���M��	��榹6!y���T:H��k�*`�![�Va�?����d�*��f�.B�q�[x]IA`�f�p�jlߗ�W��i͵>��̎"'�hK��s/]R4KG+w���c���a�I#�, c����7�$oZ�:���������
[~:���HS/�P^b~ԭ��9X���0�wLe�øMk��}Y�I�w�n�#��oj��^�k_���7)^`uJč�
N��j6hھ�XQ������- �;�*�����7���n�6�&����iy2O/q�	~��O��/�P�A�i�ҹ��d�"�+��cPOy]J��A%�d!�tf�s"q��2��������Ok��c���Ƚ�T)���M��>��|AD
�#���~4� �~([V�EC�N���K�_�0ij{|g��5]J��k]%����t{�����0>1�ݟ��yj��\�o�M�.1��+գ���[�2Mq���~]��k �}|`r��@�K�V��EQ��nbY�~�Z��)yL��lp�V1�!j�%�In�)x4G4}P8� ����+܋AІt�	ёP�8�\`rce�WM
�����^m��h�Z�Ԑ���%�<�2uԿ�4s!bf��.��UѼO���,!;�g�7(�j�WF�B��6�Ҟ#��Ŕ���Z���6�����X��*}C�c1�/������C�\��-��
����L�,�B�2��� ���_�pO4�>�<��'8�Ѣz�$eN�[���:��7��Op�*��Q���ؑ����V���-ԕ�<ZM�jH��^g 枅����f;7�Ne`:h��yȰ���n�)�9��Q%5dgZ/�Gs�4k�2������̖XCF�rǢ��ىq�L�}V�g�=8TXF��w���x0�)�-oҴ�&�W�Z\����I�@����3����*�~a�]
}�CJjj�vjV�jG����3�������i�Ih<s~�޽{�R�D�"Z��[���p����ertx�D�� ��:H�T���G��F�o���y��)^N�ި��;3f��ٜ���H�`��a77��T����¼R�G攏��ֶ,a�K��.4��g���K-�>��q���B��#f	��L��R�݁��XϰǠ�g��ll���,c����y@A�3�D��
N�esS�2����3:������zp̫w	aZw����@��n�d����{����}#�9>܁��A�a�FH�+�3�Z�L5(<鞵�.���p����e�!�r��9E�6���K�������N��y<�,[������ED�S�Ac�nn��*2�W~�Q�E0������J]0i�W�C�����m�����|�*�&y�U�v��qr(�=�^!���o��A�������U�j(�\V(��a&
�]7����W�|��Cu ֚Ji��(���O%����6���xl�����ĉ��M�Zn6�b�frʮa�O20��UA��� ��v���R�.=kI�pm��T��EÁ��I�����K��7��GO�+�P�9�՟F�Zu�)�+(���b�.ڋ"憨��ު�C����4-�_	�J�8{�M���2]������Ć!���[+ߘ���Cn�l�U�=������ o[�H� *ŸH����dr�άB���B����+t��#T����M�� 1r��Z8�G]G�D��:֏}�H� ��7��+�P�����o@_!o�T������X-��+kx��k� ���߅�o��Z��! /Ht��s���1`��
��	N��j�Эb$>]V)��l�� ��.L���6��:�$A� ��D��'�n��z��"��Q�k7
Ty�8;6&�P�nD�]i@+n-�xD��m�Wy�y�r��7^g:G�J�I�-�3˽���&�vCa'��)�R�fí� ��9و6,[���ݓyȔ�c�Uco�A��\Z��N[Y�g},�gJ�����['Jn~o�!	��p�*_�ڇ�Yj�]JJ
O���W�Ic�d�-�)��(:������̄�v��$�٢�^ Jt���.�¶�z���t�ӗ��ٓ?�G�!R i�L�=��T�欿�5���?�0�$i�$z�ZQm�6�9~e'&f�<-�[�x�؁��CW����So�ˍ);��ث׆�b�f�`�F�h�����x��ȍ5!e�U
�x�5�[�����gV�n ��FtP"�lz�>�V�zPj�}�6+��X����gH�U�E��qM��#�"�ٛ�1!�H�y��p�@O(���� k�&b�.���P�`m6ԕ��ͺ���:D.�C�M ���`��t�����f�aS�)�O�c�V�����;�+Gde�Z�6j��`!���������v=��D�f_�Hbq��nv6���Zd�wiĆ @�^�}��­Û.-CW])
�@{����)]F��=�v�a��������!��kn�[�a-�U���L��fnNN�G@�n�=�L��R�wiG��n{-����0��7|n��$��6���xbY]8�-_>n�m�.�
\]O�`�~g�r��I\5zDZm
�#�_�9V�(��Ő����%\}�/f�h4^����T	'%mu T���ЅGK��l��J���%V�A�`��v�l�-e�lT�"��̗O�rAU�ДF��$�feݶ\�B�F�]Fy�%�h�M!x[���M�`J��aw��$�`⇴˿�O=z���f	D�NӁn��21�00"��ޤ���ic�A�������Z'6�;��aE�|n��ʎy����5��f���*\74�X��p�x��:�z�)�r&�3�_2W��j��΂G�Qb�7D
4[�P�o��W��_�o(0�	ܰ*����5�꼮�v*k��)PI��Kf�$5���ۃ��Yk%���$�ϱ���1��Ѳ���*I���xzH�8B!�!ţu��}�;��3=#��EgoZ����Ţ���T�?����$�h�!��N8��1�$��+��h��_;ch�U��kӬ��zH���M:��K�������^ůb���{_��ܞN�w7�#�g&4��a��S��E��M�UJ��,8/��m�Y����Jij3��8G�1�{�q� *ꁁy.A�A��Q�*;��L���������Y�)ӿF lk!3/�QBz�
��<��7֔�l��!W��_�;�,�1lp�ۃ��]ͨf��ޝ�;���-g�I�����E�\�3��?=�:{��0���RM�n��3����V�gV?��r���?�^N�)6{M>�G�AC#����D�K����EP�"��r�!��:�/���$)S1�{�|�x���P xyL!|'O�* "��xSU� /H6���n4�8e�D�ٌ�6�a�G?�#;4���*f\N�v�����	����,?{bk����sc�ľH�!�:Œ�D/H7	N�*b�������E��T rg�_�hqoy�������c T�T�5�㣻��g*��\R4I�v��(]g[�|_ 7�S�s\��YR�i���2}�6;��d�qƂA����a�-�$#����虘�PE9�'̫mWڜ��dsB��4���BqߑjmL��n��2�n*K����w��$M���y9 ��WB^��Evn��Z����MfWV>O ˛�?�̸���J:z��4�&<��bPd��lyTg,d�d �Q�6���u��"�>����i`��l2�YW�ϕf�,�\΢҂�\��T����l����6E�siFv�����.NK��<��$*��nv�4�T��*����:�?|�fȿmQ�j�N$y9eY���3~����'��\G��!�Z+~L�L}�2܃�_���,(�N]=Zu�A˛�r�4}�լO���.mbݩP�޾���n����$]r��%"=��(1�w�������P�fi�_!���?g�8-Fl%���%9�Ta)�r|G	*��4E�=����b=����|�#�_���;~/ņE�9|�141��b9�5*Y�1�w0tr	̰�A�؝�����F�7'6���0��^����̖vf�=)�2(]̏a]]�0����;�$Wi��I�	����(`;���
�j}��!O2
Ȋ�������ܻ�Ťdp� �]�6y�T���ێ��ͨ�� ���9G����E�ӈ5W;oH���l9ǎ�׹~yrDv�PwT�>��d�3�ˆ�U��%$�+�f蒎-��yV��7�X�JJ��G �Iɠ;�t&?�KQ1&)G�3���'OE��)۸^8���O]��5P�w�ν��P�C�&)a���/�pk����V����$�!+��^���C��U�����K���?%k�c��.Y ��f9���SyV�|�U8<lĹ ?z���kb:G�]!I�����~z;���7��c�`޿�})�{��I��6u��^�Qƾ�]&<��e��DU��o	U�NI��U��P�rX�1N����76n��O���t?4��v.n�;��(f .9R��墌������DUjn�'@}9��*Uh����i*2ƣ��[��}�����䪤�jDU�����p�^����[��ä��89l���W|��
w�E�X�~�M|��H���RVx�w��`͒�ʢ7�ry	�X>�ta�W,o����G&��U\�Bړ�g`,�����aIJ��ʹW�ɉ��fO�`X�9�����t��;�K�l7��&��/g��x ��aX���jm]TH\�Pz��`����؆���QE߻��{�k)��P�Y(fF�_u�Q���9���<������y�CC�.H{P�<V�7W����.c����q�=w"��,�׀ڳ����`�W���S$�^VQ��%��3���0M����`!~�4��ҙ���8�	/}*`�{�g��K��V������O���R�ϴO����3���k �4zMot�<�?8�ht��E��>�:U��t@�}3�4�}���C�h�3�+�.4�~�q��oX�"������hnr�_���Q ���JT�m��5D����*[Q�F��D
�%�E&H��xAD���ZԮH��@C5� ϴ�w��02��;�p1P�h6��!kK�E��>��j=vOw��$��<�@G�TGs��ث~Z+"ws���j����}(+2��*����	�{�="H����Ҷ��}�f�����u�]��K�a��'��HNG���v�H���[#k��GGZ���	(�,}�X�L]}���
��G-�����`A�#at�g���_��$�ܡ`��j|�>VIS�B�7R؃%BLr�,<j
�0\Dc"��P
��jA?�� ��n_���HK���M��[]f�>+u��	����R��x��F4DD���������dV�]�L�62$aN������D��Տ�;+�}� .c~�<�N�l7@d�<��7mz�"�ꊑ��ˣ�������ʛۑ�+�W
h���?��1�s>�x�����v��yC-��r=�~.ǭ�đ�krFyj����ּf^��r|�5ey�טof@?��7rs|�}_d! ���S���(�OUBhG˭�
�^1.�.�X��[v��ee^/xl0lh��%wN߯�ǋ�`J�l�%uw������c9�Z(+3lb��G9��k�A+n�Tg���22��4�yY��~S�\2\����i��	ڕJg59P�:�0��d��`��F��m�|kUH.er�I�Pm��)��Dљ��5����*��_�K��8a �P��fZ"Ў/�?�JM���2�k��.��2�I���S4S���|�K�l�Jͩ��Jc���L<ge.�[i���j���dU���d�!1��[���z ��G9i?���JN)�X3P�*��U7q� '`S��9M݊��3P�����NN3�;X�ˉ8���/�{b�����@5�fYͮ��kH��E-8(S��[��P�<5{ۢ�N�c��V����߰k�h�98�vP&���`d�� }��3�ԗn��I\�8�0B"%��W���*4�@X�B8es"�.<���º��R��t�]،�W�/�rN=A�|�6X�n�B0�ؓbf�^ʢ�q�]��=��dN@M��Zq���<.
}
��{;=[�u�Y[�w�+u�ya�X������jf��0	<�H�m�gh1:��	љW�=`��T���PFR7�������FYz����pu:\��4�>r+�4_�}��3T�⣊��^i���N�-]��Uo&��ng���e��:��X^3f�N�$�$c��7�
� ��Vz�7�������C4��������
͊��$c�	 ���@:X�>�Ss�Н���\�n��Y#g������tT�vv, f���Xj�|�%ӃZc2���Hqͫ����>d|�pZ��5�fH��}y�#h'��2�� 3�SV�ze���)����e�R8�/�OS�����'{ ��Vo�EI,�|�Øpm��;d��ұ�~C�`�o6"�q<U�{��ڊT����Å^ki��n���g�����_^֥F�(V�J��PaDڦ�&���$U3�K3�4��t����+x���PH�PT)�LՊ�3E�m?�E<���T7_"$��єI��)��e���'�����[��g�1��`y$Z��3�^Ua:�X����D߯�`������.kgw��$nL����A��@G����a��`�M���<&.�٪�]&LL;��Z:(������L����a*P�n���S���e�d�(����E�g�r�+Eܵ��vt��w���.��S,�ŹPT��aP�j[���"+��2o"�S4y\U,����.��v�����ڐ���N��#��-���|��{�Y��󶳆���|�J&͖Lݸ��~��� �n!u��U��L�KIU��] ~;KMQ�8p
D�8��ţ�������&K�'���f$��.����KhJ=����Eov�f<���!2�`C���XijHƖQB`y%�C��J��*z�Y����s�#����G56�Jo R����$�i)�Y�6�[�?�8��|-�j��R���//�-ǁ��\��h)(&"��X��l@�^?nQ1�>w�hl>p����/p�q� '���)�e��Xz�8��D�P���֓��9c��I�qH��$9�of��1|��F�#� {�E5�M	p��f}�B���W�(t�Z*�q� Eƹ(7�����_nY�#7
��FiW�F=�=�v+�5~f�P�唯on��j+�-���-�F`'X>XM�E���*t'���4�;.	�t�I��n=j�V*��T�y-v�7Dn�f���'�OoKǎ*U鷸Mac�cU�M��H9(�E76�o���7L�c5Σ��yD7@ۄߩPa�Ŭ�w�b5����SÃ���TzI�E�&r�#�O.~� J��h0�Aq"�(2��A���-��� �l��o�u�L�ai:�-,̲�`�(��Al�ԕ4V��&�ʥ5�5Ƒ�ۍ p'�'��M�,?���ƷtT��.-5(H�|�NY4^O��@����!O>��k%�o�� Ԟ�	�|F'�A�rqmN���'�g��ZQ�S	u�m��py�iI����ꈤ��Aaa E��~�@�TT�F�dѷ�<5�Ȏ(H�mĪ����^OO�j��������]���Չ�^JOg�}3�[�@	a:�TP��J�2e��C�I  ��uS���]�qu�+�W�Zv���)�0y���H��e�y�awk��$�<��X_1n���Дv�����݋�A;φ0s��Om������&�D�{�U�Ud� �
��I-o+��^� ��(g�i�il�����,��B��Q=h`%��fqH_/��6��p|�84%r��K�(q��#�/$:�g��w�s^��M4z��8��",EéΈ������fˬ�y�a9��Y�QJuk��S�K6}Cw�/�V%w��8�Ne���_l��pD�2z����ۜaE	@��$p��u�n�3,Z����H[��]���^g3�6�=�Ѣ���^�̿�����E0�AB�Q%���3��f�Ha�/e�o�������v\mU$�Ȯ��$P�m�*�������^�޵CV�����(TINxخD�
�}/��m ^&N~�d"n*���
B�EC�t�+A������i;PM�LO�Oˊ������}hS*' �V�s[~���}�,��!F@�g��6��Ϛ�x����R?y�|�����g�eJ0�i$�X)��/��QpT[�RɗC{G)X��U[X��T~B��ײ�M~@��C�k�����;H�f����Qy�գ�U�<l��*/���^����;^ X���&(�F�9ܴN0��_��a���.�(L0���S�A%�$���BM`����K����%�Ejhw� �g�.�qC2��>,�w���x��L[� �W-�D�lǛ�J<��c!�B˕;�әc�)b�i�;�w@�LZ��3��=�@M�A��َ.���T'p��Em�t\�{�(�������m)�ɳ6�t��ND�c�R�7{�
�����\21}�6�l��td�]_�Ќ6,x�r�~�@g�-LU&��Bu�o��7��<1%�v���UNo�*\Lz\RU��c��hK���7���7�د^m�]/~[�WI[���Ce�8Ȼ@�Ь�w�m�G�Z/�mSŤ�¦�S:�hr/�����'�c��k�����^'Ȳ�� N"�ݮ��·o��$5�f��V�V$o�N]nS��=�* w>�7ᢎiJ.�� ~��7��:�Z��>o�x����5�si�0*pj)�8]�'�g��>m�{x+�=�w9#���g���q�t=|ȿh>l���\��n^z�����)L�����\A�>	�)Ki���U�^�Wo��;�$D�\-��tb��@>��Rrq���Yߠ��/�PW2�!6������oR%K@^�=3P� 5���UTS�+�,o%,nS�q]���0L���ÖP�������d�ln�+v�X畆vϼ2�y��?(�����]�$8Ac�'g���ƩP'L�ӫ�hC��-L$�0�D�9�Y���xjj��pƔ
�u$�O g��Cl>��J��Ln�>�7���a���x]*�[*O/�D�1W~���2a�hf�j����	�>��ĳT�s����Jku��0X�ofE���!��茔����ab'�b�@�Kߕ2����ȴ�:���$bH2��Ef��P�o��_AE�*�	���MI� �h�Ƀ��Wh��k����b����dj���7�] dE����/A�~��,F�`�Ä�'Э�d�	9\9�#��.�yp�˘ϟ�Ҳ�+�opSd �����D�.O�ݚ��5�
�q�$_@�4&$��&i#˾v|�ҋ�f��W�`�fR�j������X�?����iI�y��lJ��dH �e+
h��P��C(�ǿ!#ܛܳ5o/�,M�ސu���|x������xS�`�:�B�;���'ؤ�>o8�t�uf�\���@��{�݆2��utĂU=#$$���<����k��蝣,�H� =f�v�.ժx:qW�!��7�����*S���'c�KG*�B�T�O���?�l��AJBp7��������5���k?����幜��FfPďP��>'���^}�:n���/6v\>iswՆ
�O���P�`��tM�m,9�<�烷:Q���=X|Y�z4A#:/v5�����yKRfr���{����,��X���ps��F��Z���lIB$�։/�ȧ�#Fo����E�o�6{�Z�j�mM�����H��?j��h�?l���Kf�\�&��;Y$��>��=Mڛ�j���(�Ym�V��)��`l��_�� l;��dʦ�3��*���W�N�!j� �ۭ��a}����͘��zH�,+�Ƀ�����s��.V15�;����V��rkPf��Ŕ3�2��8/�w!��s�ޜ�_b��p�1����.ji��`��g�h�� ��#�Ԇ�3�Tf3*g�HM��2�t~���v��r�b	 WK�_>��"S���^�� ���a,���{���Q�1@�1��m�0h�Q��ylD�[�#6�^M%�6��^�2�u78A<�M%)g0�/���	���Q��'�ibg*+�u�g&ym���n+�ި7�A��D(�z��G�Z��$��/��x��Q�A�4�=�%�	�kS�d��L ���<��^aH׆g%�<�4�m!�PS%�>�k������(%G�[��Lk��iW��%�1�R|#f�_��^��#�c��0��KV�G�5��^�Ҭ֊��$��Zߎf����z/�a�9e&� ����że��7��!���n)\:�?�T1~�S�9	���_�Qe�Y���
)����_AHކ>ȺT+�d"�V	���L�f4���\�Iͭ���q��Fu:ׂ/wًǊ��Г��.6[u<g2�j�|�]Q8r��1�?@����KIm��3���ݼ�p�e�B��(U��(ݪ�*u�*���Y!�e���|��[k݈I;��d�ꉁ��d�?��^����~�0�����D:����.0\�"���X��Z�� �ވO���b�0�(>(T�W.�v�0	�L�X�]G�MM���g�{KI�� �ދ?j��@n�1��dw���M��[��%,�Q.�tҩt�y�`� UK�s-1���rP��ȏ�� Y)7S[5UEXӕ�����dTo�gT���β������z��w{��*�e�]�%�0 BB�E��0���_~|�[�\:�~�Z�Y���*<�WC��%]
�/����A���5dU�1N�+�G:��w蝗7	8s���+ϥ/3&���>��������}��}Y���bU��Fu�'�"l2����Lδ�8*k��5r)eT����<�b"\��t��Ɏ�������jj`H:��]�2$��6)wi+K]�w)gl�/VӨ��a>�*϶�=]2Ҙ���<k�!w�f��NsX	k�t�c�"fx�!�JX��+2X d{:ż�DG�W�u-K,����$>砼�<�rwأMbCB�3�ފ��g^ �1��>����ZJ��1�|�`�*�?6�O��`��wd�A���B �U���|T�!~��iC�ĶϾj�r��JH:������V��Ʀ�sJ$!Z�{��\���AI㧜��2�e��{��Tgb=�QHhM��m�i�Ӝb�����w(e�T�iO1,�4��ɖ�~�ަ��5�k�C=���aT�� 5�q�{\3Ea���Թ�d)v)�h��t�>��0��,�&ɽ�&?���b�-�!zX-�h�����e���N��O����?i���9N�X�O�&OV������֨�
\���(�*�����%��?�l>�q��.��idy�]M�}�pv;�Yn��K�c�ֲʖ�Sg#.)�����_�t����'L�"�0��r�G�-�F�Bz	�8�b|����\Z��������o/��1�L�ՓL�a����W�� I�zbO穃�Zm���%'�ު�k��������$��|��¸�ž�r.���|�Ԫ�t�a���K!�,�z�ک�3 d��\�O>Ȝ=)7�&\�_����M�֚�~(D	��킊��ݨq���4Wx;�D��m����~�.&��N!1����Fd�������ĝ��a��:@q��F�	??��Ȓ�P��*ffsZ����A�P��h�5�c��1T�0�^��X��k{�̬��`j�CvU]�� /,0#4�`w'��nQ^��P�y���,S�p��Z��g��;�����ϊ�� E��c+�0ɓ�j��Z�)�����.Z����a�/���K
A H��N�7�����޳��e��Ֆ����
d�Ѣ��ǔ��Ãh��S�TdS�uehoLJ�G��%(]yM�f t���#��s;{�H�����xy�s*�H�����FS�Ҹ�ؕ,���|3J:���Ӭ�[��q��xC�
����8x���蝢��F����a\#�͠f	wwq��^��c�nj�`P#�M����
{wk]xI�6�(%�-�g@Β��X�M��w��W�qy�T2����;K���/-����֑��� �����| ����oe���{�@��,�M�U}gv�v��Y�x�$���y|L^P)��yB�b�M�8.���Uj$�(pD[��:&��o�^Y���a��40�O���
�����*3���7�nEd��c�d�v���'�r�"N�ɑ���l]ɉw��vc�w��y�m4X���������h	��"0�4�h�$��.�!}�Љ�ƉgL�#	b� �'�po��ݡ�S���	1M�5KU�9TX�"�8��@ 0ņ�*�8�l(���D�Ľ6?����)�ϰ�pr�ܤN�W���3�a�ey<����=,�����"�?�'Mi̝/��{J�?������:x������%'�FMPf|�e!�=��G���m�< �����b���Mm�C��7��1~���u�v�8�c}�*���y9 &˔���y%/Di�_L-�[��^㊟��?�4��2��"�O�R|� ����ݯ�]�w tR�K��ސ�LB��a��\�;�*��e��O���]��C��iz�͉k��z��&�3�| ��)ɫ�ɭ������M-�%P��J��ҍ�ӌS�<��:��/����;�vR!��k}�F]L��������$@�żw��풐���P���F�br>�0'����}v�U���T���P�����1�HAS���
h	��%��3����-]'�}V+��C"����sl�5z,~TԿX��Np�i�M�l�^������@�HY����T8��@�࢓�Ռ�}��Х�Y��K�B!�?��~��9j(4.eT�6*A7���#�4xǁ]N�֯�����Z�qmK�"cŅe��*HY�N��ErAe�g��%�F����@Z��m@.os��yi�@���ۯ��²[:bGIIL)p?�E���=����2i�8��	�+���׋��<&�
?��j�B���:��Z��"�k>�/���ǆ�fC�Գx  �aZ�jl�����! ��b��g��0e-�QÊ����:���Z�
m�	zP$�X�ߨ0c	�/7zg�Έa�S?����~M���&�d�v怒̣�ت<hD���x�}a+��hR�Kk�r�e�@��8j�9v�|�����4W�ŏl�HDH֑�����|���{��A�3NE��F�$��rс�� �v�.�	.��?�|a_`.��'O�K]��a^>�@{��[&>t.o�o��}"��F�#/��}�aӬ<$Q �0�rr�L ���5�\V����Z*L���>����S	�{̦�;v�m�XH���V�"��j�T+	�+�-E��W�0��z
�c��g�<�@�zh*��I�K�g�
XnIK�����4r��b����P^����E ��`/-D�UKvld!?��G�+v@V �����{H}����Q$���]�ίKA����Ut9�pq��Ͽ�0��7 �'E��\���y���c��o+�t���1��eV�a΃ʧG���;���"J]I�ˬ�����?r�D�yQ�!!xBh��rM�Ё��������&3�UȢnK�)�&�$ryQY̎;E��	��+�F���yK�"ɲ���߾��p�8(h1��Op̳�C����%�d��i��� q�W��b�
Ǯ�Vt�+pe*B��+Ap���A��߉��:�����>�-S�o3�Y=��黗w�ha"-�����H4����iCbWD��Hji,9*�p��:Vd?�w��d��N��Y�Qw�[�ʸ��뫐M����2N@~D좥Ƿ"$Tx٫��|���+WS��i��gWK���-\�?=�^�	���E"���׹0�K�l���fc^/t�~/�����%�hTRԾ�a�nr��:�ږ�I	��+3��(F�2w	�@o����tJ٩�ZѪP���7�3~{�E>P��g��VZ]n����|[�K?)���h\ʶ�<5V}���Ĳ�l�TwU� ���~��:�Z�3��W�g�:��.]
K�yK�"��|�Q3����&�踠 ����Y� �W+��y���F�t��.�㻐S����i�����f���A\}D�F�G���I����w3�d'$6 �s�?Q�VD�0:��Ř tׇ�� z�}L�~᧴FA[�W�tZ+�G�S�O�h��ơ)��{J�"���Z������*��h>� m�O
� ڭ.��Th;X�F?v�Jj0� �L�Ι��C3�U*���6����<�TH���>�ܹ� &5�1N�Ȇ�p:�p����E�f\��rzZ�ș�ܑaą�8Q�,�3��!�I�E�I�� ��w�L9@�[�̕|��ΪR���)J�}K���4�w<e�2C떷��="؊f����x
�md���N����(��}O�+��@+��GP����+LA��[~����*p�M�J_o�^���M�m��/r��<�*D��%�Ղ�7�A�a��4���4���&e��a��sv�S��@gZ�p<���dR�<b��Z�a���5ո���#כ�[*ò�5�BHC-bS��٪p��m�;���?C���95����(��o��Ǹw����W������
7s��::.�0�}Pt�!)�Udq˾ף�q�in2-}οW�vT�^Tbf�5�9��nU���9��*+:@1����Dݜ�7��*+�b��I(��7a�p�^*.]��
~J3�zf�ǊD�ӻץ���M�ݞ�)����O.�N��J�k���c,�0i�p��TǳU�����ʟ0{�rB�PF������H���ES�(���8F�l̕�pS�����|E@�IPn��W'סk��`���Me�7؀%�w��\~!ь
���z��.���ɹc3yh&��Q�@��u�LZ�G�6bE�#��gfŴ��<@"����:�����T+��i�ck0�����w���9(���=���á�d:A�'�i�:�+"Շ�>�9"Q"M7|u0~�y�\����m껕qu�L7�~�>�Ǫ��5��xoL�H{�G�;��? ����T(6�5d�W�IT�"M���4qu�QqH�Rx5�1�`�Ɠ�*�g� ���Ne~�ʾ�p:ߎ�.�m��wcG��!!��L�nl"v1|
(�`|�P�QedQ�R��m��[C�f�K��@@�k��1ڎ���i0;"�(g81! ^{��L������G�@ߨ@�]���/����Զ=B&��=���R��B�;��MȤ��z�/� �Qh��ؾ����Ο%\o���49hd�J̷9;���qoP1�uNgD��S�w�-��`�4��ۡӕ�y��K�"�=$��C�ݟ�|8�B�� ��=*��/�gB*�K��JM��r~��q����TC��]�*&�(�y�/��,��8�)��T�m�a� ��eɶ��(��O/B]V�e6\|`L�<�<.�RA <���P����SL�>o'b��5��_D:�St �.��ʝ(u���-b	�n'B�х����>��"�G��y�;��c���92�@���=_b� [Nt8��)J?�~6�jp "<�4�/�-`;�	f!���1��x�"Ov�t�o��+�	�k��f��H'�ⱢR�Qb'S�w��{wSsUL�����j$C��Nlܗf ���ø�K^i�d�3/�㒅C6�����wi
X`|��_�;�q���?�>ו�,����u�'T4B��}����~�(�۫w�H����C��)�ϛ�_��c��T�5D���[�;��B*"����`���:=(+��P�*���CQ���X�g��<�n*jԽN�KZ>��cN2�KP��`AT����dA����6�� Y� 5����_Ԉ�v�!�x��0/��R��L�Ӗ\�L�^rղ|{p.*��������[�f��ہ��7i%�.lY�~��3⥶�C��דéD�@u1��
��B9��P*��������i>u=��������^���i�L����5�ʡ��a6��7?���j#�7������f��1Wr�����}�}W���&]�E`���/�7��5�$hG$:lW �j�	*����~߻Ό�!&�qC7�~�*p4����}s�ͳ�ᘹc��ɰ@)��B���	��Z���3���e��y}��c���[	��HF?���	�k��S���v����-��S�;�l43��H�-�^&�,ڙ��X��I����5
3ɦ/إ �����&�����1M�S$�)%i#�38:	�~��9~2�v��ST>�yNe�e n��ɥ�~�kU
���h�BlK��O��ygqZ����������y\�YwB� k����Z�N�6)^���s|��2/��(�^Wd�<]�^}���.��#�UYnf���u# b��H�gﳧ��|Ϊ�%��,W��"x�$k�ܦ܈钍���+ O\o�U��8G�rXv	
�;��ca=;�8�n~4�
T�[�Ftn��o뭊��g��|��ʳG�F�%-+D��fa�����
V�Y�2ǁ�$��!>x��8B(�5����뇓S�V�{��A���<J����9w-C��{K��6�
�7eo'a��CZT�PI�hGW1+�7 �	A·���Z&(�h�����T�{f�l.+�2�1{I��5	Ν�ß�����s���U�H*␼Q~��Ylc�sFO���4:u�v`�����N˚t������cx������vo&zMz��6��+-��~�<1���E/0�M��hx�VL��WRf�j�(z_�ΐ�3�A�0�U�S��P��a��,~oW��\�V���O�;�J���7�J��=�&�M_X�\ޜrc����T,moE1��J�C�Yc�y����	Š�:Ҁ���S�$;������"mY+<�jcj�И���.@g�|O� f��u�io\Ͼ̢/=�,�^���G���m
쌝�mm�~���E�@�GD������}��(-���_&l�λZM�MM��4gG�5Y��$	ݴ3|�ϯ����!+����u:����]��Gz���{��� �×���xE������]אYn�ږ�˦;���c�mBOi{:�D���c;���U�z�(w2����)Bk�[r�(!�Ah�N�V���ei�N�_�^	�;r,IS�ۮ��~��<�|��=`ϙ���jN��|��\��:��`e�R�e:hz|�cGT� v�L���Z�S'�����q�D�*�{Vj��}D>�&Bii䆢Q���й��b@P����!���1@ʤQ��"^�|�A��7֌$�L����0�j~�ɹRL����bgC?v/A�������EL;w�/jЀi�I�)Ʈ��y�U�_��� �[[������R��L��(g-Eq�fb��U�2�>q�r����x�Kwu��ض]��i������ �l��u����Ÿ$�ٌw�ϯ��a�Ud-K�?��6�
 �'��Id�q3�v"���-��
I�"��͛��������N��{+�JR?f	f��i�,�{��WgG%�,`n�,��t��ٿ(�H�W:3n����6�G$9�KE�R&��'�&��w�{}��7��;�VC��(�%�9�4V��<@�� �]׊�Eb�?��e�iItu�V�����swP�įF���[a�+��~":A��c���`ģҠ�t7E�7a��UZ,����jኘ�IB�m��C�.�J��"���)��@�J��5�"�߻�����~kL�J\&3��T�����M3TS�@oy��meG��zu!>�m�c�j��m	p�f\�ڂ�;7L�fǾ���nj�k�Ǽ�K��3�i#%b��`��PP�(N�#�c�7����f�J[��CM>|z5���c�=�P圄Ӧ(t1��fQWp�|�2-�A`j|�0��|$fGu�E,�j��(��6�j��;�㳟:��Ȅ�Q(,48v�]YL�ńv���n�U�wS���������P�2MnD(To1�b�Z���T	
d*�0����v��r��)�V;�kDs=��}����W�I؍�6�i�Rma������9���PUϾ@����$�y)rf��ݙ�N�#�(���x�խA�;K�#��ҧ��2U
şD���C6C��$�?�+��g�*IUN{JU`ڈ�	��&/2k����!���u�V����SՅ���D$�Β1�@��G�^����>$���훘,Zf�%0U~  O[3;��i�1
�#h-���"j�6�q�of�4���x�1��\�r]�\5A3��$���Z�Ѿx8��_X�K���H��k#���d��Sp#��f�������VF��%	7�b�W�,� �Ex�F���v���p��T�lH?�~��}#&皶(�D��^�o��8�͓�W5/�1b&�\Ee�4+A�7��Wh̑y�����
�WDjV�1���������5�ʊN�{�J�Qކ���vi�Z���K�~�L;0�����C��������w��y���Ŋ0�{j�KP�X�$+�ԣ�D~e�sDQ��G+�6⋪z~X��ɶ��֭�<�[�|��R�6⼐��@E����:��d�8���ޢ:!��R��0�gF�d�M�C��8�Ԏ�{=�� ��׾O:)O��{?�K�����|�aF{ !�-W�?��W7�-�/��р ��h�j.�*D�5ƌ��5����/x�Q���g\H`���xA��$H��n�=��m�.c�x���w�w�ڀ�ʍ���������	�vg������m�:��9:�a�&Ư��uwy^k���64A��`�����枽��w�,�Kt�ǽ��������9��֣1r_�1��a��lW�/f����cң�-�!H1��}�������T�}D��B�`H~1���)N�)�c��������Xc��<��\���h�J���ϛ� ���o>�����L@� ���~|,6�၂d;;�K0'O�l� �i%���"$=Ӫ�n��dǪ�?[�n����#K&����`4&6���ņ_tU����ѻoU<��[��+�"h�t�����͋�>�tXf�"N�.����}u�w��t%�y��&�BOl��=]�
�'��c�*TùW[���Am%Bgrb8�Ă�b�--=냴5�.<R��k���iO�:z��;L�Ԥ��XA��+ۄK�}j�38:��!�B`�	<�뮦5��$��	Sd�8+�����:���ܴv[/g����R��C֋�v��)�R�sf�R�VW�F<�?&{#�z��Vy1 �-��7S82��/�l@۰Q�ϭ�P'I��9ghمj�̊/΍,:�|R^}<�M��=����K�~<������A�6%u�dT�6iguVy�&.�z+~�@�\x�F�t����(
5�;`�{	����\M8�&ǳ}4t�Nǟ��5�!5�!�����'fo���+7�]��:�B��4u��t�����^���hg��1OG�7���JѨMvb��R/�:ߺ����!�Q���FѪ���%����
�^
%�ӧ��0�?�����W�4@c�ʨ�o��Cf�}nH'�VþO�
e�qss��b/���x�7��q}&`��?���+�Ƣ��+��G�%��At%6]��<B�(�C��˳�L]�i�j9�.)`�IƏ4�sz��m�r����ɱ�e�Ddt�e��y�8�4��o����K�p�u��\	�g̍]xVv���+O�΍r#�<�u?�
Ca�[���/V,���H�Eu>�/�P�eUZ ��&&���:\�8{��Od��F�Q�f��o�$����3	�8�J���Kj�n��u�c����k�V�ㅴq8Q~h��'MpD�L�ĉ���p�e`�0k��:X��7���
:(��������{��㮵a8��l��0<|��Ipl�&b\~�!�� �L#O�b�+u.�<��n��?�)�%�En/�7�P8,Ǻ<�-.R*Se����^�����H.p���6��n��;�U�f��(�8Ď�-}��f�Hk�L�J�Z�*v&�F��zh��<�A<�o�u:,hҺ#cY�C�]�R����mȽZ�`�Ԗ�b�?]���r��O�)�EX�/��u:;*C2ZKn�%U�d�ډ�~��r�:�5��m����LorQ���po��ڃ��
�s9��l����G�c��Hm|q� �AҮs���1v��}�/Bτ2e�-�?���*@�������A�S��_����f�/��wusu�*uWlr���ZbY4��U��1~�׊o�~{�qY$��*Z��^�x�@S�([�_�r�	�]��m�VM��,�umS|~ky{�P�\O��L^����:��aaג���O�il�
���྇��yk�X�Ө�}6�e�͔C���;�y���I���P�i�b���`*�#�
�Ƀ�.��!!A���w�h�86��4��`���u".�ڡ�\�b��?�ʏ��!��M���?�������SQ[΢�XbU�Z����L�b��b�j�O�-��P=E8��t�Z�4�n���{䃝c ���߲6�1s�����4��Ʀ��\P�C�g�JOH{�"+�T\w��FV�|�lڵ��������\Z�G�[�h~�c
����*��������k�<*RK������9Y��x�F����5�#����׌�'Ը�s(�"��� άp(��t��NsM,���*��iNc�;���4��Iv���.���(�V8 5	$���OP�N����ӉR�U���,q	q�e��d���3���3(��=ۖ9n`k2����4�H�qqN�(����r���7y��g��r���8�ƃ�m�!�_{����Y�b��h���f�=�A\�ӕ�u�42��Ҡ �B2���o��;��"�B��ø�5�/%H�G�N\����*�)�X1S���'�� �Da/<����ǌg�gg���Q1��Nm��~Z<��YEgW�����L���T41U��?����U3�>X�
�e�㚒f�j5�ʡ0�i�oŻ�e���Pl�d(�����~��c�1�>Jt�=�М	fH�7K�����4�ҫ����rϕa�gI�������i�}D���w�<l�C�˝��� {�@��|W;4������_;��+SN���	���󸆚�{�ӣ�����3���˖1�CV�`�~��>��B����FdR(��^���z^����Ԛ���c�o���^y��������,n{��D�[3&��{Ѓ{��uW���BQ6rV�R�AD|���I0�f�������I�	��9��ٜ���k�Nq&�cȼ��<��k�c��@��_;'Y(vI���닲�+�nd���	�!�=2m��3��A�<��~��z��� >+D�>k���v[�/���Ǻ� `���ǖ¼�S�z����.�rĴ�g�0C�������b����+L�Y\���Ӹ6N$P�l�/(�(�}�U?ʅe���j�S	»H:(Ñ�wd9��O�W�sn�\�pI� �;=:\LbA��L��Z�`�H4��v��ۿ�i�l�뒕��>��S�M�U8\Aϭ�W�? ��c�[�-��:�.�t���a��,�b����a���gQ���S�;"T>�����p����+��>�䉚oK�f�z`��|T���"\ӂJk��3�l/�A
J����C�H }	$���i��"�z�W#a�a�4�=�oL�"$DypSU��!@���%Ҵ�ܽi$�e�^�tPS�?�9V&�f]͐Ŭ.��[�l��sչǤ)�S������j�~m�m�S���s��?���@�	v�x A�4�}?���?�`[���cO�fkV����Ԩe����ό8����K�wG�sV4���LP$�E?�-�K�7n/%�������;.lxX��*�Э}t. ɳ�α�  f�T���yNo̞��qqcR[X �1\���V�� ��l2���B�?:o3�-��G��3h�?�3JL4��yǢ��f�fg���-i�$e2�Y�I�	���h�4���DHM�Û�r3:q�[=� �6��r<�^����G5�I�>>�+L�4�˂�9�Q�V�9Q]ac��ʦ���gw�A�Ҿ}����S�/��1TJ��gf��7����o�nQ>x��Z��S���.f�-{�\����].������ej���GO��k�y���f��+z蠑r�Xf �\�:������>�v|�A�]�?����
��o���J/J�����"�C�g�"�<���iG�����_���Nj$�ͮN�{-���>��`׹�w94(\��'��l�s�1|�KgO,�� �=�����:����SX�9f@�`�,X� �B�w~�������oВ4P◂��U���xԋ�r��|O$s�����wN��rU��}WyvF�v+�i?KZ��X`$]�����	� �qP��v�cL��e���*Mƭ��	�U~� Jjc
Ԫ_i�Ų�7Ҋ0G�/L�m3ݬ��S���qr�6��15B��V��Q7L�\|�VFۦ�{`!�L�ؑ�ښ���#��i��>
�=�����Og�����(G�fv>@�y����^���7����x=�@��/M�����[������e�R�`���_1(�Ի.�CT��e\MSp<��s�M�W�B��ǰ�?���r��[Zҥ�*���T�����A��,[�3��o�c�a�j��8_mڅ(���r�Q�*Ԍ��T�Ԧq2��A�_tuTkmo
!Ę���B1�{�%��j&g��쟠�9N�p�$��I��)�*/��>&�a�1�����Z��xS���޳
����w{�U�fy&鮍�Sg�ʊ����X�2�-�R���Zǫ��c<�Om���*��TÒ$uӗ�~9��ܾ��^��t��6�]Val��9!�NoJ������d�p)mt���"U�J������L��,ڈ�(	$��%���=�%�!w>D��r�9N ��ep��
�u�1�Ma����-��-��K�jt>���Vbi�})#�5��"2�.ȳy�幖"�8T���ɱдz\�{a�l�6x����h
V뉋73�"�d/�^9`*��X���bw��z<Q���S]��0,+A�8�%\3�C�T��7��h�_%R�^�ݵy�
���4����7���� W[���<�Om��=i�	�t��M�;���K}��є�O�� �pv�aG���ձx�Ol�<��xOJ���	���-#��Tw{'P�^�����2W�s��]�F�->�x�c�xM[�;���񋁐u5��aV�+1�n7`�:G8G��p�?�_�+J�_ ��d9����;��G}�r�S�sg�|pP�®�Gi+���ϑ�+$�i���\���8�D��V'�\��N4����Ĺ�kH�l�Liɨy))�eK�b�G�ͽWϺ�@j������w޳��O��O�5��`�2�@�s��q��&b���VM��埥l����¿���,X�Ps�.CW|$ҰJ*�+l5!�Y����Pܗ��*�n̟[5��T�+y����E`�Z�͵��WmM�luHg�JШ�5��x���-Λ��v��5��-���N'Dp���3��״�6���{ޖ��E�̕�b0�Mo{�Vj�hv��5�Gh>�z�.�oפ.H	�)�	�3<վ�ys�J�s)�D:I9����1�ƥ��]��]����12��$_d�<�j��34�j�愅s�	�u~$�X��}r���$�:,TOӝu�Su������o��@ ݀�Sv���n�<a̽��SZo��Zh��
�B�C	H�I��0zh�w!v����,	zP��؆(���Toh��,�̲bT�T�4�cO(�c}h�E!Y�NU�-`�C�$��q��Z���������,%�d<�=������F��>�0Ź�Wd�t�씱 ���i5.:���1��&��`ө��$�l�I��u���<�v��� ��S_4��)$Bx�{��Y�1�#�26�.���m��j9�a/���P�~f�1�]Ts?�	��a��u��劖`���C�f�[͏�Fͱ�o���cj�V=�?H�H��q[玹�g����Y��ۄ���F�������Tu� XC���$8ɿ�yl�S1D�~ۣ��.i�st|;f��*B�>lG����.�g���0X��F��h����sofև|�h&�#�.�����
5�˭u��wޱ5o$��N��ޮ�Y��=�V~�"��+��"o���*��k��$⏵U� ����BoQ��|/�7˪���麤P��"9���4�#]9b�R>�s��^V+]
�J������Z�o속/�:���"�s�U�6y�����u�	I�K�ASek�4U��,��@�'�m ��%C��O�Ͻ�|/#�'ۊ=������Ӳ�j��s��6�%�В�~iR��E��am��1%����9+d��ie7]�3�Q/$ � �e�=��?5]nJV� ~�'r�Y���)�-�kp�*r� ј��f���mDt>��l���GDZ����4;`�t�Lv�n�r!����]gi�O���l�s���=ו'�Q�=�=]2f�%x�6[�x��`QN��������=�3qœ<�z,��=��3%f��'/P=���l!j�V�_C쿷�w���rmHꆢ�g3��z�FC���2�vaHhgB�"�.]WN8�YG��y����PE���D�+��槐���ܯ��������ht�~�i��a��G���#��y�쇈挶�/�oJi�D��i9aE������1�5��}%o�-3��r���x7��1e��\��9�4�Q�"j ���Ϊ�����*�8��)'�RuېSI1���j���tN9��|����[�G�Beym�|�&��u���{�)x��$-Rb`�y�h]i���?Ezİ��1b.wo�@Q���M��!Y�k���m�Yp�����<rqݽg-ZG�F��[U��)͟ )���gb�򂂼�V̷����*W6��ԽS`��M�E�"#L<��Ԡ�S��U"_U`�����G���2vr8����� ��:I� ��T��z&�Q�!��V�k��LXEk9=�4o�=}��H���*g��ZV��Mض�O1jl�RBsq���F��?���d��vH��L�����c��Ʃ��V������,����Z��/W�Ƅvmݚ��+�l-e��l\M��t"T�/S�}���.{k�}��>�RsNN呄�v"I��?�ν�bT��0k���ۿ��R ԛ~�ddd�RT��cR4m����ۗI� Q �a/"*
N�����E�� Zq��<��ش�o�YC>%i��n�u�U椆-ӂ����+ЕT�B�[���F�^z��Y��qP���ژ�e��M�ɣ �O����d��Q�E8��i���U�?�1��$���GD��P�� ܨ��Ł���)ӭXyFb�rY�(� A��M��sW��E�J��&�A@�K�ɀ��:����e�-\j{�;X���=�Ox��^�`�h 	����=$B:�I��*�;�.uq��<�����Mv��L��\�,\降�^T�]d�P&vj�p\�o�ṿ3��l�k��R��q���/�m����c����!���(����;�[$ʋ��q�&>U.��o	����
�p˗@����zހO�l{5C�}�}��s9��Q�)�d�_�m)�AЖk���6��A�}�O�-�9go������ͥ����R��U�����]/���B:q2v>��[���� ���w�7�)�����<5l~�/5Jź,b�4��/|J�������=���t���3��-�>7�Yy]�����=8���m�J�v�������% ��3ˬ103�������l)�"����*=(k���,���'����4��@�=Zx���N�<X$���f[g���lށ�u~�:2�L�H#��vt$��sG���%�>W�G���'%��8�3z�`�f?q���˽|rJ�yhF��R��]���
u����t��K+��&��-�U��{uÑ�Q���:�޺�uk��.���B��t��:@KO6X�`ƹ0�t�>y]RBO j�՗�-����e �n����zs 3����fw� v7�^�+�m_I�K�u�=A�m΀�w�&[����`W��)��~T���D�H�6��ʅ���h�i��0z�S���DApdh��8s�SdO� G1\'%S~s`�C�'ӝ�Bp������6�����,�
�l��D�_!(̩!�h<0]�q����酱��H��~��Ow��/���i�		���g�|d#eorܺ�1�E�ڎ	7�+���D�$/�G��W��&�I��.u�J�θ���3��L��,�`8l�|?[e �E}FFT��U �J�tgb1F��2��]�l�������q[�3~�:N�Z>�v���EY����#�y��㹨�w�۹���6�!��W?�֞�
�24��m�����u�	ԇee��5�WPKp�ㅏGOl)mMNB}����}n^)%Jf�k��G�W��:�����Nw�sE�2(�`����%�m�?z�d�|:�vJ�v��f���y��4r(��~ جr���8[}�dz����x�c!�J�W7-�h����^S��F�l�*T;��y���R0��
 �eC)`]˺~5�e�p5�W���F!*�ʗW?�F1����dك�rYաZc'���4�.�pz�o�N��+u!Ձ�ǝ�/�+l߂��7g�]�*��2��#�R�#z��˔�h3��PP<�p_<�4��QS�>��@%��$��²S0�)���Z�>��Q�4`��g��@�),�`V��5U�Y?�8F��r��$�e'��4��e ��ن�}(ih��Um�N9�����y�K�l�|�����Z�j?\<����(��[���݃�<f�^���E,l��d�����dfW=L"��]�'L�+���hh�|J�*T�E���b�7�U�П�yf�9iX�l`x����aD�r�y���phy�w4!dv�G�X��� ����*t����u�����r�m���X�[�o��:#=La���ѧ@�oZ1����� W��q2�=\�.����5A�ɛ:���d��GL	����	�ҠE>�G�����?~�-���`8[C`����v�VP�)|�~ᗋs;V�ػ�Z�b�"}�G�����A�������+t؟�td曡�Ƹ�Տ�KPv��u!C�h�#�f���I�SkY��m�6DHr���ix���˞C�3%�-ݰ�
�c�89�Ge�p�AZ7��� �թA'�r�k��f�HR���0���z3�P��hީ��t�	�o�H�S%g�l��+O��Ƶ�S��e�7��.J�=�����`����j�t��Y�	֘X��NK�]�C�8�������h�Z�e��g�E���|nL��D<��ʫ�����r���Bd m$ }�ػ|�V�v�1^�9�?���Y�k�h��ڧ5�u�hA��1	�q�����Q�O��K�8�yl�+;ON)צ�y�0�lFjom�������l���
�=�=޵9S�f��+��V�|܎�*	���)���V8���N�� Wl�?~�p����|��,�V/B�Ɣ<�Nd�`0z) w�K�?.ܵ�!̱K	-��
�B����-d4���F���̪�Wa�2��0n;�6@��������e'Pyi����寬|%��iq�uڡtM����ы�m�>���Ʒ�����T>�m��]��7Ra�I�&��o��X{"nZ��k��[�l@���Sb�U�9�-��I��n4��e%��=4�c1�S�@���,5���:�T�q���?g�EK5�g��^�U0Hc6A�c�H58ܦ�)��`0�!�%�z���%�%��3?�eW3�	]e�i����"�BӤ�G�{#k��ak��ص����<kG�jiJ�� �s��
]ҫS��#1}*��\gS�]���r����+Ro(�}�BV
�k`�`k`GPǟ�9R.�A��jd�!�]AmU�|� H�՞CR��t<Ѳ��dVӟ>n��6��'?⩺��|e�B(����7z�.a�^�1��
ǊW�ӆٮm\b�ꖱO���/� #3�������=� 4aKȀz�,w�CT��2�!9v��,<8Ī��ςL��K��6��&���̬qfҥ#��X���F���/�$C��u��V3���2�0�\f�f����:kZ�N�c���������K����d���9JU7�Hc +y��_
�ԃ_�;ƹ�$nS�I�Z�X���c?K� W�'�S㓗ەC�mӒH��Q��s�1*T4JLT��a����h���_L��&�!#�^J��T�wQW	���uR����it-@Md� 	��
��!��g#���&��Z
ό耇�5A�`�L�B�fRq������� 5x?^n�e������fP����¬�MͶ<B�g2"��Y2Fp�a�p|6n>Ӑն\�/Y�Ɵ�~����U}�c�l�ړd�����=�LJ�����Bt
 n1	���'�+��8����?�8��^�ɬ���A��4��nP���0������]¢6��K�x�i���>�m����XOBq|r�Z7f����猙���]�s)�Gw��Af6�pǼ[�ፍy?I_��w������S����-m�U��I+�Ȇ�u�*��d�/1�����+��2���GQb������Ct̴���(=���>���勞@���lBs�kjK� ���i�ɨ{�g�UZVh��l.x5K�S��i�;r�R��C�Px8��b�k�qh���(��5����Z5��Z��g���kļ�4���0Gz"�'%:�n�#Bl"��݂����������$|�¿� ��A�{���!��w�̴�?�����a�WU�6���&��C��6�����S:���Zd΅s�!��U}\��	���J+w��y��T�#<�hy���Cr�#p*����@Zh���9�Vl)v<j"`����؉n3���>|�v�8�Uv7J!�d���^��O��k�xн����͉��(�pK=!坖?l��}�Lq�+Q|��` ��
��R��uڟBʹZn�$2\0 ?���#�چ��\8��_7�b��%�b��Ӑ���DT�w� P��nM���P";$Y��t�_�<������ ��*-�
�y�pQ�;t�X��ʉ�DFG��m��S�^p���'DaZ
ıِ��%�:$���j7P�v-z=L�4�uJSUp��cwN���Q���J���
�p�c:6��MK-�N�w̿����ݏ�x?q��(������^�.��j�珡(����R�X~C�_��ْNW+��"(��~��^�T��e[�?�t1 24�􂝕�P��o�Z�+��;]��0m]��ȑZ\���u%�mp- *4I��~GU�%?w�]��iq�Eʹ�}��|d�О��>CW���F��`�0��B:<>����G[��l��B��j�y��X̳Y���*Y��ԥ�H�� �Y(��E����F\R5vC�(�!�|�)`+��4j�b�kBH:%�X��A�A$��w������ ��b��H��r)�g�s��u�o"��Ԙ�Cp��/1�E}@�o�N��e�6uE���|[����R�F����@�;w��+ K_*�����?\�	����i��ǲ��p��̎�Qy.
��%D�Խ��O{`��V���B��m�d9� �k�������~�4b���Vs�%��)���>h6O�?,��g0L�RG}/��M���`�j~�f;�9����R�,/C��64�\,>Dտ�B�/KnSC�GC�����x���eYc�Z�� ���7om�뽮i�X�
�J�iC����;e����:���f�G\O�#�B�������/}�U*�֣����}�l�7d�,��C<�~��O��лc��[�}�.���p�5�w��z�|,,�����P�Ov�a@�����W��o��ĕÙh"�k��j˔�JP�Z]� 8e��E�e/���ƕR@nAH���q�
����47X��:KPk��އ9����e!*�s(�],�>(X*p	�63HJˇ�����䶟��l�S����la�Dyu�Hcv_�ﻕ��椡X�|��E�r�jt]7 `쀌�C��rp�ʓ�cF)�馒{]�2p��f7a��78�)?ݼ4�tiģ��0�֬ �[e�<�@M��|���H�I�X�D������z:�(��?���S�s�� "��f��b�X{���<�UN>���[G4Zʡ�UfQ���s���o[]�_|�*kz`�����ɹ�LC�^\�נ��Kx�C@ZK��uʬ3D=�����bh&��0_�r��:4��̟$�[".-AQ�Ү�QFDE{�2צ��Dx�v|kʍ"i/5���]R��W�p��`�`�%�,r��ш 6w��C��>86�PD�ʫMJ��i/X"W�F8f/G�����@��O�e���of+��5&O�Dh�����h)�Yf!��I�;�j���t#��>� �#���Ae��fN�������7���<q��Å���T�����.��S�Ħ�$�j;����Tģ�C����6�~��v�uu�_��'ix�?�y�P���]l��3�y�(���[M����3E�LӁ��O^0Q�Cf���7Y�H�������>�v)�-l�]h�?\dc~_�c7�	�Cƭcӥ˨��H�tɃi��Q6KP�5^Y����j�P�����@ײ�
U��M7k�g�t��D�u���.��O�ٕ�1y)Y����	K���s��>�i��Jo>@c����/B]�?`�h��M��9[3��E�LBY�V�ck2�9ΝA�>�В���u�U'��.tr�6�t� �0��=�ބ�
ֵc�
��I� {���qm&�J*��bU����3:G�ݼ����&C:��!X7����=�N���_xz�?�:�QU�^��7S����F��I����k�����f�Oe�Τ��:r��"�z���I�H�9����9��xjCHFTV��q)�B�1V2vʈ�Zy۵���L�eRTq���M��E<r5V��ثR��{��Ɲe`�A��-�[9bu�n
ہ�f��'ӕo��l�\�T2-҄B�3H���^���V'�<��գ�Xu�����A~~�ܰ�T9Sra�k��pj�UɀM,�z�S�E�$���]�;�ÓI�٪�\J6�[kHR$R`�G%<__�{��K�w8�\t�+��w||�V�|�b�!��H#�1樘����M�v�a�^-�6FM���)-H�3�{Mt���F�ͅI��$3v�<�mŝ�s�H�
�h����&`n��#����������hh�e���eN��t=[|���2�n��N��aH�T0�[�\K����I@�K��;��h0���y��)Fz�	�W�@)���;���y3��e��s)�ՏL�����tHr��<I]Yjѵ6�o�rմ�0WsCN�F0�Ӵ�B��⛝�p~LdL�F"hn�oY�u{�G/�,A��9?T�kd�%MJq�U3q���n_œ��*���d�l���-:Z�d��&y#=�u�H!g�1�w�K�>����JV��Nҝ,f�-^��"���E�M&�lu"�����
�
xH���+F��ש�6�P�VJ�!b,�XX~�4^��ꑏn��GJ��w����	�A�s���*i��.�����`O��WUnN�B�16�̀�w;χQfb�x��d���ׇ�qYs�k������hi�*OQ�R��r[�ћ����b��u�Wx�d��i�gD�?����R����$Fm���O����	'���'V�h+��\���D�ǺJx+�(cs��b�L �rW��j�b�W���^x~��Y�gW���Um�4��w)9Y�t*�z}�3�7���,dSE~����@~��Ғ�&�&H����-8Z
z�-�r��iB����f�|_�e�������q*��X�������4��������48Ipö���ѰN�����}d��jTz����~g���`�Fɠ�-���B�pR��+�� �?Q��$P�$
U]�<D�<��~k4<k�^y?TLQƱ�Hmp����F�İP���W�K�=~!���G�%t@At7���T^oK=��ⷽf�^�+�
�뛷=��<-1������{�2����:L�n=Y�^���O����n���8���gp�,���oSʝ5?�B+ ��k��k��ސ$b�����|_I�`q�Yײ����Gz��`+�H�.�� ƌU�R�^�]�R���P٢=�(��jLԵ���!������J�������]�m��
k^*��E�Q�X�יּk�:�?g^��u![�">�k�+�<��ݲ��w�쾑t5z��Yͯ���Z�B
%߽�p/3�a�8��[�i!�y����+Q�O�
p����@?lM/T����÷6���o��э�/���l��ֱC�WII��!�4	#��[�B�`�(j̹�&�)\-���윮���Kd����'��P������U����퓞�*H�1�g�@��o4�0)\2�_5h��=��noݐQOm�fz|A^[��MV���P�Q�ƩD�N^,�f��@����ܢ\F����"v�B�P/t����ȫi��E("*�:\`�E�8�Yo�T�I)��P�#d�#x�7�Bĥ��c6��z(�)ߗhu��s$6H�y-L�Q�Qx����m�5�p�8���##h.������jƝ��XIu�r�����,��zjt������B��M�@X4�'B�oH1|)�(�I�b��P��zںx���rZ�.y��)�:۷�`:+�ܨM0��gyu��C��~)�)���MH���?������X�sn^9$�g�P�D���2hkȍ��}b:���ﾉ����<9a��{m%Q,�y���B��\Fم��S��r�{��+;}i���dڴ�^��I��,�c��w�)c�1�$[�>�X���[p 4��`��D��+�c:��J赨H_����3�}��;��1���fX�U����r�_"�b�^�@��[�y�o Ԏ C3�ro\2�A���
l��fs3���\�]	t#��Bp|�� �'�6�H���z��f볗�9e���C,ab�n�f�τ�H����<|^�9����1^.��# O��'��B�Ln�r��9�]~`��E3NP@&-j?����z�v����o�<l��6�V���*Tߔ :�ceE6v7'���_2���M��$	�x����K�m��������4��`�t��8�೬G�k��E��ͼ���P]�W=2!���?�V+4J��Y͏��WNu���$���$��! ��z�w;`r���#E䈈��G	�h P�7<=��z�w��B��h�aJ����M8�V�@G�O�c�J~녣�kI�M��7�ID� �5��Y��s^�U��G��cVo�ȋ�1,��:L�CRi�Yz ��SK�QJղ��G򛄯�G<��� Ą�2Uyɱh+k�;�9D;� 2v�^g#s�,|9H���`m�!.�7T�5�\�wٹ��r��Jr�X���q$��}��"��jS���)?rv��?�����,;�s�]��~D�@�S� r>ջ�d�̕�����]���;��϶ d�9��cB�`OV��7���l�!���e����lf��2���,�\��R�]��a��	*�FX��T�^��$0�V�%�ļ4i(�����,��B���FGR4.=�(�Ϟ>\Y@H���� ���h�����ΡI���Id��U��K����;XS�B��[���̉X��9vu�(q�%":�D\B�m�׀�ݣ��������ٶ�U�>?��9�[ң)���{����b%�x�%�wr'r�Y��}�3Ɵ�������U����`��˅дs'����`FR�� b��5F�[⯸Gߜ��ټ���q���w���,�����W�����"`d��=OJ�b�͆���I:ޒ���.=3�5&��R\npx���a��������}Qu�*��E���pi��wr^��`�L}�-�?�=��Lz�'��W��qC�Ĳ�U~�d���M���p���5&O�/��K��;l��Z��l����"C�nS7?B1)���_ ����A�3�h��+d�YX}ii��^"�k)�.HY�=��@!�jnZ����BA5D3Y��8��=8��ZJ)B�=?�I�q,��逖2�37�����']�ܐ��z��$�����ٷ*����-��]L��B�>��5��I�T�&��?Ns���M��M,����4Ao�؁���q��CPx��@�{�^���B;pۅr8�X=�^r���2��o�Om��Z�]���`��EB�3���=��p���S�c�v�SG��_����g���N[�N�Ml!q|K9t���Y��Bmo�E����\�i��:�=��0=��
��7��+Ǹ���V�nF���P��Kz��
��X���]�_����67�z��ԁ�s+sw���	WX��o��>���~At�O'x�A�L���/�@u���|j�Б$E��c���Fkn��Z�å��59���'B�m�:�u���m+aR��G��� o�-�ln����Ҍ��oSb��sKh������h�bY?Xݖ��L�2��+���_\,\0`&��a����p6��W��rWBF�T���a�������z��� �7Y>B�I�1�s��H��6�M�ɜ67�`�R�@FV&�QV�zl ߻�g���L�>��5�?"8!�����X����U�Sh�UP�T�V�M��4Lb�<�']jd����h�On`Rf�٤1ӹGd?f7=�<=���*�V��T�y�p!�����"X�������P��;}�`�q���L�?��{��l_�d�^�/pEb��`8#�Ǡ�?� Gj�Xj��nm�f��2y�� �
f ���xc�*`�K1���C�-^��,An���5;���kf��];\��!���W���96v7ET�05v�	oǽ7G���^˱!V��P�����+��������o|6G����V89c�";�=��VT6���K-���F�ZJ���` r��� ���n�p�~H%���d���C�26�[0�0^�lD.�ſB@bh�+=�����.�����Ȃk�%z� �}��~i��G��^}�1�*r:˝��(29��=E�$��u٨=�|\}��/���]�m���>;��cg�{�8�X�q~�3��wO��u�XL���_���$F]~tk\�2�Տ���������ͣ
�G]W����_����Ȝd�e�˒�D�N��B�O�7��������6��(��Q�4�h�����)]���t<;�>��0�KI)���v�R�����f�2/�>�<&1mJ�0���v�>`�&�:F��nz ����Ʊ���L��g����2�V�J�Nc"-��ح�w����M))a͋�#ͮKj/q�䏭�_�4Ȁ���e��Q�=�rܫ�iw"�L��$��%ZsC ���-f��G-���lt�.Ԧ3��#;����iz@Bp�fh���3�f�M8�d�M��e���2u;���Q�"d��zb<e�̍����ڲ IE���Q�q"�gv���q�y������f��S���I��4���V,��5�&��=WQE����;�@���_�����=3D,U���3I&���]�8�a"Phw��S!�s�@��)�#�!~Tg�"bǞU`���{@��WF�f��SA甞x%'��yJ��Ɉ��q������0h}o�p�P*��צ���7��H-XϽWo�#�ɕ�����	�s��q�`L�������=nd��0��v�P�T�G�&�U�߫ԧ���1���
����l�K��c{��Ǐ[5*��:dz��BTk����*��P��Pq���&4���e�'�=c�H�L��G���&1�*�s Q|ҪI��S��],��<��4<`��M3��q��;�&H�7+C�Ĕ�*e�&?t�Q����}��U7�zv�R�� ���I�65S���/*r�lo��"������/�3��H��UZ�K9�~�ꍽ>Qehj3ϱ���Ԩ
�|��~Ո�ޏZ��%��aN���z[�{������	���q��M���2�$���vuK�A�#���g;@���)�u^~�f,z�-D�k��Oۓג�#��K7���L�cC	v+M;�Gl��@��~Պqɿᄮ���xdj`�:��*�����N�~S�>@ݎ' GJ�-/�����z��/*� R~���<�-�o��z^;��̰����h@���c.jl��!�nꞹ�Q!&�8!EwO��Pn�:տ/����E�j8N���W����M?K������d`D�I������X(%�D4L��U�� "̻��w����A���0S'I�؜�f{Q�j�W�C=���X�o��qv@
��h�CU$d�{0E�Er���L�u���6��
�����T1r�p�	Y�VV�����_���Ŷ�聄�Ѳ#�g�X+��O�ڶ�q��#&�i�/7!���j��hآZ lmm����k��o_ٿ������h#ƂHc$��<�#�����w:��H�}XK��H �ೌ)��qE��wbo/X�fj��[�L�XS̡� "@�r ����]���CP��I�
�(���ĪT?�s]$>w3���D���@������^��U���'�X]*�t�79:�Rz��+��j��M�QϜ	�Q���3&l�w!���_'��!�����Ngm�3���&Uw����"��l*����c�@�<��d�
��Y�ycT�!(-��2��FGA���<�ϋ�����R�uJis��A�|݉��@���7��KV�W�l~H�t�=��+8�0�;)��2�"!�G>��;�sS�[���h�j���]��������+JY	����ہ��3�A���V{�+H��慎(d��"���!�A��ʺn�F!E5Y ]�(��s�`f�-���P:P���IR�ʟɩ��³��2���ke|.b�RT�/\����v��P��d�	�y�4gx}c>/;�?�%�S;��ֿ�>�91j�_���I�J����7 ��B�.����!o�uJ#�y�6m#�'w9��ʟ0v�$L�TE�P�*����� ��j�O���B����nI���Z��`-.�q走34�FX볷��R-4,�Uą�Bl~����qw����s���%tM�Z$��r�0I��~�1���K-��+�.�B��LH��qO���Ȥ�<g��}:3����<)�V�b���u`�BC�۴�~u����Z?�b����
�z�u�X�^����R`�N၂ҶQ�)�=g0�%��k%V*�``[�k{��l�}g ����^ٸ������A�O
G��Q`��O<�_��k�}��1�� ]��������6�[�	t�������}�OYk*>��,�v�g��a>��?�^���G���D1��n;c[�7��o��O��~����V�{���B<磕�_�B6[+��=���WW�9i���}Ңr8�HQwyF2��WIN�v�8��}'�v"�vԄQZ����h���"M��z��eEk����0���w���S�At�켉D��Z��^�#����e٦:]�5UE5<�@Lkr�G.� H�Z����0+���M.���?͞&4�Y�����ډB�瀪�SBDԉ���zP���D\D�6�C^q0շV9p?�A3^�o�Q�3I�����8Z��\�kI����w������Ɂ���F���z(������*�ev)�ʲ�⹨/D ��I�qe[���C�u�JJ����T�|{��k�T���q�v{[l�/�,����9MFА�2gu0�g7&O�
z�<�w��`�fg�'�4{߻��ˇ�֋L.������� ���,�}���
2
��e�0"8�69v�k,%�Q�K�I��y�§��v��yT#����}�~�|���7��I��2`����Q�Z���y�����b�j����&{�����z���q`����R��J�� �~�L���x�/ߥ���OHPBQ�o�=s�m�q�Z�._���1a0��+"H�L ��c��:�7�*�:�cLF'�R	��z\�ڂM�t��[##"9�S:6ܢ!�Z��ٕ�o���H����<G��k�;*�e�{��h�����ɳ��)n(�<����������a���n.EE��Ϩ�Z�E���js|�&l�FH�W*�x��Rx��L�Lg#S�͕���V�� 	���P��XK�.{��uʯ����(8� �kr'�a�2�
�_�BB�#CȊ-nQa�M~PK�ֲ)ft&��W�p�Wt��qR�ىf��14�y�Q���ۢY�����<A�uF��6cMP0)�J��@<���`]6Zem�����1�+����p6Y�>���B���2� ��C��"�8��|�*�i�7�>�3�n��w�e���a-�C�z���g��V%4����@���*>ջ��k�8c��ޮơjk���a�-3`�l��5�+�kY�b^0�A�\�7��L�}�>뙌��fb�{��=y易�9��Dx��%�G���{�n�9蒆�E�sE�d*M�3�= $e����4�)��~��A[�O��T�Ÿ}l~([P�9��;Q�Y��)�sO�V� ��>9����v8�H:��䵇_�,Y�s}짦��V����+�}�����>}��b`�љ�n�S=$�dL��z?�Y�)dw&;Ynȇ�`��F��?O�WV�O�8F�ݶrK��sJ��Vo����6��D���q,hp����w��gҹ#�l��
 X����I��Z*(�V^8\t�vl�nd�ᐳ=V��:�p�֚�v�<�9���v�@a֏k�lpi�9h0O��Lu3w���aS�ȔhlӥQ��.��������\���Hz@�L��,DQ�	�S��Q��#نg+�g��
�D����n�M�4\��V�aX�vu1�֬J��tP
a@�7�]3�c�U�R3��$�������쀡� x�j� _Yٶȹ�6~�b��f8����V9�zFԈԶ%l����V`/��$OL����n�#��Rgo�A��b����`:�0�m�)���o-��QQ�}�1W!G�֩���<�Ӳ�k���B�L� f�5k�7`���\ڤ<v�9f��줉 +c̵�~��^�Q��ʸB�]�z���<wO��3��Mi��=��H����U5).7��]������I���?�Ӭ��R�+� ���x��P�?�� <�'���� �\T�a���N�e�l4�"Zg4r�����T�C|��Y)�K��aX[��;I��7H��m����2�|Н��u�K��Bs��a�z���b�-#�D�+�oFP2 �o�*@�j/�"'n�"C�z���	a�EjYz�y�LӢS�9�߅��J��{\�瞏�����"������g,RnÞ
�����Oi5���,;j{�#�Ob1LnL�J��\�3�;���M�s�}m�=�Ձ���g�J��\������3����!&��<U��
�[�X=�P�@"�v���A/������#ȴJ� L��:�P��9�5��l��N������Ê�?(5��M">d+(�Ki��J-)�|,�\�"��WکYͦ�YT��D�C�)~nq(\�N��wk\妖��q��(�6Ʋ׫s|;�V�VZt�pjFN��^�8�f ��;�۪}]oX^�i`�c+��h_$>����$�����x�#G���.Ƕ�Mx����].�pL��Z�w	��H��� �WZ%�ħ&�]n+h_�����V4�sqˎ�AZ�
q��;oމ�ޤ���t�7!P�s��eq��g��ǁyԓ�]��/� �i<�[� �é)AԌ��٣)�p��� 5͠�����ب������+�ӆ�it�Rf>?�:�Y�U�Ë����9�Q��J,���R����`��,�}i�'��԰��4�q�����#AJ>�͖�X��U�8�S BK `�Q�u}4�S
�	Ebk��m�#V�2�f�_����G�c�Z+�1��s�d�ѩ-DiN����&S��@�t�
�������.U�	 [b�-7r�\F�G�C�y��r�ڷ�^ �X��Y�F'"O��fҪ%)� ��y�������1�*��O��w$L$�舽��2�b:Nb����=Kg�Arl�����8���U�X���^�`�c��d�$��'�x��8n0{�nk�޼`Ǩ�:���J����vy�م�l�̑�&�%�ݝ��P��_j�C�� ��.^�n�a��/u�r1��ys�M:�0�gF�b�nR(��sಶ� ƑQ�f��U�
���-~ƎT�
�$��1���;ph�#�}}�v��?�D�vk?��zsH��g6�N���� %�|i������&�d*�H�è @�x��j�W�}�R�s�W�K��8����PNi�[��� lZ<M�T{v	�A	�'���vC8;����t�!4�EPS1���`�����gY��jC���3��I�To�"�}E����zts��L}W������uY���mh\Ujڦԇ�[2�8DՁ-h�{����4�����o�JY�����vu�)�0[��P���|�E�a8�N�q��e�����̿(��r7��?�rd0�I�k��y=�UwF˙��y��<���`B�f\S�c 53K�.��q���ΥEuS#p���R��9�L��I�F�s��n����^y�\61y˟+L���Êt�N0uN�*��rN��Plx3_��GEj�����D6�`��g�~�B#�w�x�MXrg���h�z  ��ß%=���	f~�M�Ż�Y\�B�I�c�H��rX�I�%Y�����6n�S������ٮ.V�z���fX�X��P�
Ah7��9i8c\?��ʚh�}Ɣ�q����٦h��р���J�tC'*��CD�#�G�%�q*��y��;Qlmy9�!�ܫa�q,F߃ȩa�}��y��+ɨ�p^R�ݠh��:C��PRq"����'�#���	%rpP݈5�7$!�s�1��b��,.�1^�����N0j*���	�[��[��^�s8C9��?E�!�S���hi�m�V���F����X��=7B~K��5`\���iT��]]�=����w9g�R~�}#�8�C$-���w+�o�+��c��9�|�*����?6����~`Hf�%�czI��s��X�*�"-�i�;����^��tQ� �1mήg𳺐�%D-�,e�Ꚕ���~[�� ��N��p�*3�Zx(�Ik�9׶p>�~�6aӹ� ��ʧ�)qXԲ�8pu0#��'��D�~�w ���|�{��ɥ^�SH=m�q���iN��3}O�i�c83,e�\��C��,]��}<�
�P8�9{�$��ێ7��	�x�2Ha�1�{�s�H���ɉrv�$^L���w���Lg��6!b��H����2��8�j�'	�����XS�hM�<��'��Kũ&��
f�I
_}�O����?|�IM��?��x���p(���rmC�ez.��.h )����F`�E�v�%C̓�n�ۏ/�����&_>}8��;o�����Y�sl��En��ð+���Me�A���ף���	��ar�5�k�Hi����V�O�`�FO��%*�c؎�Ŕ��x�
�Mzn���ؔ�����bLyߓ����SL˭�3�wA�aY�n]����hA%���lX�WQ|ppԏ'x=UY[���j[1��tq'���JAc��+���8�}��b)���/� ����Ÿͬ8�w��{�k*@-�ڰ�œG�$�N�l9^(����dO}(qG�k�w0R��j53'��O�{�B�dG+AI`=������u�������c,�,�l�g����B��[�-�N����!�����)D���Qԩ�ޔ��
4V'&�x��L۳ڬ���E��-��zX�&���$x�XD���� ���v�F��Lϝ���@|NW��:�����%�P;�e��Tdc(�r�������{"������n&�E(;��w_�Y(!�s�:q@�,�Y�76��X���x,�4�Tᆖ�D�YP!�金tT�x_���c�D|1��/�fMv����k�;�s]*0G��t��Uֺ�{���?��Vޯ� )�	�=y�,1�b�"ꬒ��̽�J���n�t�ۭ/"�yF���q�s�n?�a��I}r�ŐqN�Ce��<�����$p$�I�s�ӍYȈ��(^��d94/�������b�t���&|$��.1=�Ĝ�|�&��$YZX��E\ J�ۣ���5$��?%a�.�i)y ���0BEa���+�N�zCk�k�I]�_��`NZ�΁ܰ�`/��G�j��H;��R�8�@�.?��f��[j� �:#��0�ТnYT�xL�jq�%)vFl��E௭��mM[%4�m��#���!��_y>O�T�㲌~(2�+;���^e[/�� ��\}���W���@7?פ,j�.��������i�8_)�D��m̆�h�V�j���B�TF������x�&��/:u�.&�a��fO\���E���J^���e�b�=B�m����q�8_q��vy�Z;e�->�T}w� ���A��Eu� ]9�Pd������B���	�������FR�ŮW�f2BF�������_��Cms8`���jҳ���Ltm��5{?C���\��v�a�@Y�}33��7{�׳���N�`��\�����}7�K�'o�h��KQN_�r�)wS�i�=����1Oh�?��	�[(���y`��S6D��N�V��Qc���;�X� ��g�&�?N�yZ���_��kb#6%ґ���"��f@���21�e<��9���H.�,�O�91ø\I=A)���˾�H��u@�u�lY/.����Mu�vV�4e�ܺK�����6[R��m�#-<Z˹�,�`<�r�a�������~j�M��6h��eX�0�f?gXH��_iHDn�lP\��A�`뛹�����/�+W���f�c�]e�>O���p����/�*�~g��y��j��-ra����DT��S�N��N8�ʑ�'�X���p�VS8͐Ar��c��� Lf=�Д��Rs��ʏ8�����:_P���Vq,L=>��rZ��v�P�<z|T'��;�l �o�D:�d>��1&�ݩ
��m��bs�-!��O��!(��y_J0�����8�8�:i
�l�2z˫��>:hfLQT'G�}�B��O �f;	�����`�����u)�xb���k蒞o|�Xmt\;4`x�lʔu)��d� ��2;��圹�] �/�P@�๟o5ʮ�ЬǞ3Ï>c����oV�O)��Vr#�D7�; ��w�o�"���%���?L'F��7Ȉ�'�&1#����$�g<�9���H@�zτ��/R���V��ɖV��9��[�.��P7
5�E
���3��W`>�R��Q~S<��&�2q\2t	?�'&��=N�_!��g�c)�^:�l���p̥�I���i�j['�p�.w��Ǫ�5�|�"�QN�G/� ;Y���v5GI=nIG!+�-5Iٳ��z�����]Y��p��U#��ZZ�-�}�U�,�V�qB��cd[1AR(G�iM@�ʧB9�M�*$pWk���4�KF?w���1:�Q�n��2O�W�������Y�<��;r��ohX��S�I7�DJ��9�y@�%F��&��F�^̦Ѧ��]U��@28��ؒe��4Z���m�+�/T��ꑣ�N���� �,�Pm;Z8�F���b���1qFZK����w�^���z8K�[�5~W�}����G�!D��2���b ���nH�A�3y�F!�_��7v��>����O�07EWG�\�Ub�Z�m��$���EnN������)U����_9�}q.����ΑҒ�qxanS3/��{���nD�+��5K�H7�|��n�>Ք���L�&w����S�qO�.wE�������#x�pt���89֤�A�l.�;5A�,����k��F�Xn�eO�Q'?(x&�> �hS��[����30��لu����/��)J�U��"B�Y��gk��P!�?bX����
wd�)5��,D���	�ŉ�z[����#�;�_m��z�O7�;�ZT�$�8��J?�_2-#�i�/~���>-'�>��.�����5�y�b5�xa�N� �������jT�n�݊��C_�srZT.��Ɇ!~jh�b�����k��z�Z��K�	٘k�ZaŰÍ~��m�b�Ё]�5^��|�1����\�v_ ��G97��U���L�C=�p�J�3W��6���Uk]j`�a�`&[jE�Dl>4H^�J�B\��φg�1�X�Tkx�`k��K�kceM�k��O�AM@>��	ϓsiW�ђ&�;�����V�|��<��ew:�����SX8�:&&���!_#�$
'[8�8��	3iѮ����x;�xu� h�>1LJ'�
SA�$�K�{�7�e&����f �x
w��a=�Z�����(d7Q�}K�V--�=ơ�@�����AD������R}�E�V�,� �%jл��D��}�����Ʌ�Ǟnc�
�����џh�������]�:/�g���߿,&̌�;��8|�n���+#+M�u���#\2��S�|r��1�^px��D-��\��Ӛߎj�M	�O�G�$"��B}�<���Ԫ;�0g�R���Y��0�%�/Ɛ���Z�r��6-l4=z�T=є�Z�LsO��t�]篱�i��"w����H���]~���|���V������ ,�C���x�%-hX��hj�RN������N,��*T9&'+iG����0!�V5�Pξ5������x�YZ�EvX��'�����CDS�F�e����
�a{���R������a�C(b�����GT7^¦���,U:�QL [};���ѨH�YD"��ħ*�=-3�*���5x�G�ae�2����ҷ����W��r�O�Ӑ�	L�wj�B�]&ͻ���������"��������>Ҍ����F��=pkOP�͍�ȯ��ʿf&S�H���D��>|�5����}Af@))�4���Xl���b�C��%6�D$qF��V.l���n2���m�^o�<�\/����m�S
�Y�|���v���f�׾ZE'�=$ܡ���#��]
�\���E|��\���a'��@L,&��uE�HHb ��~{ۯ�Φ�g5㹱F0�B��2 j�49�?�T�q��f�ju����Ԥzux�����w��	pg�0��t��PI%���B\���g�U;�'�*���6��J�bS�u�w�;��mL��Q5�{5qB!Y�ʗ7���s���u�`�7 D௺�S����X\�;:�n=~��P�}�#@�^��fnE��ҰP!���Α��NC�+�
`ֵjQ����b[Fֈit��x�_�o���"�^lp���p��h�65x-��}�����x�v?ޭ�m���{+��nY?ݥ�\+?����2������9}ȉ+(�xՁ�ӛ1g	�|,,�ԉ���^�����H�L��|��M�Ef��H_�J��ں�\Pb;�-:]�J�厁�xV:m+�d㤪�$�.�`+`긋�B�\���-D)�꓎��J��<�B ԅ�7����������[�v]7@�ɾLl��'9��_��0�,��?���J�@~�ҳ��JwF,��&��n����׼_�ίʴ��mh�[(ş�����tG��N�BäLpӢ����Y�O��4X��@\d��iP~�����*H�%��8	�Ki�p=a��F�U_��y_,�D�`վ�$~� P`yy�2G��$ ���<Ux٩G#�?�a�hS��>�貰�ۂ��{�s��6p��J$���*=�E��_���w/,$���d�K<���( �-D���;Z��ps��팥�'���2�6� �J�}9����^u6?5��k���r�K1�gwng:����g�.R��e��xk�U_��T���� ���>��
�;�!���^���C�$s)NYXglX�"����9�|8�:Kvx�P|��V��Hlw���s�0���Ɓ�|�г�B����α�nM���������лZ�M'��=I�r�<9��ҳ��	=��׳V��6L�9e�?��k6���)JU�y��#��Ѓ���>����QI�ZΔHE�r2���En큹�|m���\�߷֏�Q<v�O4�o��ʃ)y3��dI'Ҕm3^���j�%�SM����F�����ޘ��q������gω��V�'g:a��57�s�9k|�T���4V<�7�Um�]Ҧ9Q;@\�(�0R�8ˋ��I����
�L�f��&��^��]���g �3z��SY~!S�3;8��I 
��r_�J�V�6�dyς�"�w`u�Z���ܩr��R1���A�v�椺ʑ�:�Υe�!f9^P�l�:���Yx4�]}��?�- D�e%�X/<��S	&�[�O� E��dl� ��L��%�C��sV�M~���;^\)�(A��I��YO�l^njv�vA�?�B cgX��H���D9��{!��iԳ{�Ć�	O]�k<w��<���V4�{*��?ϒs�ѫ�G!8���	�wk\�!`(����2oV�GGt�љ)�)�"i[K�d�gA�"mj}ݙ�+��.���t)�6S�G���G����ԟ��N�X퍞'��)>�͑=Z@^p���vT������H�y�׳Tt��X�. E1EX�?.;�N���R�Z���Nsj�i4����4ǫ�H�c=�����p�m�Y���X��+��Rz`ύ�������.~��R☑y2� ������?��b�m�CY�9�?�7R���k$�ts�G6��lYlٶLI�~�!�OO���ӑ9}���T_ (����t���s$��Z�K����i0ѸI��[�2�z;�+�%�����#	���P�8�&�l�a��M7�uH}�R�PE���|%�F�K���+^�@І7�)�7�Kg�� R�1y��s!x�/_r�ޭ���7�֫M�r7m����L��@�c��*�k7-dݗ}s�� 3_���>݅ ��5�w��$�� ��o�bɾ��>*��u� 2�{�Ǩ�{j��  �n{�2S��P�֩��%ɻ?_�x����4- *�H�~>U�1o�q��pkL7��4�x�9J�ljw�)�Ϲ�e;��[��'���^ ��r�%3l�Η��M`��*��Ѯ���[e�A"��>��nj���X�=�O��Ċ
*�u\��w��>'��M�X!����ie��@gN-ѿ՟� �3�{+��W��ј�iꪡ-}� Z��9wqBI,ޭ���~�`~8��t�W��FH\�Ԡ���֏�/�X�kQ��
�.~6buL
�AG�~�����Y���B11֎�ۢ��x)Yã^�m����_���Pbf8S���
)����I[o?�V��LR�&��ȣ 
�����Y���c=ä��P����5	Un�&12��������J1 ��3��%�� c�M�DB��>�D��N�T��}���Y�U����C�	b'�����4Z�0}�V��b~��*���:��3B:��3=�%���\�\<�տ@a lz��۳#4*S}�K�<.e�逸c2�^ɰ`��ny���]���͝�8a�Y���`)�Ĵb}��Ǚ�N�9���!'�y$���ir��;�\3)h�v4�&l<9lA�w�ceS�'���BNs߁���
B����#zh��嗜��Y�tfV���!�0m�
%�t�^�l-�x՞�+ҳړT���ܨ��u��-�]1�)h���u�%�Z	���ޱF���$�����Q�\�e���b�n�,$>���N~��\)�����PYV�ژ�W��)�x��!A��U���ݦ��kv���.�P-yFu�1�L#�I;<�!o����G|g��eS)�&�Cl�p��!�AO�\��.�)�Y_�u-��^��<��B�+� ��g�� q�ƪs�����ҥ�1����Z>W.L��mmx���N8�mu_�K��}������3��`=�eC+����(���)A\ �.��:s4#�*����?��>hba�ЂKW�6`_�U�dn��5�8A�7!�V9�M��u%�8�g&����(���'B�� ��>RL��˛���[<Я8���?Rwg���0_�%6����*�f*� �����4o���w3���=+G)܃��q髱d3�n��J�~���Z!��Y!��hͯK%�m�֡�Pq�3Cm"�ï\��ɰ3�bM�,n!f�$�5Ox�6��߄�`���N����N�~���O��'����劒p1�ę�rZ7"q)8Al��Ρ���̞�p}D���nN���`�X�k'�M*}����}�O���|a��?�ufB<��OdLUb�X%	s�lK�C!�p���a��&��:e+NbAdc�&����6Ɗ2�w��K�fF���SO��w�	׻j��E@�G t��y��l2���rX:Uqc(�O�}�;����i���c8��z�7u�x�#��̑�$�z;R��Ǐ�t_Mc2a��.�d���P'�W�guI��{U��^�
�4o��8N��[� �RP!�D_@�Sa�-�\�~L݇�d�(���ä���^�~�nG��]�A�mN"����}|�KI{�ŪpBo�Ў�Ӂ��y�b[�D������ԂƇ:޹�AX��=��T��J��̳usC�����b+�����E��W4ZMZI�9�����_�Ӿ�?�K��sa��	�Q{��TZ̧����݅Ɉg
#~���i�.�X�/)�^�'V��O�3l��%���6h̜��5��#�c���+2ʲQ!�P|�(:\fm��dZ�n!���UN�d��6��f�`aҘo��r���E���9���&6k�5�[��*ZS"�\�?����v�B@ߏTC�2u�����:{c���`U�Fȇ	�[Uwq��.�Qm�G[-d�^�j�{����\O�ERmN�_ M:sp��kh��s�y�����R���@�9���W���}�:mK�!f�k������лjR{x��Z�ƣ0np��'��,~�t���p�����D�Zʒ-*�����[L�z�mk&s����K��bQt;��������\?�S�����.
��o�_�r�*;�ML��.u�T���\:?*[��ؗ�%F��ҝ���)<�}�e���Enf�r]�w����&7�.욮�n]@̡�������x$I�a�$�����/����v��pw;����^[��F����7�������@�<�g��ǜ��+���9����)?;�C�1�:s��.m�F��]
��N'e��q��b�������2��Sf%{���p�+e��ర��}�RR��{�A(�gL�g	�h��<��ء���{�4*��Я ���L0��k�x�l�c
>0���Y�Gm�1a��Ź�BEH����?n8�շ�oW��6T��AW�܌�f���,zj��Ŗ'�`��&��"�#���\��Zq�T�:������ƨ��{>��d�z���\V�Eɽ�|eD��O#ד0�q��t/��}�o�G�[�q$��e��eC��/M��"r���w����ض϶��h��0J�#�$Ω,!vD���D�v��������7;�J� �ޝ��X���g�����g�W��)��ĤJ���ߨ�æ!3��s(��tK�S3�&����k5T���0F{B�� ��8�	߳�o���[�:D-�]H��S�������d͟�o�^-r)��.S鵙p
��!A�Y����ʮ�;�B!��p�5M��=�1c_f����:�SV��;���1������&T�
"�-��%��r�`��b9{��Z���N���á"��0eB�v�)F���>�Rg!�{f�Nv0&T�B���I-}޼x���/F��ӗ��3�e-�	s�
M���x�}���C|��0�EeA��1
jP�����ا�C�\�^Y菗��E#!7���v;�`���"�RoSB����!R  �lE��)���f��l+�dO�1�"(�w�������>�s��d�q��S�E ������WjN��|�bj�(ӂSY���[e�� ��oˇ!�ހ���my�d;k.�'*��:�t�S�''�[����c�T&����ҁ#�E��ի�p��V���J�Q�!=K���F+��EI�Z�>P��!\�7�18�n��06�?k��d��Dm��g`߇&�dvkћ���p"���z0�2��]��s*j��:lC�H��ӿgK���`b ٻÀ��r%~{=�����!� R�H��aj�{[�,m1g���y�0��ċ*�ς<r��N��w�R���l���B}��b"�@x%N|z�h8��Y�X(Xugӧ/�名1"�u�r��0>[U}nՏ�pMn� �o��%�֭�E�Ç�i�[�.�^[(\7�݌pO/��<G�̃�u~�b�S����r\�� �W����!�A,BG-�K>W<��3���`�]����`g�������B�rh���� �L�u�Z��L�n����:Zp�T����Mҗ������1Do�����4T\������|�wv�rRU��VLWlk���1� ��Y�S��Ċ�A왵��û��Q�a�������߉˶�OR���D�����6\��`Q��4M�Ѕㇵ{�<~lv�:.AI*h8?L�������BS)]��H���u�c
t�=�̀�/�}�Sy��<'�L����{5j4^��6�W�?	�_Ӑ%)�P$Uf��C-�����>׫���!s~���v��-> F3[6z�����%qV����XU���> �2�%:'O�P��%I�AsJ�,��PA���i�1Y�0M��Jv�/���Vs��N�\���Cl���>7�b�b��y����Q޸������VLu��&@K�R#�`ա;��Hd��,9��ٶ�'�3�hsPn=(Ĭ��x�v�+���~�#h��=���hU)���X@�m�s$}=n�`qᆹ��)|��z�Z%�����^�yx~�����y�[eG��Lf�r޼V?#3�� S��u3�O�q�8]}'��MO$��Ҽ�VX�$Qe_�m��o՟��ć��ŵjF��l�J�
�-\]�����9zz�O�U5�\�*���O��Q A�G�6c�0�U�BH'2I4��������*ݣx<Q��DvK��̃��E�d�d�Z�C���������d/�*�$���%)%�?0;aB-�2����Aβ��Ŵ ��a��f����2��y�-�w�`�Tk��S�잳��Q�/[a��O�_o �,Vl0�;$�V��A:~�s0�� �<�H�Faǐz�[-b�׮,�8i0'v��u��95��g5�#s�D�j������<��	�I��ک����/�:�R���\�%�B��r�y�f��^��/�ҮqB����|8�:Z�+����;����������@S�3�T���G�����/�y���"��U:ps�?����&khK�_�����x���PL�1���ͯ^�4?b�V��H�R��<&ި	��+�s�����YZ��9ɚ>X���Vlm�3kV�W�M����
�G���k���t��j=g"���bV���^�A��
����h�������iC�\Y����
�	��#�Oj�eM�x1#%��Kӽ�*�BS�Uh���NBO4k1)C����ϱ`�ƗE���� �/'�BW�!bb����O��,�� �_�Z?u�恫�5n_��D���ސscT�?��!Wx]��q'<�.����Sp���M4w��{�݀��(�&Jo����@	ʥ�Ϊ7�=;xwCB�+���]�g��dup��z��1��k�Zk��A�V��(��"�0[|_�σn6r9���l�zuڢ�1Қ�VE��WK���F�b:lg�鞔Dk���J�|QB�2l�g	S����S~?e�����lT�[P�LO� ��(��̠ҩ�4<�"st��uj�.j�7�-|�NlנK^�ڞ�L�f8���<*=*��C_,�u�2�J�?R��ܱև�2���V�d��o��tf���x���D���d�z�� r��)����/M�{tk@3D#.R�5�G�����/qvS�]�G�xI:��ԳUY�b�u����+�HDA|�FP�͎\�0.!��Z���� L��\�N�R���ûN��z19:���IJ!�yCm�䃚�w&�2`Jl�,����a�&��&_�x�a��r���3'��H�0s\��{=�61�o�O��2����v�[:��;���ؿ��z�P[���N�Ex�� ������:kEy�?APY���޲��&A��9e�&�_�sx�m��3~O�.��ƁG��^5�\�X��պ�����-:������[|�b>_�݃<\�����TY�;#M����)tGF>��]�!�RSǾ�@4P!(�W���<͊2bs>E��=��Dݙ�U�-U lp4�H�w���۪��]�|�o������@�k��	�y�n4�Z�K�Mu�*��rf�bY�����3�x��U�7�R�i�>N�	���>���0�+�Z
�M�z����4��Z�����Li2M��ڐ��T�x�� #T߭�2�QRE6<� T�w��4�K%��p�Rx[Y8�,Y�Qs�%�H�3�#2c�	�
GN�����x�ܽGc���g'�Jɇ4�D~j�J��N�r]�y��Fn*�i�5��޶�D���mL`�O����C4��H=�k�`٠������ro��+���;���O����2W��#�և�q��S�x <4Vt�_W���}�𱐘6��# ȈEן����=>Nf�ㆭ���2���b7��>O74`2���I	��I[v�O����e�5�A���V���B�M��W�<���M��|��&�c�O/$E��p�/��?Ah�(s_彰o��	��ѶĪcp] �;�.Jb ^rHX��ay��p� V��v�1,6'���T�v�e�*��H���& ĉ�a�'�AƗɖ��ah�����q�QH�D�R�:����'�'՜8���n/�n�p��c2������}�V�����C�1���ځƁ6=q�ns�����$��n�&��m�;.�?�q��o�>ZX���F�����=���x�I����{֌d��H��b=��͡���ޥM�Ay�\�gq9����}�2�&��a���ar�@�8��*��#�.7BD_����w�]�d?�5,vJʵ/BT��[£�3Q��^X��<v��������qXEJ[*h���a�,gʉw 91���:n����w>@\U�=���O�٬��Ş��e�oc58���Ag�T�e��.�.����⌅��]¦�^s�^�h5���"Ȇ]��l�8n9*`u���d%FI�	�Z�Nj�<5s����P_�/g���~�r�SxN@7�Ṕ%rl&���p���~���x�f�#�������J:��N���`�;[ͨвSA�P[��}�G�h��IÑ_b�Y+خV�������E�'M��R!l~�^%��hN!>�*{��BD��q��w�C?�̿�'%F�Pq�i"��R�{E����X��t&�ڰ{w�<��&L�!�JV�U��ȹ�l��e�����Ѹ�k5F~����S�f��,+���:�r�i����������w�ؕmU�
f$dX���aW'�P�-�Y��u���f\;�Z^��Q<��ݵڠD�Ĕ#���x��K�+~_�L�E��CpYϓ.�JV��k��n]WUӷd� �S�n5�ֳ?D��I 0#Cq��u�J�w���f�"Ħ��z:I{���[D|׬Z�����_�Wsw6 ��Ȇ��u�,@.��!��ZxE�M�@�� �'a`�"����arT����;Pi Ԕ�}�5ނ��)��v�2���x�MwjB�p����7v�?[��_�	�u�� D��+��*nno�9�b��ڛ@k����=(�81O�jӨ�ͼOP �1!��\�ѹ���MV=��ιE��xP�E#{�]��>k�^"��?���w3�R�w��@�s�,�f�!X
��Af�����|o�U�@t��o�r��#d�NO�`�&���t��ƅ�s�p���o8F,�1�n}X�7Fj����cq�SY�>�&¢�Qv���r+�K�NS�A��ZU�'!wNU�}%b�MC	�Y����#{5pS�H)A����OziM8+���ۍ�t ��b��@����ͦ���c����׎K��|����P� "Q�����	Ų�	ǠM���>�u�N��ʩ��#�����<z�����r�>,/4�(������Lʶ�5���:C�R�q��97!,����3R-�T���A�{�,w���8 u���g��`K$�m�ӤZh�4n�_�S��5�n�D��ԝ���.b^dD���� w2��yw�$�z�\�KY �?QPxF/=�-NE4��u�S<-F���7J9Ռ�d��/��YV��)�sl��9� �����& "vI�o{���S��>�k� 53U�8֗��{��w������!�F�_�Ͱ���i��3 ����Em%�<*��Γ9�J�+�Ch��umH�!��u=Bf�����V_�AQ�{�v5���}�*F)٦QX��k�h=�������|\8���u��w�A5�F��̜���?�^��_e _�uk3���n�Ig*p�Iiä/Ɋ#�ZC���<����(:8��/a���i�wY�Q� x9_	�������8'��?���Po2#�#�WZ�z��v����>�%2�`��"s��V]}\�����h�8�LI�y`;����<az���8�����6|g�U�'3�3�R9��6
�4 �*(�'V�s����.�5�����ʤ.\/. ��5�Js|�)3�"j��b��U�-�G+ b�u�b�z��<�q +!ӯ�e��q6ߡ 	��?��O@�hg|.*�"�Biy��6����%*1fQ:�끺�Q�ܰ��?�9��[���g	i���bu��R�^{�@�+�Y�>�� y���Qrl*6#�r�����@*ثGȆ0iXp-{���?x���'��U�T0�Ad�=����<��|ɫ�$�+�J�.�nfh�Z��� x_C�sD��8�������Z�yj�"�֙5R��!Ű��M|��u�7����d�	1D��X$2ǵZֲ���3n��5qx�1Q�V��,)�joF9��x6ah���~��i�u��@WaS5�md�FC���+@3����P�9��rw�̄ӸѰ�,��&������ų��;2n]h�L[� -����jI�x���Q�Q�_���=ϴfl1HݑW�E�@�U�F�ӄ\��V�����`麜500��!�=�E��x��J�� іmd��h�c�ɯ���;4�5` ޵1������l=�YQ�o�KϓoJ�_�C@���w팎��8l�%V��c�KQ��.e��JM�vD��y�R�U�X�KBI��^�?�VU�U{P����ɸ.]c�`������o��D]��� ���Yݶ���:���qo����o=FR:�.BH��+�ﬄ�^�u�3�v7�,\�+Q�t��1N�����t
d��~�P���#lv O�/״3Ĥ��t���[q� ���N�ei�zie��ڼ/����	��uH ȹ.�a�?��ݔ���։EYkC偻ө;&[N��D���~���^�^� z!�����@����� ����٭�\��'�������Ma)�*�Y��@3�Gf��h��,��KK�'Њxp��F�<�M���m;'ڪ�!#.q^2 v�����Ak���<�U�[	.�:RAo8�!?6R �sHP����ݢ�d3t�i��*�C�Cov��B��o"�K��LC��U�̕���'�uH�ȹ�����J�i�(���m����p�����}П/MP���$�3����V㞭�-���U�8W� f�Yh57*�۷�25���sh6��m��jN<��>���^酄xq͎dN���o��ud�"|�>�l���O:T�� S��{Ŏ׻��xl�Թ&�J�27���c���O���wy�O|@(��
��M�!�H@Ih5~3u�.�!CV��2��͓SϰELV���-V���TЩ���|?vU���h�8�i�N-~�S��l+�-�f�T�^�Jp�m��/&/�b�BYx>IkD��R��|ϡ�V˲G��K0iz0�"i�ӈ2n�q%�wWX�%���Yieς��`��>\K���K	�<z�L�:��rT�l��������W/Qq�(��.���Ҥ0��a.M���LU��F9k�ET�כr�π`��M����fy�����Fi���y^!&�s�� ���`�>^�FH�w�+��������&���;��M$�"���M�����$VL��Oe=��ٻ�@�{��l,pl0R����U���0E�����S0�R�51Z������r�+$����TFW�5i�4�w�/{LT$jC��>V6��3#*�%�z��׃#M:� �u��l��צ��IVU���=

ܹuY��o�uFE��a��,~���z��V�8��2�5澶�S{�	T)��|Tḫ"���O�偲��l�c�+���pl��1 �Pp�P����U��xf��<T0R�D��dXЀ��Eօl���%]|���r�&�����s�8]��H�+��G�Zo� �I�)�łL�6CObp�pM�B�&C��A��\%�7�w��d���Ȍy�L�ѥ� �	;�$�DE%d�p͍�Ӊ�}BM��@.�#�g�bi��^�t[h�/)����U���'k������$ܠW1i?��gp|���*�p���YX*��������	z� �mu!V������
��:YtJ��`'���5�>8ҏk���Isu]n����At�9Z[�L,-���3:5��J,l�%��9w��\��`��+
�=䫡)8�0G�a2ӄsY��V����9v�>��=�>���=ȗu65�|A*N�w�Tw����_M].aӪ�wZ5	$���!����Я3�Ra��L=r�jRXxJ��:�'\�h��]��j�}�Z����~�� ���T��#y��s<�^9\s �o��Y>*�3� =�����sL(L6��F�;�ͷ��{@��X~}�&%�K��vƯ���%�m��zm��n43�0P��z�������o�[���d���d�翆�d�2'(���{����B'sN��1�qy�ƕ���_�ͥ�d9\�J!�����J"�/o������w6>�n�������;\T�u�u�M�/�f���mm���{\��9$�P&�n�<<ʒ�i�[ub��k[�#�u_��Y �%��8�����T��� e�~��z������~��G�V>UC3���{�r���߂Nsa�
�]�CL��5������āu�+$����M<�?ׁ{1G�H�.�E�2��ͭ?�dC�Y��+���,wM����ׇ��N%�=�.y陠e�G��r���Q8�1Y4��XM>w���kx��2�\w��}����N`wS����پf�KZ��;ݳ�*����h�b���nE�m9��=O��vg��(��06ާ��&1�2�|����Y�hu��:M�
d[1����H���n^!7��p��h������О��C����K���^*]�>&`I�m\�тr�F�c�_F��D1S��y$���4%��^���}��w�*_��Ѓ��@.��]�	n��AOU�-�N��ǵ�r �8m���O֑2=�_v����L����Q
�Mb(g@����_����=�8Ⱥ	�	ѡ�S�Zt(r�Qwo�v�e��GZ��e�R��7Q /��/Z"�0n��Hw�r�;�ȑBVr�r�SI_N{E���ai���%�s���iK��R��%:�.��lɶj�ʈ203�py$�.�^����3W�@	����Ҍ�aj���0�k�ۂ���J�Iu8� �-�y�r4n�͏-2�|؀�I=.��m���\+4��X�,�"5W��oK˝�ݍ�: \MU_��Xo(�%=CR���.����wg��e��/f[��೗��е���փ�9���O
��J�֔������V������>��ʰeS��Q,���5�dI��]�1.�NvS!D�t��Mw�����b�`��� �v|*c����?�*�t�����BAR\ݹ��sf�6;p�����yV�%�0ĠcFS�b�y��Z_kA��$��#^o"�jv�����L���W��XF��Iq�M����+Z�e������3�aÈaY�G�C	�)>R��(���mY6��]quרor�������n��\M�&f���7dp����z2���/�O�̥w��F�G�O�V�%�~|��G�6�>�1G:�!���=8�2C큩�}H_-˺�U�T�8�0�smǹڿf2�Tq�qd�(r���k���ύX�v������I¡8E\	��վ��{�v>|���y=���L�ѡ^���'�א������7a�n��:9b����fd�}	�����<P��>�D��}E Q�}�0���h�e�f�md��leyDfa7��c�<��#�A�L�NsLV������X��/�y�	bv�=��j�&��>�w��M�Y �tE�H_.O7��Sr��9ǻ$3ak/0\�Lt�2c[�	����8S�Ė�|�Յ�pM}D`,\�u��}+��-mo�9���!s�m�p3H��6a���T��m������w��;�BI���w(wZN�nA^��iT��X�c9/�<�P@�$�%��_ˢ��{����&�
7�]kSR��Dn|[ݫ��Q�R2CªV+���]�WpHG�4�Uk���Ž+�N����	fB���މsM��4ة��Ms�H]��n�?�����b������6�D%@����E�Ҫ�"��:�:���/��9;��SK�<�Nh9Ay�EJ�O����-��T+Ϥ�	:	<����^[ϕ��)_��ʬ$\%�cQ675P�f��-dP3�hR�ͪb@�hM�4�+�$N��@m{�\y[f�������������ʜŧ � 5Y"�: �~L/�΋�?i�>I�KhIx�
D�̲�<�����������Yeӳ�P�y䲢���u���q�7�#�96���Uۄ���P���W���!Z�m�YF���FRь�8��i�{+ۋ&��-���䘱I�!�e��q�T]#*s��.(��ʘ�E���8}����w��]&�Iw�5k�#��5�y��C�>^O�'�2ăE"�D杊E�FX�ɇ��c g�_b��t�[�V#��퀒O�S:M�}bi�@�"���ޯ1���5MSS��c�r�߫M.�	���~���U-�6��*X�B���B*�j�:,����Ō{Xe �Z͙������C�s�.ܤY5�4V��>�c��U~���s﹐�\����Do��/٩/��o��Yg�G��z��d�nlf�z���˩�)/L��j��"�&Z�Z��K�Oh}�1S�����#)%��Y�M����:2zk �z�<��W�]�H�����}���}�M臭 �������&P��Q5��B��I�o/�AQ�@F�-�Ш�?J!���8_�ܞ�Ӽ����?�Aa�
"��Vq�0�F���i��ѕ������W%~ zm��K�y8 ���BF�n�U��l��]*��8�WܚQނ��i���Vc��R�*��\�����❛���i¬B����l�ת0������6=6:�Z@/�Tf�ʓlrc��N����0{��7@ >k���\��G�)~�� V��C�e<]���P�n��q�M���R߄|�]�X��BS+��#�,�.Q�_~Qv�cа��N�_��|����FN��� J��;2��B��S�;!\�yf���T.�
�/<.}m{��o'V�L,�B�L&��4_Ÿ�gr p[K�5���������P�����v���78�EU�M̂��t���3wí��%���M��(굆�/f�+^�k���ݼcIb}gQ��x�0������G���
S)#ilu �q�2G�Zvh�^zh�#~�M����?��1tJb������m��M�'$X����[�F#r�L��7�������~tF��t jO;��@8	Dl�%����2�y��"�[��"�=��Na��Wf�4䖖hd\�L�^���{ �[W��o���WUk ~�Y=�e��|V�$��#�-�ud�`�?�O��<��Յ�b��e�_qi��d�x�) ��d��q��Ql�FZ�W��N��/���*g��,�5���&�C�y�/7�َ�t�ib.>�����%إѯ�'�Y��i���'���p��q��K2�m��:&�r�)9Qh���\�`t�O���1#�UUq:��Z�l�U�F��<�� �w9�<��j�:���E���d���o't��O+�WQ�f!��q����y E� #r�\&')r���B@֙�A�[S���k���8L�S`ED]����!����--93D���{�������c/������G�:$�&$�ʨ�_���8l���թ70#Z�ϓUj���(
��'�ݲ�7���iTv����E/�.�[
A��i�=<K=@��� �e`��x-/u%6��VR��q�0N����]eY��.3�q��R�k<�ǝm���P(���{9,�n'LHC�'O����<�._D���[J��d�F��HJ䪩Z{�Tw���{����LS��%��f~<���Lƚ�ϥ�F_���nC_h�p�gm���.x��;���98"��ǃ����Ɠ��v+���X5��'�5����(�����Ԋ����gA�^�;J��%6q�@��sz�	�3[��*�������u-fַ�"� ��T�5�:9i]w�ȋ��wm`��]l͎���E�����Jg�t
L��E@LRPe(���|�^^�� ����<$&!�`�cY��.�6�A�GR3J�"GNk
�(��톰eJ�;�7�K8i~��yX_�J��V���uC��P\I$ńN2n~�`�%�� �1V�����|������_�=���2w7�J��1i �,��]LD�"� I7T�ޫq�'ݣZ]w5�~@YgNu�C�o�P�%��=�FƼ�$g�-���׋&1�AP�-'�����*f�4y)�޸�ʅ���v$_�]>�ʐ~�٢�4Յ����~.7��ٌIW�!{2.	h�BwLy���\3Ev(�4N"�q��5u��>x;-��EU\vnG��	͏K�)_�++��N������g�o��N#�(�@D,K��^Qc�V[P�iv�Snpĕz��_�i=2�!q��������r�a��z�]sU,fs����E�X�H�s������ �JE�'�5��:����Md�9@���fO��uM��K`��AV�	1�~h0���9 5�ʮd�=�@�0�`=#{U@�?YM/M�?v_Ы^�hX8Oï���DI+�*�Dh�^B��;���`��g���$��{����l�J�����Ζ�L��҉�POX]A�2v����,���FM���M|������GN��:=�b�&殆�:Fk�~�O�;�mF��w�ql<9�����1�<]�ω��Y`WS��&�r<���1S8P-���tL:���ꪮ�:��ԙfտ�e�Ir���&`f�<v"�T���*m��[.?�Ew�k�62�z���k�0\�l" hr��H|c��޾������?{C@
&8���r��:�T���PUg.S
����⎥$�Zs������W @��� ��C҅�$Q^2?̿��fۨ���� �h���.� 5���1]�3o|��)R�A�o����n��񻸎�IY�_�B�����|�!���N��AQS8�X��{���d
�y����,pt��OMwm�_W�.�FSk��Sc� ���/Ҭ���`R�eȹ�阔f}5��p�>�J��	��r-q�l�����Z<��`V��9,���mPIΫTЊQ�Xz}=��0H��'U�5�`�NU6$��ڨ����H��-�c��p�3+���Hbf�f�����|9Nf^)�2��Y|S\B�=]��R���M�I���m�O��a�G���{�O~O�,�	�3���$����_/������8��~��P�+[�oßﳗC�L�q��EPP�����V׉W�};@�� c9���ko��0z?
_��_�]Z��TVW%�*c���P��;h_g�S F���ė�8Gp<. ��r��۠�$z,�9@g��#�Bm�{&1O��(Ğ�'�g^��[qmǐv��%���?S��d\�0��nHc���mLYj�C�E���gE����<ξ�CI�z�,J��Ġ���KMш˛m�}a(�6R�|�g��f_���-�X+��9���EH+�[)-;y�D��s���Q!p>�y�����+$�0�U5�pdR���S�*7=�Z�mo΍����*&�� �Ԙ*K[d�Y��yjt^6n\�5�0�˜�Wl�-a�����i�Ի�W�IK� Ҷ]P란�V��nI�Ϛ�|�쎢�Ly�3In�K7|�@N�6�Y��m7%�Ek����q{��5�}p��F<�f�mr��h�Q��&�_�'�f��"@?� (���h��C!Yʰf��#~�����i\��aG�_4׈�F����S��)ې8������1�&�RE�P��@l�S�~P�O0T�=�k�N˥�G�-G�d��ZN+�"KƄg�-"�b]
,�ŷoK��.e�4(�(�/M�H��(6�ɗ��D�V�D	����Q�[��Fe����I��qƿw2g���rx�%�Րw߁��1BS��m�E/D���_g��l������?�s�)%ۦZ����Ȣ�@���
��l�m�<�hބ<=�ȱB�� ojCZ��2]ɤE��!�b<�!�1�w���QG8S���ץqw�a䐋M�|�(��:����xp�7�%��4�|©t1w�M���;Q<��$Őn)��Q�^��>�X�'EL�n>d��s�5��S�4T�:��w*W r��閙"mP;����9[K��M�;N�~��Hk�EM��mS�EU����Wo�S?8�N�#����gyI� �q�׹i����b� �������*��7� *�`���tA:�l� mz*�I� و��K}D��[7��&�e��]#�7��*�d���6F��������~
�G���D*�f���;������n�W���3�� *4,r����8��%كE�2u�݀+�r����(wPO��>łn�%�~�!�;d㏰k
�"���)f2
��
T�ē�r��,�� 	4�e}ڻb��b�"�4�<�q�����'���7���ŵf̘���a�RD8ΰ��F8�uNO�_~�O�*C�����辂b�㰂}�=�1��CS
565eU�\"����ٙ�m��Ѱ�܈LR�a}�����0s�M����B��k��!��yQ-�@G4��:L�Ȃ�%:�5";�}O��.<����@��^%���v5r��?�_i��;��4$���R��,w��CS;k��Ңن�>/A3{)O%�
ucd]o��|����.W��/v�e�R쨣,��;��,�7�Śչ
<o<��U���D�m�@�]J��q��,9�}���(�H!1e��l��S��`��(� 9�r�����u/{S�$w�M4�t.�"�5�g�"���,�4�{HpFNhc�]�:;��6��C|�Y�G�� �7��K�kk�z��S���J�>'F!ZL��7��I�J��x�Q��;+ﺶ�]����/��^�� cv�k�����1��Ő>��É-Ü�1��s�@�Q�euoTu�U�~]z�	A3g�
�����O�jR�U��
�����1���!E�ɾ8򢐊�%��ͺ�6[�p�/i�z瀥���2]گ�;ZE�}�`�0�K7�@�u{���y�{t�E,/ �!�fP|\�,����}BH&3�����k7%%�HlM�Z�.Ǆ<��&�퀒(;4L �!#ql�"6Rǯ�Npw�����}c�cr5iXI�5��B���𾂀�����X�C��h�����@E��@J"�1�\�`7C��+�Za:�	k�M�;a�r	0��4�Zկ��zAhb�M����h���o�}��y�0L�Zz�W1i�O�'ܨ!�����޿p���Z9M��~�X��	
��mp�p�*��Г�yǭ} x��((�MP���F~95<<(�B�tϼq9�f������k��@����L �r��A?�&/z2��w�:"���Ԣ�h��@�a�U����ia��wTo���Q~�R��s���|7C���K۳K�����Z�/��\�k�+�8[灬�ũ�b~L�њ��
V�S�#�Am<m�����	�劜�JqO���by�|Zk7��t"-I9;���^>O���f�?DE��1Q3� �.���9ԞNx^j//O����<T�n�Ɯz��}���*{scn 2��&���	[$�m�����R>�mF����Oqx�o@<��,r���>��X��|&T�6�X�pݭzYâ�T�������o��R����D���*�{����;�h��|���A�"PCl�w�Io����!{Y���}𣒍�_�����y��E*�oQ�yU���=(��':�/͇I'w������~��[�Q�nq��;a���s�Yp�>{��S�QS<_�يă��!��_:D�g���������O���=�8�^����G���0��}F��o���Ѭ��gᚰ�ネ_�XI�l<�1���
PT�&��Z-2p3S1@_���:͝�GF���4-���O� �n>�Y��i�peIz��^yجY2l��[�uD0΀$�Ϝ3�3ӛ��Nr�N��z�������5�-�dC"+�	o~�}"��'�T�L���F�_�LN�Zn��<���VGǽ����n!�R5�[[A<��Atz�������������{[Q�1���Hb#�N�z?�Z��4?Tm�}�FThnCo)?@s�݉�AH��r�`$G��J�X����;f�0���ݏ
:�$LC��2�_�ۘ�kg��p���wS�ۑ`%)���X|Dߵ�/5ӬSJSWr�c���˳'�>���(�?W�?�#h�L��X����y�F���7VWv�S|���Z:g�v��{v�Q/�
�$�+c#�i���}5x��,���:��ȟ���
.;�^�+��AI|$�r-6_z�j-�2�55���	�D�t )�1�`Ê��;� FQHf�A�ʪ_��\�H�:� �W�8��kފ�6>���R�<k�U6�Vvc��(� 8M�J�ּ&��~�t�O�?��T�u�:#�A��a���8�M����gR8p�R�P.(c"@���"�&�T�A�U��_��s��3;�8�Qyٔ����^ڛAo&c������5^��^�_�`�Y�Nd�9�?�>��uQtq��Q�F~e^J@[|����̅�B�r�'�s`�u~"��*{�ׂԒ���/��] �@��P����!�*Iq���K�?�=�$n�e^_y�� ��V�����V'n�/@����h�}��`��%S�M�A8Q�FӍ�\U��o.�@��B�Q
ZB5����;�H��.ɤ6Q��=Ɔ�����yܨK
��mǳ*	�i��kmٙ�W��l8PmC�O�co]0&�V_ ��Kzh���Z�qL�F�pDi�'c� S3MaR�1��R�E����YN��0�bR�?T�>J'��е>�(ސ�v����\��d���d��l%T��!��&����n�I�˾��D�U�ǃ�ς%'Q�U�L����;��Ʉ�\��B�06tN����5�8;`�M7��e���n��ԣ�kN)��#�=�B� w��_�2"m}a�,c[rfhJZ�2�yZڇ��?]����G���^P���;[W�X��n�����8	�41��D�w��H]��s1"JǼI�ꃒ��1ϐ'��ºF*���hR�m�W8�s��.���!.��u�+����]��?�y>�Bg9���1�W�d�i��p���%D|lANi�p2�@��L�{�՞�c�n������(ipέ�Z���N�9�;����2��B޽�>mX����L�đ�51!�ub�A&�]*��K1�\�TU��P�s�^T�_�AM�V!h�'�x��Q���K��?���W�u�����ŗ�X,�[�6�/��Uζ��!�+&ڠʜ��z�<8����ʠ�>��ou����G���8I��_i��-N1���o #�	���M,T՗�
�M^�b鼊��M�u�lB��ٲ��(�X�ˣ�Ȃ��i�b��B��X-XA��O}��77=f#��1���Ky.�.
e��!*�.�a��UG��:Y��t�\l�!��.ba�K[�:��}�#!�Ue܍�U��^��B��`Н�K�T+����`rq�!0��Ņ"�d��c�E��p+�I����V �V��?�
�����Z�p�[MX�Ԙ�x�Z�aBqv�����/,X/y#�Nz�gD\&�uIj_R�O�z<EP���Wc|8C�ct���M��n��/�$V�Px����Ui�졪k�Q�֢"\S�i9�uRG����/�C\�M���B@�C$�p��S�NN)!�5�z�r����`�[��Y7z������ß"�0��!���?�����'_`*���9�)�,hdVt[�9,�N�[}��?06�\�i�9����[�N%�B=��������NpF�/���[^�	�BL��R�N7�����v��*z-a�N��Jŏ�ת*� �Aʇ�����b���2iw��m�;���\���Ak�+=��O���%��H�>٬���������V�7Ѡ��m)jW�"�p�V�z=Y�E��7�RZ3bE�#���2�ej��z�%��1q��Ԉ�zr`�4,>���7��W=W�ѡ���U��R��
�_��~�~�>�!�$��<�A>]�(`���Y��3�2�P��d�(���MK���Ț|���V�����>3FeO����/߯2��/� Z׺q�����"F��4�^QNP����ʈA�s���!ohΤ�%�G���M��{!������D�Ge�$5�~�����Y~L�Ń:/!�����^4�;����^��ıZ�p�(^d+�UK�e�1{Pgu��BPVjpә�dϨ�E=y(g$�B�ҠX�f/K"Mo���U�~�m�N��� �jנ��c	W �l���r��0�l8��L��c�����y<�qh�: ]6�ɏ�"FΌnK����j王�?�/ň�� �Z��4a#�zh�و��������~�8(A���ɾ14f�����s�l�?|�n.�C��s��|ّ�"oz���f׎<|�_�
��jƲ��Y�9--+Q�ر�9��Տ;Wgw7�A)̫�_�@C�0�������]�T-b�J]Ph���v�R�]�I5+�����^��8}�h��J<�9Z5�:� 5`���Y����<��$Q܄Zy�($����n1�q�C��n�Q�A_?��m¡[���LP�mI~�2^F����׊�S�?�%/ːa���_�
������
W9�������?��a�N��˿'�O�}H�������oO�)t�O��t��	0C������j&��{oBǃ�� �R˚�U:��3;�G�"\Ep�{�hE��ۊ�\����,k�*���v��Ǉ�t<�3�)�?��ħ;�*D-\��4I�z�}q�?���sT/��N�p�
~�T��\X.n�Q(���$�2�R��p�o.R}�O8��w��I-_�wRc<Gb�V��!�|�;]�o��;酫Ț�o����)���W5������I_f�Ks��7���q	2���U$#JlWu�!s���58���������o2�����m*;�D�9P���H�\"v������\�U�������+ɡ�V<#5�K����ؙ��A
�p}���>V�<�r��e����Erp����Pm�<�C@nEl����a~�X�TXK?<5�dFj(]x5	K��:��'�����`A׹�ʧ�y�	:�p	��i_1��AQ5J�NN&CKw&}�p�	o��7���TVu/Λ��#�t�Ȅ��<��v�^'�K�9��d��_��� .<�p���m�J����У[Ս��R/J~�"9�e;���� `�Zz�k��M��������מ-�{V>���''*���a0=:������U"a��K�-�s��Q/�A����
Px�r�q����6�A]���m%xy�x�`f�
��E��P1+�lBw��zN�L�f�����2��=&���o� D�~�̳U#H46�_i�5SyQ<���������LM:UD.f@>�!V<1j����d��Q����dr?�<;�6YQ��2�{j��{&8*��.Y�0�K�J��Z�<��`����iű�R�&Ҟ؛I#c�XIM\Ė0���g�ywKXu�%�]�"}���}2��r,J�|P(Ecb�w��R~��6�$3�s��-��k\�S���䳹U����>�Vw�%�0�N�"Q�؟�
#~X��<�Jy����kَ��D��ݛV�?fʔ֙&�Q�Y(	�S�����8b�L�_t?����3v���K6--���mv�`�C�#}#��`���W����:fma�靹W�'��|�Β�=��<���;"=pi�����m���X�|�yrJ3�7�"�X��g|Y��H�Cm�X6T{��C5�%��Yw�	|�L�U��!�����a˯�s�^VQ�E�t�)�"m�U!Ed�(T򰖐�{��h��F�(秆K=@E`k�'-�r�@sl�|���K� ���
\�[$DnH�-��ہ��-�;fK���&v�T���Ͻo:�\V~T�W�����WG5����}��3v�Jʥs98��ɫ_��)#���p�ٞD<��W��tQ
d�r��~Ri3^/���	9`��pL��!��C��k�Ѻ���>(ݞ��o�l8#�[�yfW��&R�_���?V�d��zߓ�O�T䁁�����
�,�XK�	��r1���p�֚�0g�7�^Ĥ@R)��.��V3�t��_~�KMd�
5q闠�{?�#�_#�D?~��������O�	�?%��i� 4;�?�Yl����|qF���6���t��,,�1�*�!�iP*a�����]�����hbj�r����8���D�F	���$�����LJ6���9m�|� y7E��T"x6����5����V~g6�2�/+�����tI���å?��v��WOL$�����D�NTB\>F�R����P�l�������q~���mvF��]�e�a��СlW�C��M9y���I�'J�ĝ���%��YA��a�鯣�o�\׎���G�6����H��lW�	���FF\(����x�+�����U[�uZ�Wo��.�f�3��W�F��j;�:��֣.�6���@l2K&|������б�������u��t����t����?-d:�)���p<�b{�h@���v5�mB��.��u9	�ĝ^��&����&GՙA����j\���o�$,���O`��El`�]kS=���:����ٮ9�hZw@��y\$� ��IV�n���4<��*Ò�ܝ������f��`g�¨z:tO�:[�=h�=9�I7�]�)��El、.��X�Y�+d�eS��d�==~�h\�3x=�֜�N�|��M����Y�s��Z�^�:��w	G���ڐ9��񒩍�nIBn�vcƣL�f�:�1�2���l*Ə��� 5��M�/����:V�+,�P�\$c�0ZMaܯ<��Zؐ���� ?C���u7�pOPG	"�����}h{����g�P+��+%g�]��k������N��9
/FzE�Vf�@�ЗLW����W)�4�v�`�҄�{!�J��|�׹��'�ZHȔ����5�[���[��UrR�tAMçWX�	1(<t���jbQ����!����i��'m�8����|A��12�,
�Du�VJ��(/&� ڨ�ǈ��`f#A�O��ǚ�mU�N`���`�N����ʴ�tB�b�}��v7GM�	�9?�� I�)�����D����P��b�E�]�>qw;���`�< .�����bN�p�ü� �(9��R�:�=��I����\dj�Fd��/��)�1,�ci�'d�VF5)ɐ�\Ȫ|q$Q�Z*$�%$ۜ���ޝ���dHX@��z��$j���ԝ=o%�Eq�i��M���ɫ�e|����������ߔXa��V���=��B���W���$�T����<�p�φ-�/���g?�CtSm�߼:A���z.{HR�=D=�8���{���}xq�|��:G��@(\�v�P���3�I��(�����F�p#:P���?�V��g����ۥ��W���Z�'��o[����~~Z��� 7V�:i�q���`�J>6��i���wN�z!_��)\'D�Zy�j�,5�~�X�&�d��Еfd�ح&�Td���q4Ə�y�|�������]��KF9���sn�0j�	�a�b]jL���R��M6r�����,N�����7�o����O�8���3�b��թ�$ �R�g&�G%c�:A٧�é~�Q�a6T^�+K��e��c��F�f���4�m�����8x[?+�ٟ��H���X�f�>��+��~T9�O�g��z�Z�9X�P�O��֦i�i�U�Y��y#X�oO*����چ�����bd{�S N1ٵ�R�m�ⲏc���Gc�x�^]L	(9o��횤z�P���LR�|b�
+��m��]@�Z3���T<�M*�*K��<�{���
@$ߨ��0��ƫyKm��{��fTޗ)PȻ��+�����奋�o��ɣs��sF��O9V���G�:/�z��D*�?O�8'�+�������9ǐ���9�Ѣ��¹	�����ӗC�2�����O��1�R .��֢�����.S{Ul�ho�{�G&v�6!�*�@2��s��5{)���YP�S��B!����q>�k��Xݼ�AQ8L��kz{�5$��mǚ�D?L����N���qܴ���f��t$L� ���5�4�k^���=W����8����h�(/�$s�O�lKp�%|�j���n��u��8٨��F.&GUK=X�	eU��iIO���d����D 1��~���KC��8�8c��$��G��	�L��nB7�}ßr�9�	�/?�=�g|x@��r�1;yj�G�K>�ݠ,�
T�{K�\ n m�]M��>i�,�(Ev�t4�H����:�q��QwBL��"�&7�)K��#z�C�u�N��F�[_�<9߁��t�Rb�Z�{*O�䬱+]Kx#$-(����r�"w������8{�
��X��1�Oi�7�
�q\�����c��Mtuj��.����2����gl��p]m ��
�J!��P�J�h�Y3��??5-�8����̔�V�.�������m�e��1+�p����ʦh�?7���܌�������J�,(*���4�|O�}�	R_�ܢ�4.«�j�H C�Ll��+,��sG�L5J�_6���cH��9jN��[���A�͗��@&����+t5h�zSP�ò	Z:�ec��McSj@*�"؁��~*Q��ީ|q ��~8L��b.�6�vM��T�[�q��gQ��q�^�>��V�Ҥ@��Y�?(�C�)����*�zG��ydQ���!�T-��"�G�gY�X�Y�d?�|(,�u�����X-^o�a#d(z�����|>�N��r?����`^�:�j�JO�_�'-��3��\���Z��4��	��ė�]&�Q�S���6�@���II��#�����y|�>C�|2��4�{���A��ǒ#�Jeܛ�P�O�����\؉Q�[�e;��ԫ�lqRU�"�	���52|��?Z�#��C���ҭ�ݳp�^���x�]��H>V>�R3ܳ���RO�w1_x���H�Zh����,��[��D�։�%�]§�BA�u�~\�u���Z�f>�W�<d0b�Q��[�y]_����{��djZD�����LR�𰴖$؁K>��	��k<�+}#��H@���1#�A�%I��3!�xY�5���D�ޥ]��e��X����
Xg��#��Qw��iӞD�r��j����?�$��u(��������W�L�Y+��#�mT�#�����"�W����*g����I+b�*�f��h��3�;���U�!��~�}�}��t쏡��0>^9;C-�؃�%�LZ��	�=�������5�����m���Kϳ�pM�n��[F�B����:��3U�1����i��Hi�#�`(���	���J>�xԕ!������A3�R��dݥx�KH;b�d�ָ>�&��M$JA����7Tu�%��j��t'�PJ_%��Σ5O��jD�l��'���J��ؼH0�o�<��Xl��U)���v<F9��!����uˁ�`Մ{�@J�.��K�έ+���cw��n,�Z�N���&OJ&�{2�����P��O���J��2e�=˪d��#��!�B�,�y�1Pૹ�yC/Ȟ�VǤ膽�~�=M��o�3�qU,b^_��ѓ����\�鼀b����&����N�L���v��j����[5s"��g2��'�81�nm@#_���`�}�G�����S����ՒCE񥺑E���.�����S@U���}�i�!�Ge����vlS!�qф��`������ ��L�z+��O�%�C��C���DJ�9@�8�Z<�/�JA�N��������bz8p/�/!�U<)�?<�@��E/�T���Kk�-�:e��V@O3"ʓ�_�LQ�4*�G�b�����3�������}�d���G�䈑�~��J�B"]�n�X+;۬��bp��x\L+�N��.���x���A}f��l1�#�MM���6RȒ~�I�l�>td����cORW�+e˧��ݚc�r�r���Χ������������+Y�;D����� ch���/*�Ng�����S�)y����o�4�H&,6���vQ"�^������^�Y"������HP���zS<ұ�d���G��p��G@-�ƕ�Q�rz�IH���a�tpt�4]@Cs쓨0�8Z�;�_�J�r�!�����P���F�6~�z5����LK�_g����?钊�%p�x�.�y�uڬ�g���<� �:x�+������t���!�w3x��D���)tI�ZwYP8�QkG���^�ٍ�|�`Su�����k�'(.�O�4_{I'&*>1`\ZL'�Ro �y�s��|��9��G���g���toV���Ak `G
�bR�+O��{vq�D285q�>�H�SJǀ�h�с
/�KY�tJ*�ǖ�k�k�L�u�����5(��4v����IO�:߰�O���� ڀ�6��#Z�$z����)���Ϗ�lz�5���`�M�+�r?):iR \�s�-��~mzf$P2�+�%��6��%<#�<�x�]�.���Y�i$�������(I>�-���@�=`qI�2��3����D^� 2���:��A4��A���)B�U��Z�df'TK����N�v=:�
���� r�YK:K�9��*��mʭd�LF�Q(�#5vm�b��q^h��":����f��	 ��j(�z�?k��H:m�}!�pM�N
hC_v|"b>3.���0���
��Xd�������	EO�BF���#O�����dC����* \���$�	q���n�l���1�D��(m���,T ��`"��た�u|�d���w M-����3�}���a)��
�s3ޑ�q��C��'�������'l���5b��Y^A���0o��D���i�V0!DV�]	����}|E��;h���]���.�U$H��e�q.�wtU���a %����"kO2��6Ӷ��v�F�^�C?
��3M�����$ɏ
r	��*���3؀�x�yTd[�n�4����榿a�KHϵ�@��3,�T�b��@�T��]�FR@M�(����O��m�����Ȱ\��$�O�Ǵ:P��n9Ϥ�h�p�8�jV����ˆ�0�Z2,��X�$W���:8&t���~�A~��X��Ts�p,.������F��&t�Ϛ<���ݞ��a��[�W��P��ɔ�LS��v����gɧ_