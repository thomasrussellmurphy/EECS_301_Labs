��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��/��Q�w���a5P��B�~�/�'̙���S{���^�qѝz��'�hřD~dVr�F�!5�=��[�\�bYzy��d�(5���*������j M����J����Cw&�u����Dg��>_�,��o��3�9=]�sn��5���A<�-��Y�,���AU�G���̻N�	�Ϩ�g�ϵ�w�Ω�k���R�9HO�o�u�(v�W�T�yVL �q^�Q�0/�����)1�cڵ�E
�W�D�t/�Ș���~x��R�X7�]0|��?ͭ�m׭��e��%\rN���H�i��8A(_�P��0];�ű
�0y�����
�F�(�}�����6�o
\�Tf�,d���b�$,d-�OƂ�^��seI�@����
���F��#Ru�F��Xϵ;h�oAv]ChQ���:����m��v+V�xV�W�Y)X��� m��wv���
�3�VRHO�-8�+����Rs �����c�C�������h�qb��6��ηd�<�:��P�Lz�2���E���{]ޚ"J�^�_~��x9�r4�\��D������%�.��u �iU���������.�Qiv�IG�2��v��K/�2!l׉w̫'�nS]>�)_
�op%���ku���BӴ��9,���HH��P�su�2V�W�M|ni�Ά+���HB�}qX��Mˬ%�`D/�`��>�=ꅌ4D�\s�°h��R��/87�D"���`,"�����9�
s��L�f� �]�R�G���6ǝʄW��R���(�ʦcW��(�?~i[fJߐ��<Y�I�ҙ��K<V(U�<�|ƽ7��x�j���)@V�HA�bj����iX�C�@};�!��ۘ��k.WKAh�Ԭ �g_��M�
r����=M�zA�ˊ@�����TѨ�i�4kدYt![�y$3�+�޺����c^-�R������L:�a��Z�����B�
�u�#�qt�",M����g$ F�ٱ�*��Ⱦ��0�Ps`��y��vN�j�&Q1E�4��Yڲ��J��S�n����*���q�G4SI\��w�[��@��U�8dp�3�)�u���1���x*�[�("���,|g�G5��q D����tI^��nK�0����b����n�Y�6�]��UP�|^y��a����^4�n�C�]d�E_?Ԡ���H��F���.gn�j��w��8���0{<�	v��Sm���h�v?S�@\x.�J��nư9Fx��Řg`́p��T�P��9�I)�E7����$�} �������=Ǹ���qf��O��	�PI��`�~B��c����
PEp#��퓰G1ء�hLgWN��RBJ��+d����/�m��Z.����Gy&P­�,/��I���i�W?�Y��)N��*�xB���o
עT:ڠ�50���]��`�Fd �Z�A�d�"NdK�_��l� _�p��n�2ƺ'N��9��S�CM7�L-I?��1Hg���n=����;t�}��r�DRϽ����{_�(F�� 7m�6UyC��^t�`퀃��"S��P���f�x˷�5OL�ۈP��U� �H�N����x��V�!�,C%�P2p�I?�B?�ȇI�T%�=�33��pd�o����\ƈ0�{MHXB3 �-�Ű��[��6i��b��蔽}T`��C�B� �4�B~���X
�^*�Ęd����ZM�-@�"g:��J�ޞ�$E᪮"�X�hٷ�/$���X��Kj���S�t�����cC�~�Y���j�[�����a2�$m�u�L=���V?
st�O.R�����]D6K�� o[(3� N~+�_Iu�a䢂�u1�D���;1^-鼙� ŽȜ���y��R�ogr�2Ŵ�^z�q?K����X��HF�N��}����-X�*`8�k�'GkEV>��y�N���L�ky��f!�e��)�I��,�c	�W�� 5F��5m�$X�2V��n(�H�ݲ��n�RQ)�00X����3@��T4�Q� �kQ�� hU a�s�2
�V15�׍�U��UE؋����*�$K�đ���E�xz�������vϦ6�9�r4���k����|^����љY=4�'!K])s��P�'_!-�W�E-ī�3����Ly5_3�T{>�Lf��F�Mu�D��u3A�FW�
B)
��h,Y���iX�mRS\X_{ӈܪ�B>�ڭ�����*�8C	p��0�Tn�s��A|b�t	�f"3k�3�6;�<1!&~f3" �y��R;C<T�� ������0��4�r!���YOSvN�k�7F�D� ��k�>i��Q���(Oۃ=���c�v��HXbYX�,1�$���E�e�ݳ��A114�v�_u��W�����dzs�f��5HC�ɸH-m �d�̬�k~Pbʍ�7��u:Q8U��6=�{��,� ��[��Gـ՗��lǸܵ������Q�Y�,���ۗs��{
߾���A�A����W�7���9N�����3�1�*M,�Ѓ5�-x\�$qۜB�@,�Y�4C�����/�^p^��b@l�9>vJ��L��d �EK��u&�3?�nRy^#�@%��A�Pf����I��+�fK+Yk.�&�d��k���1��؂�� ���y2b��TcI��Z���+8�晣3bj-��K�(&"�x��P���=$�щ�洞Z!Hn�y�����ħ�s9�<k���W� (�˼C:���a�M�nE�au0ϵ���~�rhţ�����)_1đ���ss�~$o��
��n���z�q�x@s�n�uMᜩ����zZu)��b�ie=J�#�%�DiS�˹:>[bqi�2��pe��d��Q�����7��� vwv�[Ӱ\Oi�,���G��D_m,��š"���7���y)�S8�vk"&�q�Gʛ�ɗ�q&���F |��$��v��#��Gcj�M|�	�Pr��)��O�8�
Wis��'YP�f�+Lb�+��MB;~Μ������ja�V;<j�4W��Fl̓P��t�[p�{VL�6e�vAj%_3SvB�cb�a|�W�����8�����Mu�"��N>��憲��b"E	DTHL4m���N� y���8�	�Z�4m{���)���@7%���k4���:�i�\���l�V�t|�Mg��ԇ�-{y���b�%�H�t�h8��&خ����'�JN�#gB\l#�y�!��d��}���A������>��'b?ШM��a��f[����釳�;O�&>Ox]�mD��(��Gy-�	/9#+b룘�b��R7��l�߅r��,���:���?�����_ѫ$&e(}(_8mW��F��3���Y�RV���ױ��|�)�g.K��������=���CvYk�}����ĥ��ȯ8�������������'�0�c8��t��+�-t��x��!��&3Z`̒��?��h��ZC���ҧ�~�}%�����IRI��x �7|��5�6������r�"��m�N�Q�(���y�!���r��4��;˒������ ���J��_ow�$M^7�i'�fT�B������
���I-G|�\&Ɔ�������؞��-�`���oW-B�����P4=�t�N$�RB��h䩈@R�Tn����� 9��_���x|C�q -8ʦS$	9�~	fr�L�jVXe�N<Ш>��p��0�:2;Q1ҳq���aG�Z��g(�O��c�=;�=��c!���S<��hڻ����BrY�D�uM�	-MC�0��Hm���a|Hy�Y2v���93��ӧ��u�+V���/qi���.3����b����f� ���?|��;�	)55����e��,����R*J��֒�3�%��GA��/6c�DD�l=A|ddX3�ႨG(GلiΊ܄�4:�LU�Ra�_�m(�e���]@�mY3?v�B�3A��p�A?lE(�t+DG�0�~k8UT>�+K9uQĄ�� ���Bp��ӯr�_b�c������4�B��So�� M��ȧ���փ~, b��5���<@q�4���\��:8�f���:�c5p�K
C�?�>��~�Չ؊"WhhE��^��>�|����,��5a8l�ӗwS�S4�.�zA�Xi�3��y����F"-A���"Oxc��p�l����C'a�)���m�J�Nr���9/������oJ��t:�ɠ&��e8)#��9u�~��`ʺ|�ߥW��wz��]m_��wD蔺/�Wܽ�J�"�$i�sy��d�.��bD]���-RDgT���$OT,4ҷ�T�:��������s�����	`@c�ռ�nmH)iWشXP䒬!��M`���Ӟ�-Š<�@��-������J���o ~�Mc�XxrĬO������������������#���}E˕�{�j|���p���d/�3
�<5:�wg�M����V:3"�L���u3c9l�{ܩ�6��έ��S���o���d�j'�� �i�o���WsJ͂.s��}�=�+sY�iM�1B�y~�$wA� ����S���C$��ᓽK��4M�d�Dݛڒ>}��K�S-�+�^<�x�=Ih��F��M	�RҜkXt TD�C������l'��Z��.���OɊ7��������ҧ� qE��fK!�os�
�%�6�P�3CY�=W������HҽHCe�g���4�3�\�*Ua�?�����1�$o���ځL^�	�L�D'�
��U
㯼��q�F�1^�P#�^SJFfK��L�"��,z�<�Э�U9��Y���߇C����5Ol�fԕ �`9��5�?ކ�����+4���y�LÖ]�n5�D{��`&ϗ<Z���̚��w�#�߇��kb.D�r��?~�u�C���C)�F���/+=t�vl%^�#��{��3݇���[�&�lJ�<��҂���?Xj����@��}{6oD^x3{�M{K�}8���b�o�n�X�$EC֭��c'���F��>X���`{�����aY�CO��u
��ku���-q��5S��^VV�`���c+�q Q=��$C��C;�X;J�W����#<��e��J`7��xn߯+7�n��ɰ����d��+����4�v��`&z��zG�3��b��g�U����lF����gw�r��P�{E�r�x��N��%�t%6M�#;an]#��$_��ϸf��o�8o�mpZ��@�$7`Er¦ŋO�K�,/�u8*Y˰D���>�gXh�{-�{Y���J��(|r�v�#;�A�2!���Y�>p��M�����)�)�$�;c�g�����=i;��={԰�Ya�����a2�.�ޤ|�*��
0D����HT��t��&���-)g,�썢�jq"�Tb�U��j4�.� 	�Z�|��8��x_�5����ق&�_Z	��Y�㱙�KRYd�v/H۲����Tp!O�_�A4�92v��=��.�Up�^��fl�0O����ߔ�0��B�9P��7�4�|�����\�H(�G�K��Xu]�7�a��c�`�U��� }^@��a�k�����t��jp���L�81�f��}�Y=��-�6����|�Ш��,�W '������C]��yJ'ǟY:0���eYZBwA�%��S-V턙��׭0cC.]����{^!�M;�K����E�5H��:2cM"C�t
uxi��|���n���(_-v�,�������h�sX�Rϧ���%�VX���ǒ�������j���ⳃ�lV�m�S,/�2�}s�
*-H;p�h5�������\���>O0y̏�<s��?��u��?<Y�ǯ�.���`u�yHy�%S��8s�5�'�L���L�)*b�R�ۃ~\��-�.'�M[�b�O/�'@�i��n̙�*p@`����
)3��N�W�\�C�(�;�ʱ�����e�)�����B��T������O�R!r�*\���U/��njwhF��D8��/r���%�4��j�l
	�)�Y���l�k��g!w��9�Y�$����z��c@8� 1YJ�h��,U	T��n5�fQ�+o���M�J<��Y��Ѐ@F�s�-g�F=Ng<�G�C	�r��&=7E�*n.b~O�.����PZD�u�z)��[�X�B����Ɵ��7���J��W�(}V���h�!��J6%h:.�#��c^P�d�d�C��2��D�z?�JXA �B2_��_P��z�f �ꚫ��[$��{/�@(qf���ƨ1W�W�TR�@� ���4t�ȟq+v-���p%uf�\Y���\��6��M�/��co?���?��K V����G��ěb�(�6�K�֦�7k;�hQ��d��΃O:rBXQb��$;6�epPf����dV�,��#>v�5N���	uz�́�"&�nA�Ȁy�{������q�"�
+
�GZV���@��v�l�&�5�P���,�Y�@g�`���G|v�/�xT&>���x�e�~=��lڣ�y�g�"�E��\�}q�'��	��������`H�l�7lDם3�5*GF��-���L!�i	��2�(�����Σ��%	���`|��esׂ!N��ú�$1��7Wo�����c�|�ˉ�v<M��39�t�qA��h�|8�a�1&�>	9c~���b!���?��G���#�3U5����r�]��ݓW8��@P�q8[L�|3_r�3aK��ă��xG���V}�=���F����׶�lر+0��rp9��r�n+�W�2���!�鏽��ŉ��i�y�9����Y4[`vʝ�W����,�8!���(j�5g=��w���?:K�F��M�IWt��<�y�c������Eʪ�v.$��m� �oQ�d���(W	�����[f�t"���3�GǂUUY�ԃܼ�J�_,�j]2��R`iXm}����F�!@�y�)�A�k|����v>�02����LXhO(�R��l��{�=2E�9��魑��C���K����A98G$�<�\P<��fvq�s�A���Ŵ@�ժ�XO�qi�<~o�aS/5X�n��d�X�3�f��`~|}Q`��@ӾnY}�f)h`��* so�A��A�ĆL���yc�v�ή�W.)1�[�i�#% ����������Y�T��c�����)�r���Mh	=u������Ǵĥ� )�s���,p��l��-j��G����/���JwF�.J�:�����6�-�~��W����`�cvU$7��㵘��7P��edF�Xž���W���O��X��R�- �CJ���vɵJ��|TZ�F${p����11ŸI��q��Йqi�H�R�}D||�̛��VAUq:�{\MǊ��3A�r#6.������r^��lh�X�"���^���Y��`)2  ���������u�یgʲ�*��p�;�c����w��H�h���$pim8�V"�����}�E5훥Қ,������^v���$��9<�c�X��G�q��@��G*
�3N۵B`��C��A�Jc����,��~Z9?�©T����l�pm�����2��x�4d|�)y�B{S8�]�F�x�A�Ǒǧ{�r���a��)/��/��>�`颶�T�`Le*�?�t�w�_� ���x��$�8���������A����^��7��Ym�3GP��˳�gyϥ̩�Y��z�,���]%�3u�JI���Pu,�Fn��Z9m��-F�b�RԀ(�&���hC�%�yu�J��@�ȴB3;_ �@\��H?X��tZ���1Fתf�>a��J�t$PfמFo/,kUݙ�@B�R�XYFH%q�d�
:>1HD��̇�#X��������eIw���kgjN��q�.if�<'�W�z���l��F�m&��2�49�	����&�,"���p%�{V�
�=���rև(�\�3!=�R��(��O���������lj����;����_���'�*����C�u���W6���� +,���a����L��D�����c�.>@��r�:w��oCѶ��'��`��ש��������n�"����9Ÿ�F�L����J��B�i�Q_Y6w��'���{��iR�h%����1����a��#F2PIΑՉ{N�ȅ'b;;��Z:}5��?(�*N�?�,*�̀�Dא�@a�[4�w1�ĉ�-�̔��h���HS3� VP���T��\��	l���!��*оG+�'fkI��T��͟�L�Ǽ %W9e?�z�}bGNB�L֥v�h_X�GuаD�3�q0���-��U�b�ṯ�!�r`�q�#��YT�<���|~��5�lz�@��#E��}Ϻ�q-����<TOZ�gg����K,M7��$��
{�S��dI�gkX[�p�]?A���IT2�$ͩL��e�"͙�%�H����A?[��r�D��^'�m~��5!��i+�Y�U�YI�UyY�F��ҽ9��6B�o|���#��$��tw)l$���v%�j���K��,z'[���Г_�e�&�3���:oC�z�~�Ao._�J�qu�R�[����':$lD:Q�a֐�+�F���o��r��f��U~xQ<p�b����3���A��XO��R��'�X�s3�7�1.u�^}�3����1Z���ɓ��-��r��5�96kr� _�F�"Gt
�IQL;��Zj<l�*vP�����<G����9���6�v5*+9͘��/;����T���alA%lF_�!d����r+6��Ss;�E!�H(�"�0�@��&�q{0�:��������`���PTF�Jh����9x�Sh9mK8l���<��_F�b��eZ?��7b�Q7�vxXP}A�dZ��u��I�Z^�M�*YK�@�-�������0sN�?�ч�1�c����X=h�f=��dL�Q��~)� g�����lNaˆ}
/Y��Gr&Z�Z0L�.���m{XvrKâIe�i]���.�Uq�d�<A#������D���ٽZ��-i�'g���Â6x��B����I�V���q�y��:qf��;�{��x0�S�L��}"���N�G��/�51E�6�7M8LNIR$��q�6��CP�?�{l|��_���/;�f}j��J�`�1��Bm�P��>`p�,��<K��Cw�������w䖄4('V����cc������|��&�c���l�,�d64$Q��y�A�2��K���r�a���ȿ/�,��Q����N�BCR���
0�a��G�Z��ZpW�BMDSb��3FDUX�����ܻ�v?#����W�-z���"�㕍���jk�Y0�&;{�h�:^�b�O��WI�9}�a8Ir��"p�{����i�<���P0,���L�]�^�)�T]��Dz���tۛ��-у?5'w^{yE� yZ��>a=��1��ח�DԨ�3�z��^����n{XT�Z!F�S�U+<	_Mq~x��l�r��}Y����7V��5!+�|y�#�AA�uC��Ɣ�i;��٘�6s��$���%���� ��1R��aX�^��������Z���+�|�ی��~�Ki'��ٗ�|��z�.�`w������2�X�L����b�K]��v�m��/O!�����a܊�'Oh5׿�xݼA*�r+�*�/�Zwօ�`SEtl��>ALg�**�Z
��o�U�3ap�t�C����[L�U+��ml� ���:Bݝ�V����⋃�NPr���b�t�^{m)V����N��gf��U�Ց�1���оp�	������J��m��v_�:5��;J
,���P�}m���m�i�ڟ'���uQ��ﳁ �3��;����5����>!:� y��uTH�$7��/��Y��ztOqdS���܌�2���$0�5IS�Է����u@R7n�SO߹O���s�򲜂F*=������a�����<�g$o�_�?�S������Xh�o���~�6'�Ha;��9�ÙJk_w�����%���jnЊ���|E9
�vm�9᪀E���K�d70�x��OD�-Ǉ�n1 �r��6]�7/*���	R^19>�@K��
k�]��ô������:z;�������)��Ґ?�~�{�����!Q
Q�$�P�{!��aat�e��jFU�����+���D���b��̷&hb4���A�=����=��b�CN��H�U)��:�¾O#ʫo*�\mڐ�psn<�p3�jـ��w��s��!�𺔾k��v��� �>��!mrT��\��^\�i�����>�2�s�s�=/����l,̣6���p~Y Y6�JB#L�L}�I�,|5O�d��)��
�T`�Q<�[KEǲ��H�z��ڦ�#��g���`�	>J�n�/��PB5ۡ�}���:�H�6��)���LF���s���!W��:`+[`.` �ۈ ���\[���^J�->����ol�~v;�g���wVf�ۊ���ulP�Z|���y�<�	+7v�8�ټg�畏I������'b����a�]V��q��E}�;CۼW�]s襯��1�߷$i�W}EE&Ϸ'R���k��%o����1�LV<rn,��ÏcS�.�bu~(Vg��U�2�����~�N��JMed��I��>G<���rp�Q@�C-6N�7�� �A�v�{=;�걃�%g�2`IPic����"�E��v���M_h4��/�]4:(��'#���c�y		z��$��qiEh�tHa�H��C'"��$�֒T���
w1����7/�㮷~".ش����v7��_^�/�
�%ٯ�\����;�eW��i�;��1C�I�����㓣r8@4�mb@����T�_&��Q��Z~J�r���Ѝ$�7u��46��Av�T'Fi����%�
�i��}vyWڍwJ�i���Ew9��e=EY�P6ۤ	�7i�t�@c2Q%fR*<�/���U������l[`&EiVC�I������f��$�[m��4P�+���V�ݫƣ�]���q�z���>�8��N�;M�=���2'v_0�u�����qі�S�Z0t�\�"+vS�_3:�9������D㳗���B��e�0ve����5Q0�s�g~�tX'0�ʱ���:T�+�.*�ݮ��jh��H�C�^�.��&�E���񼚷�Q�DD�����y������� X9~��*�V(Qe}b�F��%��Y�"]Awk��z~������=�K��5�u�V_�����%�R%�ln���зt�FPkS�>��dƖ�H��v�9 ��+�_rӭ�1��uK����[��:�����β>n��C�^�q(D(���H5�������i����ۦe�Th�;\�f�EDQ?(��t2��l�U rf�n�x|����QNX��y�й�c���CwL�m�.�X����{����������HB��:ԍy�*�TA���*�n�T��=��х��g���׃W�۰��$DH�6?����-�W̳�ъ߂�s�
��e�7���Az�R���=�(�Y�Ë��AJ�+[��Y'6r����{.��Q]JF�A���rDԆo�^ޕ�ݽ�Q���t3��p,gu��e�2�YLp�!���l����/r*m�?��~r��n�$��թچ�+�#�,�V
-DT��>ڛD������:*I&Q�A�{#j���&"/�	�~H� ����� :5�����yu�Mb��R7��i�a�I��yT�6�(d��� �g8\�lDI6�CQ3b��W��㿯����'�X��̞���+�ԦT�Xa�yC���x5��n吹�+Y�Θ"ȓ�W��y�#j�y]��n&�"�Q^��23�I��]�;��_���!�d(i�:*��x��#�o5:�Z٠C#O�:b~ԁ)���H[��yL��	��H��|ufcJ!��ֿ8�F��y�ˋ*ڀ~������y�n�)_�a����V�QUOP���T��w���i�?�}�~����/�ж%�u�V*sy&^HI>�_7�U���:��Ԃ�n����A�]ο�ם���ȻX*����9����}��o�-��{v�/󰫆�G�5v3��dٯӗ���2�g�#�9u�ηE�X�lN�P`
q�I�y�I}�8��<W�Eq��)��<�g�Z��r������Xb7�����~��旀]�f��3]n$ry(=��6s���"`Y�=i����m1��1�^ʣBT�m��:��"�āj�|<��C�dۮ���^T�~�{g�M�z�ٟy�gR�����Gf��M~�����YeGtwW���k��}�?���mtĆn
̛�I��]=#(fE��8�B��j���+�l�\E�8�%���$smr���SH�h^�V��&�z%�Ȼp�wMuN$2�j�'8��M��m�d^o�;�[W@AT'ui�~oP��q�6w���A<R��j�+���ȼ�9�
!%}J8�
���N�`�i��A�R�l�a�%����z���W�Bc�Cл��c��n�;-'�SB5���U1�W߆E�K�,5 �H�E�h0m&+)�=)������iU�~n���1��E�o__Jrb��]�N� A	X�~�
J��J
uN�.`�=#��w}^�#_����/4g���'6�ea�������N)${ˏ�L�xH)�;Re�8o�qO	Տ4��PSs  �pDuzI��`]a@2��e�ju<����8|B�%A�%�z��f�T��~��=�+aB5cȿ�\8r&5,��d�z쮥WoH0!��x6̀�F�t8�8�oAp����M�,?:�ə�_?^���1�v�����@�nE� ��8LF�Uŵ\:���T�Fw�~�"L]�R���Ƞ��b���F�yqp��;���CE�����C>_BΫ�� >?��M��?���&�H��eS�E��9����m��g :��AM&���0�aQ[c�#������S�m�-02�d��#z�^��ͥ���9z\̐$�����p���F0���U� i͛��e:��&o&Ufl�����rB�\n�+Fp���V
��[|��c���XL�١��xʦ�6��F�!"ن+����^S�1���G��d�Q�l�P��OŒKi�����8�lf=��rM�#��g��Pf�v��OR겎���y,ښ��!�	�S�[Y���@�c�K]�W�ӑ�+\�炨V+�Y�z�>Z��_q*Q}�С}�?KD�[	�(G����9v��R�8��.W< O��V�N���t}��sʸ��|��2��H�=n����UD���0n	@�q���m'!���4�,8&�{!r~��Jua�%��%Ei��_
��e&۠�x&`�@ �g2��c9�U��%���}M�����NB`�a���ab$��*Pdd�����f>yu��q��Z��fސFꜴ$V�8��ŌLB�^ s��@-�`EOJH'� ��_�ޕ����L��ת�uD7��ͬ�0�q���~+|����k����� �!�E���L~���Y���V�����gl4]��&�p��zDIܒ� e�4�GN)�pc��g�B�;��������Y�AN��������4W���D�P�Ա������ �RB�Z�[�E1�<�C��!�)��٧YX[�.{Sh�2�w�8_&$�A�&���9v"
lЃj���tP���X+��p���'��XZh60o��R�1�Lb�+���[�b��u�!��^��f�� �ݛ5���S�h�ً���%҉Z:vs��W�Pμd����7�"�y���|�g��~PW���$��u�Sb�jJ�O���[�UC��Of�u�=OK�5�Ϳߠ������do��6|g�����E۟}��C�=_M*;߯e�� ��O�}���_����]}�2L�r���D�d�*l�R�'��.ꯅ�J�ꪝ����$@p�|Q����%L����9��-f�!�q�p#ʞ�R�!2>l���ݛM,���-
���+��Ѥ2�'�@1֥�L����9 @9Bѥ�AqkƗ�{c�ZxK��r���m�z��~EJ�0%����Ի+}6H���sYk�e���E�Ty���26�
N������~`���2�k��j-H\�'csK���EL�|��)+��J(��[������5fgrp���`=t]0�(�lX>�C�Z�DoƘ.���C$#�a�x�����a����)��*\q�C���95�Y�3�/5C�+�l�����	��V�M��K:�ުu�I)9@���j���Y�	!ng�*3���!.�����a�aƞ��K����I���2aL����v�ƗYl�?�?�#˼'T�a�=XM�͋��鰴D$�U-K��eD4��]e��7u�A��C����S>u�3\�w$g��RyN�p���~���n�YU�����W�n������rN��[��`����1y��"!vDK�#�OM�⏥ᗍ!33��{�_���D�����:�l����%)��BH��7ܪ�G��n+�LF��x���m5�͑���#�uOӖ�Z��̏f9僛r#�L2�T�tꆢ����y2��P#�"0[%�¶�R��!��
�U�h�WY��Y��.5n�"V6ۀ�J������I���yon<������P�������Ԩ�ӿ�{L	5�Ts��	|��4��E9�z�^� ��9�E��)Vm�:%�k5�mv���w��"�x����矦9_	�qn	��T�������L�ИBy�!0�)��MÀ�#~��&Q��ɭ��;Q��Q&a_�y��)?4d:B��(|����޹Akd����c�����������f���%�����U�p��5_-��_s�S3Z����=��sx2��O��Ye/DV�Ģ&���zv�iY�������Jb�c��&�=�q֧ϱ�<NumDj�^�4���qJ_�T��9g��f�!���O5w^�9>:�k�܆8[
��qh��%"�<��73�h��F�I
g/8z�!�ط�zkX5���۵o�dh��	�f:�w�IO���[_��V��NH�y�J���
r���*I[(� �W�>�x�DA���gF=��U����/ Ed*�6+��#�K�BZ`P�;O����f��mh�ѵ�E���4|%��&x�Ð;�B��}�t�#��K_f��)����joGU�̫q�
�5m����+V���0%f�<�E���"��F�0��TZ
�8�/x	�_��)����R<b6�z̥e�nf�j�j~�Fx�(*/�3����Ȇ�nf�M���rA� E/g�P�S-��n�X��b����"m!�c��x�	��㊰��C�)?/��Cָ����w>`xK���P-�]D��|�2�T��ѡ��]�@��B-�ۨ��I.F�e�&l�^p2�5��ʱ���p���B�N�3mf��ofx���MmV��-��q~����6us!�XR�q��N�!"������zGӭ��x�:c�u�ڻ�U�=x��e}�����݁𴧴FJ���!���6l�>�a�-���/�&� ��pQ}�rIË�]w�Q�i��yS�.�����˖\O-a��������e��@ݘ����� �V=�NArR��#E�H��i���0��7A�ߏΪ���N9s)�.���]ە��	�	e��y8��>�_kX��>���l��9��Y� `��eb��I$�B�������+!�*�~,;��f-S�韜Үn01�ϴ����������QL���#=�@(0M^�@:r�a�(�?#�N����X$��	\Nn��`H�ȍ��~a�,���u��|�w������[I-H4r�럹ɾa��R����a��=So� k F�
%�◒����R���{������dEI���c�G�������p�K!��N���rpȈ��J�E���
� �|�$���	�Yvx)��?~T$RU8�ܸ<�I-��Zt�E:����k�&�]�l�^��TT^����T�Ʒ\��s�*�[5\�U�vi�Y�l��}��Z�V��u���{��)	���"����rmW��py70�<~�>�zD+x��د4l��]V@��{*Hy.[�?.�	�q�gZ}ڔT�^P�6� ��x�ד��v�=��U���P`d��͒^��Z��j�L
O�a: �����3�~w�ۻ��N����^X`�?�ĉ�����(��B>XKЄ~��'B�@���w��.?W����Z�&/�~����{��6��㹐ZDy|�Z"�b��Yp���T��KZ�:C�@���f��̹%�<+�g5}%\���!�
ߖJ>g� 7{A���x�gd�)b���.��Y$\�*$�%���n�D}��P?$��;�.����ZZ={K�wtL�����Z�ͷ3�\\tl�b`�U�r0e�/%=�w\E�~M�������4�/���X���<}�8�Њ�'�וL�.:v.) ��NP�/�~�K�>���C���-^�Fo�=��D)�I9G���Z3
��.ͣ�p(i����p�;�5H���⹭�"�6��8���'0���}b���š����T����wڈoOm� ��'O�H'�F܅�+�.Pl{�x���s���mK�G��
�'~���+Ig*+����R#"�a)�B/:L��b��o�S��@�1��-��B�D�aݧ�"�Lu�8�f��4�ս��1W\����O��" ���%f%kb0kjy͌uN�_D
n�CF�#<��̋��Tn*$��+D��12إ�SPj�}r�2�M�<G��Wy���ᭆ1�hm���}d�7�
�^C,��f��槥A �3灋k!��pW{r_����Zc�A�WI\��z��T�OwO���0;?h����U	��ϛg/�f=����g�)Z����Ꙛ�Uh	����z(拜 �]qk4V2������Bܜ���ʵ��ѡ�f=�jG3���L�A�pxC\�I<"�"��dga�����l�s ���39ǽ�w�j�mVv����]�O���)(��Z5���#���)�y%�	Q��܈����C�t���3J�j�����N�pE۠���Zy�x �$�:,P
�L<7�8ד5ݼ!Mi�"�Ч��}Ԡ�q���v43�ҋ������m�X�y���Ӝ�H|�3kJ�1n_n�����m�@BNJlHQ�Q�:[���L�F��wDr뜽�?M���+L>���W8<��xX�w�5/�"��-�:EOp�������M�wV�w��Z^��y���/�fk���{Ӑ�n��vE����LZ�S�u��I�p�]�N�\�L_t6@�-Tcc�նl�"����v����'}P���1��N�H�ѵ��[6��-n%?��i
WL��O���L7�E�R/:���m����X�!	��hX��O��/�N�6|IJ�+ƫ�䫨���0W'��L����k��T����<���]țl�e���h=�C�?j'��	�1kPC���%L3B�,f>��+���^=��/(�?��A�,�x�6�^��B�6f,	}�z� ������q�c���*M�vr�aۑ��_t�
�&W��9����D���D}X�|p�.孨��%k=��1�N�� �����5�I�F�w��v-��fp��U�yoǮ��e(����r(����V���X��h���!5Z�&/�|_L6�h'OJpz$�J� �/X���#��R�e�K�%��J��xH�v7���V Gũ����P�(�d,,�<������p���;����z�̴e�!�������������jz(Ī?�*5�ڒ-�6&���+�Ev�H �h�����>q�~��:'�<�]
��>��g{ɣA6BK�Hh!>����e�LU\zȽT�O�uƜ�,��dV}m���Z��"�����Y�g15�9I{Rn�x6�'�`���;�X�g�%y�_+Y�o��1pԓ��Q�1>k�F�n�f��lɹ���Oj�v/!�*uIɖ�M��(�݅^x��w{���/):2oVbǴ�~=�wqIS���M04���]j��?��e�5)P���=^󠮡�L����*�@ڑd�0���ea�ᣚĮ-�V�p��t�q#�P_���R�$C�ſlvTLh�2��}�"���}���Q�IW�`��-�(%�� ��(7��F-A�O&���"iW>�L��Mh����ߪ�ޢ۷�]�������F4eTN���g<�zE���N�`���jt�$�ύ�HLYGg��Q4
)E�AgV1H}J뿄�Өb>b��VL�$˅���u4&�^t��y�ї�"�|A�pe��<���9�X{�KZ�o�Z��A�ȁŭ����bz�NB��ۈ����i����C7����h���n=N��	�/C|B�4W.�Z����;�9l��sӗ��_�l�X��H��|V�� ��Elh���`�cl�No|�n�X��/x�l�lH(Z��8�)���.:=i���(ͪ�j��>�@��0�j�χU5$ �#nׁ��L)Zl[�p�O��=���:�"���5K
d�|�F��#jQ$[�Q�ժ�0Z#��<\�1�w2��G葂3�'���:,:6��
��/W�����J���ł��C������=�/2��}��iV�W��W��'�d��3�[u~���R�|/������$��MJV}=������H-���2���W�ItBo��0�8��h��m楌�ϛ�+uP�j�v��ڱ͎����a��ڂw�W�0Kd�~^�����]566�Ͷ��#��Ϧ��	*G�'P �'%� ���tL��ˡܿ`�� k�OP����T�ӎ��D�+��Sp͸	hgW��c:��e��t l��w`wޘc�]\��fm$!{Q���F���J��?�:Wm�b�{�7�������"-_�WB���Tv�#�����V��{@���!N�E���\�1��"��~�|c񰄶� ��0J��oɮ���0[�lS�\����������$v��� ����2ՙu����z/��(gTM{�bؤ$ͷn��7��oɟnǘ��'�'E�����!ˆ>ݩ.��18^a.���w���-X��uV�KC>+��P�h��������riO�i�:�}
��r� ���X��u}[�]q
�V�y� �������u���͞	�S�d|�r��=�&�z-PYT��"�f	U�b�\��)�Z����+_�W�zc�(�!���|.j� ��tח�g!F��|b�`�a��<���hz��sI�iV-x��=�Qd���捱R4Yo�r��5�������[,p�	�1�.�S.�Ղ�������o�s��0������
���˃�e�B`�
 ]�0�ؓ�C}IaoqrgI؃�
��]" ���J-���k����+��q��!}�B���P��������%��)��eH`�e<�%���%V�B�x�����F��&�<��9��S���C2��P9�M�)��'�2����Krt��ϜPm�L�t@��:�N|c#�X`��~$��Dy�XD���u�V�r�ɝ�̠�?�|�G�k��Z4ܸ/�o�����M��=��;��0_�~t��P�v��b��C��+����.��"��z�k�0Ŏ��!�9��{�J���I���m��:k�m�LB�Xb]��P8�ﮤhS���sf���Ta�*d����l�_'���*,�=�+tv��w��Y���
<U	��`%���p��_����g��Y[^Q�y���%��)�;~�X+w��nj���.%T���Nt�а�����*�}#t4�lVT ʙC�4IL�1�]�p��7����˝�F��DO�&�?q�s;$~'�):�9,U�%5�	Uk��_��H��	�i�ɋ\"�O�ge�B`���N���*��#'��|2={^�k_��>e���u����PH0�����>+R�ћ�����
1��m��L�ȳ6��r��p����'��F �@3��bz�oץ����1d&`/���=~qbB3�T�#+��d�!��ȟl�,�'r2����U�f�o���	2���)s�!�J�Ѵ�����ro;�¿�JaE�!j])L�Y����Fj߇�-�0%q��A��w5�|��Q���Dy�dM
V���_5L�2� ���~�zU���0M�ǌ��������V|$�v)'��A"��.�*��oo#��Ҟ�o�����/�Zs�ˡ����'�%}��[���S�&lb/��y������+|N@��Zz߿��+}m(���u���n�JUB1����}tΌc=hf���ʹ](��B+�,u�u�:PC��|s��Օ���#hA0��:�=�q��5u[��f��;�ӌ��#5���m��؋*{��p�����|�&��8��?��ϺE��#�{���[w�P��f�0<�_[e�#	��
x�fc)3l��4[:nw11��峠}����h�*�������MߨA�ѩ�9Ԋ �5�綟#W!�8�m���xC���'D �ݾd����B59�^l�\�A�bgz��F�`=,X�t�_�����{.o4�Q���0y��8��2�&8����>���s�r�m�"u����̔ �|��i��$ 8���������<KeovK��"` �"����i~�ࢸE�|R��[Z����T�"R����ʌ���RKH"t,<������z-j���=�����.�Ҵ-`r2�KD򉂁\�U����b��;Y,2t�!w�Ia8K�<W.��|f nm�g�඙��X1��Ї�T�,Ad��KBUZ}����R�pu� ς��g�����V�Zh粲��D+A�����W:P��v82݇m���i/*Y�}�����O,����0T�\_�|7��{���+<��}�F���(*v^O��V���џ�����wk�k/���h5�j���IƯ��8,��+8ɀ^�
A������/���ܻ��4�����˟���g�]�٧�#|���e���P ~t�W�vI���Jٞ�?)x�
ڤ/#b�xP����Q>~���H��R4<8��;���C�z�?��m/����I��q(�gtg̋�Isa�{��p��^�nt;<�w�t�j*.��y(*l�nz���L�6���~ۯSl��}O��U�J֭L{6/A�0����I�'AJ��R϶��>�J��W����/�=.Fp][W�f��Ʃj�D7�������?� ܉���Ef7��N4��C�ӋϺ�D�fo�����WLiүyVQ��!r:[��,�F�r;E��P<��bDB;��H������|d<�Ju�:� ]E�{���M7��3e��~@K�Znw�G�A�G- �~I�&Oi%�n�-��l��V���eė�1��\��O=�3T|D�q��!1�}�@J���V�wg7g;{�h�N���7�E�y����
�l	���M2k�V¨�Cߩ��s��,e�!�A��
yS�zgY^j�&����2
e��0@��LÅ_p7$��,�I&u�5v��X�{3d`� 4*�����_!��d"׵� ��yE��'F��(��0�I����d
ZH�=�ݷxla��R���|Z�睊�XB33���S��ߔY�8%e98[�|F���Ylv�vp��X��{ w��ȳ;��� �Hđ~V���ⶤH�*g�^MS�,=��X�mr�#��6���2|~�������t�7�h~�����zA��1�� �Q+����Z���_��LJF��j/�Nw�p^V�K�e)��澤,�҆��Z�s�M�iB9VC$H�[m��n��%ڢ/�Tu��!&��KF����Vk�E`��o_^?Pg�Q�!���7L���ܘ�R�9��C�F�,j�{��#i��+�h��W�LǞ�
�s�Ã�.�]�lSw�a��5�Ԝ�>\2��m,9f�9���������@ߧ����9e�mA�r!��B?�l*�e��Ca(B�Y%�*w����P�}�^n�&	h=����@Iڨ�d�g��:h��m\�% ���$Ⱥ�o���	9|pΟTc�2Y�'�̆j�G����׆muY�{��"nݝ�U�p^C�qIJyEJ����'J[ː��������#=�+�� Y֢~7��
̞��<��Y��.Qw�<�U%��Ng�v9<\����T�n^���/W��ͺ���$������q��[�C�mU�_	�0�j�%,�@�z�e4O�Al�4��Rw"as�6���F�$é�u|n�r^�X����M��w;R�%8t��lɳT�#��6LM�L�<zs Of�{�g�5+���p�P^Q���<!�)����5��UـJ�*Q5��|DVq��Q�~e�9��z�@6�M&id���hkw�s��ߊ��ZM9t�y: ��ޏe��^��|x��=�)4k��V_���$��?P���@��Ul��~�"�K��b���'YQ���6��O����uV䆁$��fc<o@�6.�$¬�
gI�_�±�o(����rŞ��!�P	��
ǠɷS�^B;lRH;��鵑�v����o����k�n�M[�z�Q�a	�Xv��q]�e�y�m~c��AR������w���f�c�_}D�0�Ph�������e���NHE	:�*c�c�%����2\��6�bdtf�!a�X(X�'=yH���l��%h�D��1i=�e�RA��ӟ�E~'�!BI���Mg�6�n�U��û��_pѢ�����5��w�D��od:�WMJ9l�u��m�jTؠ�>
��x��X[Tr���Ȝ��t��tݎ�T�Bи�.�粻ر�$S�t�(������V�ߡ��_��q�,c�*.9QLc'�ȼ�Q�Vݟ��}xy�����|�/�N�>����g'T\2�ht��zQb5�5�{�Z �g�4J��a�AF��ĥ��?���F}i��HqL�i΃�>k�#����H�L+���p
�w�gT<�i�
;�w�-�|�xW���
	Ǘ����S�1�(�Oa[-�bf�"��(*�����,7J��c4"��>�v)�![5,��X2��C``�/�b�����L\��T�-��$"+���M��S���C'�c�%�Ap�'��̗C'"��H-�t��k�&iE d	��vZ�����'�K����H;��W1'�mi�qc�ZB�ը���z�x�!]����'>X$}�&s��� _	Q���5���Ѵ|���?Z�3�YK֠7S�U�����@���s}<��({���#l��ݶ:�A�5?���q�r��zH�e2�x�������G�����ً%{��^=�Q�G�T�粕`]w�n�v���t�/bs�v�k�FU��]��X�m��s�rTf�+?`�^5�M��w`����A���&����q�-D����Pހ*jD~?DI+
8@������9�J9�!�|��|=�?,@�w���+j
h�ե�D�Q��X �KX���	;Ծ��<b@?���=�}{|'��H���f�I|��C�h�M��q�.��B���A��A/s���� ���1j����3 N���(&��]�Xq8#��}o�񝡤1&����4�[Z� O���OL��F���:M�k)C>朲q���� ���:Ջ~i%��!j�����6�,ޙ�ҷ]Z��#������b��M𧣎\�p�L�sg�4�lx��g���,m��J����7���Z�x��ыS�|�<B��t�K��ֵ�H����~i�'�ļ:���P_wN�e:� �HЈ�Ɵs�a��DZ�����$�)f@;��$l
�`c��8��� b
�j���X�����:�ŉ�6�C���Hc+���,�؆W����G�%�d��L��F����=�<�5.Ŏ�(�!H����lvܳ6�|�f�
�-k|��߳�:���P�Kk���$Ю?s����Q<UWjv�aR�ڈ#�y���k��"���O�/U��lX8��mz�@^�=��s�wmb�}�Qy�a^\m�#Qb���͎b�
#�.=g}�����^�\��|`K��Y�����RF��8st^��(�^�B����"���m���Wp��0Dw����%�1���F�ʼ|�����ul������UeI�A�G-�zU����ٱ/|�:}�"�6�%�������"/Gh�(����Rr�cH�뱩���r�фV*�R��Ì3��XW�g�%dYsd�"���ܒZW��ixu��VاAqpq��=���7T7/��R|kf�ˌ>���B~𑮎X
�K�5e�>�>��_G�gSZ>L�~�7Ke˲�Gn�=�%CN�h�d�|g��\����O��)�4e8C���݆+�[����~�԰���j�ǍS4��I³���xTW��Y��v����fT�6��9:L#�B��Bjge��ӑ�-���-gb��0�ԟ�Gs�h�_��:��S��*J��>��9D�*�c��SOw*�cO���M!�@�	
��*؊ܶ/i��K�(�� ݙR�������m���&���6k��C�i��^��G�O��v�~��'��F	H���/:� Z���׏�1�t�,�=Q��3č�����3����(��Mn�i�4��;]I��%{�Ӥ�G��q6Da}����t���J�oV�ͰA��v��q��O�?v�=��׮Uc�i�w��{!GUu!���i�M�Y��̦ �`��Az�0&RK�(�Γӣ�@<k�>����hl����gbt][�@�R�f-9�Y	IU�	㵜+��t����I,��Fy�#�̉.G����IR��5�&��	��M�j{"�r^���U�ds�iK��j��<���fk��$hp��L��ǠEeٸ�rJzm��>�_)/d \�����d�Y5��$B"]D�x��T��L�+�m�ν��i~;A��\d�7G�J�9Qܹv�!���X� � y�v
�md1Я4���V۹�ba|�,�"��g��^g�v�ڹ���T����w���0�iİ!�	����C>IB��^`���1ߏ�?�����n�pdc����X�����)!3�\����07�'�\�9p������#[��#��!�R��B.��NL�|f�5ǑəЖ?�/yM�)���4�u!~��OM��=�H4&kP|<��7ݚ� C.���Y@�F���n�I��������4Պ٣���H���|�S{��}3�C8�� ͯh���� `�n�8s%�xX-�$Ct�<������H��zp��6(��'�#D)Y�UY���%'�W�~{f]��բ
c��75 ��H�Qn�� ��s,�*��N�$ݕ�lr����7��6���`��g�6�ʑ��rJQ8�uU���#���Ɓq��kb5����	������3օ���dlaE����	b��B欿x�.�9[5� ��T�"�;k�%����!���O��A��$���v'�M����9�X�O�~rj&"�rqEA��$��ԇt�RG�+�Ux�%�e�0��ݎ�rO�yD>�N�S���
��D���mO�y��c�Xr��^~
���nm��>�]���q����s�Î��E��2䞼��7�n���z%;)�r3,�Ƅ5�+@��>��0�XH�����io\۪�$�C�g;���X��.��l6k�"��x��C�MҍVwHµ��?�nID�K�řn���
b�Ԓ�m���]H�H�0IJ����<�����e?�X�9(����b�ً�� ��R�0���=��*�nn��sp&J��"ҚӠ!޶� �(n�&�tr
aN7��zb�0��j���w	'�0~�����$5�Q�t0-y���$���y�Y����=�V����\��3T�6H��c�l���3���R4�/뤆�z�tp�mF.b�{^�ޜ��j�+�}���o\P�N"7�8՘�!g���~g΂���(�]�{��L���m�09����ij��ה+��$����I��]t �w�=D��C ʷ�1�+ƥ퍾C��T洢��wP�l�5�t6�zo�6Ws��|Ei'�>s�G�{�'E7*#7���H/�z+�W�.}���y��x_��J>x�AUe� *E����O (ֵ{>bV�dHf[�]w���$A���5��'e^1��պ��N�:~�5�+hz(�vҰdILb>R"��^�P�I��`yK	��%j��PLh2�ӡ�U���?��������٢e���Od@����J4BQ9D60��_��e��q}�y&(�#�kG�i�(�-2�S�B�6rXrb�	�P�����C�������t�Ɩ����C��f�+��<���dZ��rz/X��Hd8رDi��p�������.<������a�ua�Ӛ}5�D�@r��Q)����t��q�
 �;��ܿ�I���S��kp�����'r�;<ⶪ\�qS\�����[��T�ͻVer�����
�Y����G`:*~#��?`��B|v�B��ޘ���!��lY_��.>�op!�d�g�k����s�>���{�11ZӤ�%��$\k��I��Ԗ,u��0�*7���4A��w�fZ__F� 7FD�q�gy��ʓl}���O�>@��s��;-Q�(���4V�-+ �'��kF���Hco��v�x���sS�zu&��}��f�֊K��$�i�z��>�}�NE5�=��En_��6�C��'3Y����� ܋�zQ>�y&��Rb��YiF!�b��~h'ߍ���퀦��d��X�(ק?{����*�'q;h��������\N
6a�ẽ�t$�.��8k�.���È��IA���:�_f*4�~n�[*�	 �����D3�9ei��D���;����� �mmA���4���L���sSp7�ojk���zU��B-�gC��w#��m!V�*�TxA��|�Z�a�t�N6�v��[r���Yk�&u����w���U+Vy��Ns.� �7�9;�D��)�.ݹ����m�d٦wiD���q�"=0���`AOU�l����@��}?�?�,�x���My'	+i�h�n>#_�BP��	x_��^���W=@9���W�r�y��M�j��Q�L�E���!p������;�&w3`˷�)c��pibQC2B#�<2�T`p���>ٻCq��	���"/|U��8����S�R��5�d�Z�|`[��ѝ8��%�MW?�tZ��6�=��]�:k��~�O+���~��3�8�	�i��TKI�溽y8֝m?ܦ��5�$�2#�i�ق�>+Aj�p3P<�Bڜ"���ąH��W��I�z��6>,��Q����`�g����V9���{�l/�$��0��6��� ���7�4o�9�j��3�톍�|��#�\�6T�͑��!2�׮a[=پ&�V��мK,W����hE^�M]
��~�DXj�-o����R�>��Su)�z;���=0۪C�K�I��W����U�{p+���ܬ��H�I���ש��r��� �~��:�-��0�wa	���ٴb����qL~lm�M�b���.6qF�d�
�늛^�&".��p~�Ղ���Y�,�F��$g$�c���Pɻs�4cǐ�&&�H�V� J�z�~�0��}f	pEP�5q3�hnž�n�cу̫5�O�p�'��h�:�L�5h�	��M�(�m����0V��7��1_
���#��T��C[W�H�щt �:��Q,����q�X����&=��d�����]�l��g`7;L}H>>[�Tv�]{��b��{|n��[���jL���%�����0OL�����&!�K��:��cq�{���	�.��fEqq��d���.��5��t��3NdF�Ȁ;/����N��yf���S�������U�<,�tW-��q4�I�?�+�϶�<���]�C��� ��t����b��<�؟�
ݷ�j�%X_g�݋(,�����I	����/s�LwK��Ctr*�.��)��>�>9j���D������3A)3�hU�uj�Wr%pPR�5����qq�	��}��Ҭ���C��,������;H�`�G	��L�,��:�����L�+7��?�GU䇘���
3��I8��AH-�P���=���;���#�y۽�lv�5�E,��A�;ԉ�zVBiGX�I,������5���D!�����Lh�}8wϬ�*3��B�	5�C��3%.�����l�Ϻ�]�\�F�L�*�������u};����5
b��=�Ǫ7s���ߪ��N./="u9���t��!�&�{+�3��s�L�_"'����7M#�{	��y"���Q=�O���$S-�����U�_��XmH3��θ����+��>lN��n�['���+ԃ2�dj|���A51��a�7���a��6���j(�lƌ� o]?Z��Q�b�h~��E��+�#�QH��.��}�cA��A�y_TI�nb��A�C�{� ��e�`�q�U���x@4{#a��#�xAy�����		� YU��
K��J�B��%t�V����E2tF��Y������oC��-u�OY���7
&Q	�T�Ux�]��[�ӗJ�ѻ8LԾ� �U�Q"y$�ܺҭ]ȭd��l�-�o�/��1;�8�Zu���=�Q�ׯ|�щ8��[OK�ȇ���R����x1�0�Ӑ]Λe��VX�~s�:�y�*�R�+�b������^�ަ��z?s�T���8��ʜxs]��R��,cU�0{gO��T�K��d>�F�`�ʰ�^m{K"�^��jլ4�{{{]��Ph"�>CB�N�k� 5�0�:+	�.f>Ss<B��oTVq/�lp|<<΋��dI�\"��L���5	�9_�ݢۼ�
�ʠ�c=Qe*ޠ׶��Q3�5Gx�
o�q�Cm���Q?Pe�a��LO]�S�� �;�J�����u�|F�NJe˒K��մ��ϐ]+a��bd��9e��5�s�n�^({��@ӳA`�M��7�sp"x�e8�L���i��$>B��o�7gPW�S
믑���cku	 ���BA P��屃Ҏ3���?��~y*"#��O�糘^�Ô�"�n�(CXB�d�kFTjR��`<f# ��hw�І7v{D���;K�G��7��}��I��'o(X��)=�Ѯ;p	���T���@"h�������� k�%�f��0?��;���6F[�$�"g:n��t�� H�Y�а @����y��Ĕ�j��<�W��H�^�,���z\gِ�c��$�/M]��x���r2�I�l=���s�BX_��]�4�F#�`}l�.�����&���/��˥j|�Q��&��Gtxr��o��BѮ~�	��!1	x�5�A���ښ�ő6��W�����o���{�Qk/\?r���N�=ko��5����,)|�eH׼<�_���rE��f�c�TS�$uy�0�{��δ�9�����<�5'ҵ�~�6���� ������<���B��!����5�Û�`�
�ƭ���1|nK`T����nm�˧���(��
�Pz�7�l�j��&"��k�PƓ�Q=�_˻&	�P�H�]k4�'O�G�F��]�a�3-8:ܴ�+��'z�m�1L.�,�٬f��xn�d4�������%8�}���rL�-�K��N�c�
�tP��y�8��Fﲼ���u����t��`&DD�n��g�'�J��C�������B�Sw|������-#�]IsĄ�K��꫉���6��1~�\iW$�|�s����?y*
d7�����#���Ӊ��jM�a�����Š��c<�],r����zg��A/~8���D=`s��ȳ_D�J����ƨ�T��q��xC(�f�%�J���h�U��T�h��Onz��� ��q?�׿H�7�;V'��kP��B�$w��N�כ?�lJ��%��?��y������'V-�'���AH�p��m����p��`]��nQ׼�MU�?>����A��Q�,�G��q�+�R������kn*�N���k��]A��x
{%}C���%� 叇4�b�tN�h�W^���r�(MLƣ�6��(�Q���9�~yV��u�d��a�0�vS�G/��(I����_zrxM8�퀻��R��b�+�8��OF�Hд��{��V����\z^��m�.۹��_���m��!�q2u�*ǯ��7�դ���(~�C����z�e;9�/s	y(�#'�ܧ����ͪ=H��^x�g�����\�ɶ�8%3�	ѭ4eAk��I�X�%�m�)�&��܃�
R(1���tӁ	��@�B����)b�YLL�W�K'��Q�Gq��!IC'O?�~̯gP�k���ld�B�{$�#��r���pjp*\�Ѓ����Yjjr�+�����U��lJ���IvE�C��B^��1Fr������&�nK���g~��;�e3F�W��3�Z$�+',ᬔ��2s��G*}�f����l�lJ~���*	�!q�䬨zQB���TBdIQ�^�'ݏD.e�S�%��H�LV��G�������Y��˩��J�/2��N���T�*��J��e��D�����;47��F5�r��t��mr%X���T	��� *
̼��{Z�����֥.:�w`Q��MH�I��,)GDB�RU M$ӫaȿ�ٷkf=!��&�n$���}���6�[v��I�D�`p�GL���.�ޘ�L�UH%oq�����������{�>���Pz��<#�Q���eK�?"�I���sSL���t�bg��P'D��1��i輔B<l����D����R#�{Ho��6��>	�3�%�sWcS؆���t�3\V!�?#,z�~�3$?5.F��H�E�:�q�"�X�Z�eZ;$�H*�-eW9�9��I4���<m��Ͷ�pb�#0E��1$ۦ��b�IB��l����g"Wi�f[W/f�j���[�l'~H��a+��ZO�!2	��!�tB|g�7y�Gm��N��x��c�����lT B��+K�3Y�����!k�� �?{�R�:����oϋ�u��|i(K4)�
�8ġيwlR<K�Ze�-���R�M24��fYT�F8����Y)�iՊ]t��|���3g��g�=>��h>COf0F%Z!Q�a�/>M7�=Iɻ��i��eq�z�SR��h�`�װ���/Ù�����b���V@�Y,����U}l���遾/����z�i���m����pD��;��Z0�ozZ���_j_/i��@�AU	7�A���פ;�F�#p�`����6���'
�/��+��M�ܞ�k�e)`�D��^˼�C�@��K�gN�$�M�SSt)ފW�b�C�[�(����z*��G�ה�aKA�V���Y��?�پ(o9YcC��'i�#��oi���>x՛ZṬ8H�g�3ܶ�Ь�4~�ae��T`H�UA�nH�w��.���t)����V�:�<������@bd��܇LZ�[ `��t�:����ohr���I�Z&戰��E:�*R4�����|u$�z�=���t��hd�;ԨfiE*�^�gnA����h���nk�7k�����D���b���3`8����/:E�}0�Î�7��7�Ϩj��@$�A2U!���5�e���
�e�)�ch�rA3I�Ѷ�*��u���ZN`й9F*ptrEL
��jI�q����[��]KQ;y��/0��1lo2"�8`�zF���,�y��ػ �F�h�D����(�����.MRO�lt����<���	vs|Cw�S��c��NP�4x�I[3���#N⺻%7ގ桰m�~����Zy-����+sί�Y&�T
^_5��u����o(}�q�\{Ql8�>#�Zn���A� (I�h?CZ��H�H�p~�b6����q���k؉f��B�Ǟ��vYC��$���כR}�Ḥ��b�I�9��lɒ�Hl��ʱꌍ�܆j�kV����*^�����'�]�	Ί\7-$qh&�w���l�2DLq�F����x��Mt���Ti���+<���_u�q@�R��@��_�Iƽɛm̾��l�`��"QP�l��"g�_&�hQ9Ɉ��6ȏj�(�9�/��<��� ��V`�ZԞ0ƍ���N%Pq��뒾*�\�$B��p�@6�ש�����b9��Y6��K&������̅��x;�:w4h���o���ܫ�H�L�Sc��˻˸v��RQ-��$���R��b��b���?w.�(V @���X }��J���o�K~��d�֟Df>�PU���_��o#0Mr'��c��*Jx�w�n��'/E�	���1)�+[��\)��&��7��o���,sȬ8{�%p���ѱ�����%7��Տ� �Ip3�y!D �6���UZT,}���ʎlK��֛��!h_/��3���z�HX�q}�{,�9��N��Q�=�"��sR5_�_#B}���9��̻���r���#��]�$/��2��n6T���ɰ� �f�#�^Px0����e���R8hiC	 D:�0�rP��M��˛Dؿ�+�C��p��|�W�"��`!�Q��+a�,��A��z΢c�����{��̎PhD�B���&�߅1��W�񽲁��l�:8��$k�/�J�d�U��Eg�s�"���S����ˠ�7K�����˃o!>���g���a1���=\���&ݶ�do)����V��>�tN��Nܽ�?mj��O�Rg	�>��c^ϕ��T�`;[X��\��� �W�3�ah{��ml_��h�� zT6�5<������O�ڴ�2�hj�1�J�t`cE���Wf('����Ĩ�G�z��h�W�H��¾��\?���!J2���#Wq���\(c���TGl���o"lN�/P>�H�}C�,*�WX��'������� ��?�s�����e���$~;7��c ����[t8ZS�<�?4냎H�gC�I���}=��w���m���Hb�uX����V��O~�k�<v u��t'��L�#��<�FF�#˳}��6:�b��S	��`�]l>|yܝ��-f���~��"�9�J;��:u�33���,��n��~zQ|�F �F�7cz�]ǈ3��ut��W�s�@!jucdu�[�`8M'p��R�8�nT�-���Z�t�/LR���.݃�������k�C����T;
5`�H0�𰫡�VXA1����ϐܧ���1z���S��Ƈ#�z����N�qA�n����d�!�������fR�pxeIe��\6�t�A&�u{�N��h����7�.���n1Q�d��>�Q���~�=��(�tM����Z������@��Fq��&�֜����7#�����4�D���Q�HJ*
FS���I�ә(=�o�j��>�)X�%ы��n�G\�[g\�=�~ۥɀV6�M9_':[�U���~~(��mА�kG�4�$�jYXJ��س��k�lH�7H�O 0�k�il_�i�\��+"K{.���q�h��5�w0,���9�����L��O.��mӈ�����f�Υ%J��U�� �`�_�
�uwV�-L�,��n���G�O
�.I��f��|�3�AIr�,u"�+v�W�O[F�o^z�0���,��Q��Y���ًi�jGrA�����Q�E��+��x��R_�V�`r-)����}�ۄ�ZPNg�缦^��8��l�I����'�8��4�+*ζ���CDO��N��sĉr� F�H�硆(aJ��(Ӄ3��Ʊ-&[y�߹�z}+�b `�!�~T �D1�Ox��ۆ����L,]��n������7'��V��LDh�8T��k^�Iٍ�Ϝz=��c�x��{G�3[g��MK�2a��*<>]�E�o�9x�Cw�����jx+|L[�n�1��2�`U�v��mi�@��7.� ��ݳeH|T���-M]岠��VJ�9!)'�D��ׇPe�!L&gǱ�}z	pTD��n���u��!���>ft+�f�k2q
�����ϒ��?c&
��A�hѭṬX'�#ܵ��aE��@�-2��'5O-f���
��J��I�Gk"pUH?4��ί�!
��N�F6��7��Gb�U߃ٽ�i�01�����K����R��4�}��Koz��<�z.��?Z1lN�e��'a�Љ6.y߲���Z�����|~tz2t�I%]�v�ឫ_-8{��k���nN����*��n��4���J�8}:�fW���-��=շ�.
��>�/{�]
.�_'\q�d�Q��*	{7Cy�ɣ06��V�7���
�Ps��{6=����G���A�X��Ʒ�i7QƸ�%>ETaF�F=�
�Gȗ���	���ƕ!�}�&�C;Ԁ�%��.Fc�	g�"������1��h�!�d~�|L ��^v�Q7������r�.Ϥ��r�g+�0�TL���Ê�#�n
s>�=_Wj��"���yzM,L;�7��W�x�+$����<zlK..�����=�������*S�~V�!1D�5bB����˨���g�V�o��ʰ���MJ��;��_��Q�[g�qAܠ����U��t�Nm[A��,0s6O>$旭����5��2y7Q�l�x�	�ޞ���a�>f�G!��h���+B�h�&M��$%�f�z�Y�>(%i��mҽ���{J'��OD�
�=��0�<��|�QE��T'�87��c����14�*0��F�7�
q0�3��T>��촹�_@���HƱ_1�QlX�+�a��G�u�C�K-��u���8f��H4�*����ۉx�*�7�Ř'f1�y����:#KNo�P���IO@HmČrw ��r��1�n�eK�[�F5��3�(ē[Z'����F8�n��6��E�����Q�k�o,���O_y�3�AE-���ƞ��nS�H��`0���%g>� y[^Z��F�̥q�Y�ӻ�P�L�aAu� hD���.2����S!���8��r**KRo�\�|�c����4�-E�0p��u��Fl���:N:��=��P��7Ȥ����i�QFj����_�.i5-�QO��u8�Pb�y�6�+z�����3�=�l|&m��Yz��N�����m�2n�_j��)�%�ZMP��u��Ȝ� )ҟ~���@��	�d�`�`�=�qbÿ4����������Iʵ�D��gm�4��-��a�άdo����r7�ٛޅ{*I�
1�9�Q��e���D�o;��������r�O�vlCy�"��DK��@��6	�3&��m���ۚc�E�o��i:o4��M
�k?͂ݦ���_�u6���I�!�A��g*:�EA3�o��0ȱys��rR㗈���E
��2 ��(��O�L2�)�'7�c�3H���s����^N)��
��z�1�_���J�}���*��t�]�6�FYC�jA�����0�?�Յ_���pG��M��cA��lg��˦7���M��p�6]�t7�<�i�
̅�:�'w~nNx��]Le���� C� i�X�� _N���T_{c��Å!?|_��P�s�UoN�5�r���A�]��T��~�3޸CQga���W(�1���1a�dE=�}0kg� �҂J�fh�����㜛"X1�N16�֞hA�mQщg���M� 7�KU�,�p���tc0Z;/�hF�!���)���	��0Y.���Q�P!����F�H������%);|4�fIN�`t������G���R�=�e��!�.7v�ej�J��-q�R��r�Hӹ�u���;�p*�;�i���sD�K:!��]�����M���r%���IEw�1�N�����w䋸�8��Sh���DR)��#0��X�
2��H�ͦ�:T��r>)CN�)�9���{�Cw�݃�@���G��?�	�����|c����6�����\�ΓL!Qo�}ˢmI�b�u"%��\<�{�]xJ_��	=�
5E���K�|���:�6Ψo��{" )wZ�wH����fBE�6Z䯈p�O����K��O�L�����R��4��6rr����1ܯDMz:8�|���e�*ȧ�Y6�KH�-f?AHT�34B�^Vʧբ�_�F��r�&u�S,T,ۨ]�M�C;��N+�Y���"20-���j���J�&���p�=�*.��̍G�S*��^��3t�O6[IBt����ŗi ���-1��T���+2�#��h��z��v��[�;VYA���(A籋)�XKj?�m޽ZWH+����7IK�|".�฿B��n�o��S�/����y�,�7�ƀ���d.1���+>z![,aEYK=�|5E�7���{X;/�b �%nJ�Kb���0ϩ��>�T�"1��X����r��sc9G�ir�N����)��ߵ�I~��\u
q�	������[��*�,�@ls�ղ�ro¬|�M�>P���=m!�� �ڑr&�Y��P��U�E�""9u�{���Yȍ+#9~P�G�)e�շ��N��0c'�G��k��E�$7!v���X��>1�
'(d��uo�3;�2���Z��u�|��̗�^ي��o v�pL����n�4�u�y>u�5�R��'��	��P'�Y�����O�{Z��"⣂��s�!�fW�1F�ߖ���] (ӝ�{��X�ͅ��va�B��W1�"}O�6����2U�D�j*�H�K��[�xm&/Ӌ�܂��V�a�Bl�+9��Dz5�
.�0��7�F�����������?bX3l7��q�B��������6ZP�����xa���Rk�Q���tv�'ޤ�0�<��^[7*�� ;���DU����|y��y�9a�s�;D'�0t.�Ȕ)���E����G"v?�*H�
�E� �.:�5W!��L�Ֆ?���q����ݘ�l�q._����b>lӀ�t{Gk7��Q�O�&�RZ7�A9�b������]��k��C�1��F�Կ�Y�iI��Tn�7��=G�c��Q!'�A^J-ED�]�b0��>��10���Nd|���'y�(%]R��{A0��х7s	���A8\�'h�<fQKç8��MpCj���|{p�\`ֹ��Ӗ����SˋP<��?�L��L%�nt��h�!{f�J2�2^�^���D���!~7i��ap�G���^*�A���K"�Zp�px����<X>�qQ��%[K����G���?Es$]mD
�Q��E%���W�7���s��Gy�w'�
��::���ʫz��;�4�[�q,<@����+SFvt�G~j�u_j�鞄��dlm��s�����qU<C���`�2�o���.�H��^r��z�؈r�ľ0E�]k�+q5�M�B�î�M��߳�TjՒg���#�eE�9���Xt�3�����V��|�a/����0��yūn�-�gM��ʤ���e0�<A��V���ƞm.���0"�q�^�L��}��$\0F3�� ��:�7�T�2e�0�S�[B��Bn<��K߾�#�i� � ������D/�h�S�?�MFA@Ƭ�������ڱlOP��pa�
���7�<Wܺ�F��[�)w���%Ha�������W��n�xbr;� t��5A
��xB0�k�Ӿ�u��w����	4�J.j*�x�A�#�7sD�a�l��U����3(%�'Q����>5���v�c���b�}>�'�E��TSL������T�2Wi���28������j̏FR|r4)���0/��`�̴��A�1�0:�I.���tq>7k
E7�Z�`��tx�rɦ.���b]�֘9���rC@5�̾OE�G7˟BR�V�x�m��h0�Y��Oj���p��>|"yb���֨�?��*G�BL<f:��Z5ՌLb������:��&�`=���D*OY
?��U����{O�b=i���Z�!�[H7����'���%��	���&�!�y����6��J����^��c��5�"�]d�봐�^�ꆺ����:�.��Y~�̙3�Sk��W��%b�b�J0�s3w/Om��5J�尌*F��������p��y-]����sne��9	G\&��H�B������{	���l�nk�V�I�͏�X�d�-��#Fs?w��b�2TP��M��>T�Pp) �a̷"$�l�=z�4���ߘ��w	��g%D���0�-�<3��o�oje] �uBk���^J���S�Y���_1�q�\ac���障7��|J���FI��q�!2§�zYV����N�V��_����'.Z���>6���zȟ`i
h��n�4cj�
�q��������ԵM�6ǧ���|�{&&�y� �8��������Gt��x��<Jݽ-V��7���I|B�dע^�[�I� �l'a��K� r���ER���M���7������6��։M��YN��\�rJ@�Kڥ�b|�$B���EĪ4���Sz�f��}r�{L|.��ֹ�?�H� �.�+�� �ڡQ�H���	v]�ھ�evD��h*�
'���������� �f$[���_c/;��������I�8O w}�����B�+G�{ d���?mJ���奺��%)oܳ"��=��O!gx�&�t�v�.l���ƫ�sVh�ò%:�#y���zx��b?�ʖ;KeX�x"Y�\��k��l��ޡ���0j۸78jR���3o�@�a��2������P�,,�)�Ț�9$F�͒j�~δT��A�Q�֒Ֆ�|�8���u�vh����OV��BFؗ�t����/��.Y%�i��Q�L~M�%.H4�n�������y�rqюFi��:�C0DV��F�b�!�_I�o�`��A�����>, p�'j!W�.uƼ�u��2�0�us�j��(N��������@�-�~��~�f���Ӛ��&V�/W3�i`|B��(Tv�c�u)�[	�#^Ed�b��\z�C1Ԣ%`��n������}����_�]$n��<i:�@�ԏ	�A�E���G�0�a�����}D7Y!�ݍx�!�C��pF�@��:�C�
�7"�gtR�r�}r(��(���L�d�R0~wf�7���n�6�N�s���0��	oF!��?�f/�ܑ�/�L���|:������Jݥ+^���U��T�V4�t�u�Hf��!m�_n*ek�����
p.O`�ʆXg��E�\v��6�;��O�P�O�@���yj�N{�w���,��4���)X�ΰR���_�Pd�D}�&5|��DSI���"�=L�/���\�~��B]�:���3���a}���p�����yc#�����ۤIzޝ���g��}�sH�� }��idl�(�F-sLh�� B��w�h�vd��T/d3��(��P���"S� ���P��ӋD�E�m���$=@��|+�á����~g���{&�Q��L��Ny��2U<��A"�N�F��E?a}O�hU2?�����=Fu46��-��˿�h�~���[3��ʰ�JA��,I.[ug]!�֢~i�^�i�τ=�،7��n�f���[�Y(��
z�ܵc1u�5���/���	���>¹T�;5���%��2�G��������{QXZ2�Qʔ ��<A����fR��z�~���#�&��f�xF|�蔍f��7
I��鳿e�Ȝ����3�,�5q�7���� �˓4.�O���LF��a�5��B�(��G�׆s}���1�$�%Lzdc��&"�	��nԓw,*�o+xM9g�N��`U8�e�u9��G����a1������ݬ(�Mm�Xz�~w	���.����H�~�OV�K�h�3�.c��EG��&k��Qz4�0�*������*��"F>/�$x;..W�`fj�i}���K 8���e6��N��2z��+j{�����I�>�Bc��K>�q�������*n~�
5zb��i��m�=�FAiɍ�ZiW�a!���AC�����:#T4�*��;��$0���m��S�Ǿ�|��"��q_��P��c;s�1x^��Ϡ�x��6@L`_��#q����$||M*�Ƙ	nq�s�bh;g.����Sڱ�\���V�)!K�O�0X�֚���Dn�Ě���Bo��ӛ�P���Q&z�j���3p��%�pH��؈����;V[q�jexe�H?��ͥ+��`rꐄyѢ�7ƽ���"�Np�b�}bm"���8Np���Bu������r�fRIG��ua���JfX&>-m!H^����7����4�/9�p���bt,�`8bn[J���{?�c�<��[<��ꗜ��z�p_�h4H��w0GkK&����x=�C������(`D�r	���xC0��Z\pG��cx+'=S!�9B�oB$�"�SK�9�&\Z(�cE����:���ӡ~@��h��@�]e�A	�\ҳ����e�5����5Pk}��yT�o�$�~4���KL��$ �m��RV�+
R�6���y���l��Gs�����.$n4��#OG�0y���Gudُ����TA��1�����*��n����KO�[4<V��kr�R�"r٬D=qDm�h�б\/#�f�����ˎ��b8�?����7�G��"���,�vR�tW��;���#��+=.��C�ֽ*���ʅc����,��@�d��I�K;�\s��W���[�Z��\D r�.��(^��z���v:�Y��"�T��AƊL�(�r�9��`����\|�{P)�v����ݽ*�b����.w�o��؜��oA4*����_G�u8�B��]_ª1���̩,�~�zd�J�@�])�m�`?	����>�S1/�4���b�g�E/ӟH� ,� [ޢ,�����sL!�����+"�fZ�<ʕ�^��(|�r��q����3�tY]�]h�ӻ+H:���6��N�-�"�����^(Z*���O6g�)?v�4]ZHW毾����w/'�\���#O&N�Xp�ѵ�I��d�/�tS��<P���h�Ͽ҉T�#l���	x)+�7��H��MN�p���Y�uE���O:,���>f��c@��b��P޼�����C�(W���¡���M�8�=�~�aJ %�P��x�$�n�o'�p@���3=n�Ef� +����=3Y!݌^p_�7���m���ݍ�x�v�7��є�vV.r_j��uo���H�q�6�.A���fm[��Q��"�7-0}�d�|.��3�+�J�yWmn�z�f�EI����]'���@����M��XӬ�1��Ŷ��9L8����Qb���G�N�-1n�FΑ���ߋ�?	?|:"�� 3'�|�S�<K��F�K=�V�0d,�g�m��NN�ҁF�C�K߶��{�ױT��" ��v��w��tT�T���!���;ei��į Z�!Ql��T�Q���Ow��=�C��:��r�f�)��M��b?p4�@:��u%�n��>`k��Ae�JC�&�����;���Y\sQIFa�A��u����ͳ��4�A��[-�@,)�#s	.4ɗ��v}-�����4�}�B�S��*х�O��~e���͛z^Җ��7��5���Te�r�L�dl�,��N�Q�P��c�.Η��k4��e�g��^�/?��P����w�!���aZ��?�a�:V�d��|(>)����������K��P�w�V�*��!6��0���c��QA�]׋�w.?�+�^�����1��9������<(��Ӳ(���G�����~��lb�*��+�8��fw�)�:�U�(�F�p�C��WE�P����`a���xBu�LE�ea�ˣ����0�AC� N�P�	}��%A �è_X�^E=�to�k�r�F)E���9I��S�M�>:�C�vV����^�[	�ۭ��$r&��4uʹtb�g���_��D��}�:������$]2Q=^1�w����#�����l�?G	�8,"�g2h��]����G�f��YvcR��U�qW�F1�$m��~�SwZ�H8ǂn@����i׋�EN�z$4(VE�e�&[K�Ŋt�@߃��-�7*Ln/�m�1+�7{
Q�,O��?=F��Ŗ���A����@3� J���r�\s� SK�T�J�)7!L���#o)1�6����j%"\��,����h.�!��P��䌇n�P�1O�i[7=MC�_��{�4��w����*\6K�~j��b����ׅcR���#O���k�ӥ�)_�Y�^��������Ld��.>S��e���r��*:��[��w��`���P])�e��2�Ա���ro�/���=eM�99����b5����Hq�F������yc��C�m�TQ�]�`r��p}��)���p�c��6݉���V�{p��ox���4�d���k?
�%1����i[ES"b��i�%i�E38�]B����^Qԉ��.;�j��@�	[ƭ��رR�AE�	��\�{ql���m1�'�肊|=8�{��R���̟�@�%W�o��3Y�#n�s�b~H�U�Õ��G���M nM�H{�vj�����/N��x.ٓ6�+�(�n���(b;��Z$e���F֨������� 6@X�ۈ�Xrf��pA�Y-MIz�)ZJ�Ţ����b �����n���D�<�B�����C�ߺ��y��äy��m"oT��'o��H��`������
\%������d���ѫr/P*�������FӐ q|KRsH�Y����GP��|�U��dW�&&�G`���NxH[C���a?�њ(?vX��H%�˽��;�cШ�A��}��ߋG�	d�_��Nz<�\�˦�x_Q���m=���e&g޽�T�Q�O���|}�2�dǘ��C|v`�o�9k��+M���"���h��B#�-,�����%��!&zq�$.�Rg��3ã
	jk��t�S�ý�q��6�m|�s��e����Mk�F��|�y5���FcX��i��k}�SO�Wbc5��m#9f��3�FJ"�
��:��ۓ�c߾g%wV�y���F�T�I�"��<=JE�q���0 �5ֲ�0Q�a�#!l"�D��H�>Z�UT�֭
����UcԐ��r�Ls�4�JP�-�^&>f��#�J	v����;%n���Z���L4ǼgE��h��� �戽�L��fj9�Rf#��Z�UQV5߰v�٧b����[��§	6O�z�ڳ�x�Y�Ǫ�7�7��T+R�]O}���4u�TƴU����BMvN�d�����%���������Pf�"��"+D�wY�9��u��*��?�~���J�L-������@K8��d'�?�I�korِ$��"kafqK��ĂA�={b���tȕ�4w�O�%�t��hhe@�D#�əg�[�����Ȁl4���l{Q�����V��x8�kM�0˾�����H���0��P���a���l��?�{F���-����X�N��h�a��K}(}�A^ �:"	��a4��1-ipl�}��rƝHhֹ?$�o?���&y���6�yp�v�,��l[%�6P���'��f5��e���0����p���ZG��O�1��7����I�����@G�� %
]R4Xl�Hf`B!��D�k \X�c ߢ�����k�ǫpq���` ��!��(�	�F5%nQ׫�4�\V�̯J+�����#u���rb��"o��,>��DW��ڥ��\%�}�=�(=�1b7X@Z���P2!=��kN<�yB0ҥI�e$s�,�X�J�c,�L�����7�2]���w�O��1Q��ʲ�N2��%k��T ��VI3yL~�~;�ݼcA6��)��{�I�Z�%��oO]���y�y�{6�: �-���:N��]�?pj9�0���fZ���=��F��N�b[v�"����z#A���e� S�٭i�]r���͑�N,/�[[��ph��q~�_����?�L�D��������aK�҂yp�>Z�	^N9���g(�y9�Xa:�d`��T��y�O�[a$����lH�%�Y	+�Y?d�;��(Z��V�qXhi鞬W����;�>��9
�����2-�I��ߪ|V��(2*1U�������`��Mk�@���*�rRX҉����U_|\$�ajkq��V��:1�WоF$�z����2U�C|W�N��U��L��U8��"Ct�6$p ��K���a(�������z�~m���JХ%7��� hU�~�WN\����6��0����nY�2&���@ ���5��8���6������)O,����M���bSq@���#漎ȱX<���l^��B5�%��/z�nIC]_.1I����unY�
����E�W�D���?D0ko��Ӝ� �q�r���1����''
N^{k�4�"�0S��:������Y��!��۞�!u{m:�����2f+��e����p�{��,���P�_�ջ`X�(c����� m2�e�m�L�y�77�M�֣�0+w�]�o�pD��}����.��0|�P�+�Ig�@ƜsF����({j��/��qb;�)��wh��*i$#ƨ���E �]N�䏦�^�ڮ
�ݑ�*,ַ��{[)w��$?j4<{�lĈ'�R)�h\"�+���!��oGd�$�8C�2�7OX9�-w!�O<�iW>�R����DUs�񨽝�VP2n��K��X��s���&~C_��f!d���#���-La(�����%�I�)JE�Sl|#�"��b��.���	��V�~t'6��EJ��v�>�W\����ʶ���٩}O�ո�(cf�'o�&�)�/��_�j+��b��W=(��F��U[�|b��gLƞ�"4��8�J�<LĆ�&�ii�K��P.Ђsjw���'e�;�'�r����P| *Ek��}�^Pt�rAvH�=��r��]���Ձ��i|+	��g=9���@��au|�Vz(8���r%��ᄓ�9�:��,���.�A���A�������[���ť��O�+��1�"X�����*^+�Lw�0w����	��vtXp���݂�>��<nsy�{Ԣ`^���*�'�z�& ;"&�<�� �)�B�+��w�?�n�V$���G1,��H��ܨl�1�Hu��Ljץ��ݞ%��k��k�g�:��}�
4�M�8 T�	@��#U�޻۰��7�4l�ऱa1��PeWm��l1p�JƎ��L�@*O`����~U�B�ΔzԷ}&��@dH	�@k'P��x��+�9ֆX�.x��dk�������AGQ?�����ښ�Ѻ����G	bfD k2.�8�!Ϧ�k7��{?���xDT�>�3��x�i'�m6��v��/$I�&�u��,��V�$#���k/L��{�V� ��4�h����kJr����(�8�-k
 +;��t-65Flk��s��<��S�efA�+�x��4޳��)�@S�O�����a7wC95R�tE� t�U/��8un��u�Mb�� �b:K�
"/E4���i�9�$x��x��Yzx�/�n˽u=��c@t\��21:v����b�,$�t��_cNb���y9�Ot�#�oa$�:4�`T��Lp����	��jX� /��r?��6[$X�=�5��!T�?>1��^Wܦi�/�jᇍ�z���+#Q����&�~����BBA���2�h�����m��G+�"YU��Auf����I��;0
N�ea�D�).��:��=L���5�Z-�1����3���+��l���J@U�����ڤ�1"j��P��{�ɝʶ��>�+�#BP�s�ٔ� >�f�7m���3�XB'�.׺��T��ˬ�=6e<�b���`s6��jWZ�ޟ�u��D35�i�'b`��c���0��<x*J�e�p�����0�P.TY0���FN fcϤv~�(��PӘ�<��8f\$_�:oC��N���ا��#�kb/�ƛ�bB�P൉�)�Y_�	�H*�u�N���$�,e�G�{/���/;hO�_pj�#�a�����"�'f\ԃ��R�fD���-��P�%*��-[Vm�|��d���,�k��=$T�yjT@Awif�P�śP)E�u�WӤ�$����`�e@:8j�lY��Bn%��t jl���6�k~@���%6���,U�s38Y�h?�Kr���U���p�i2y�������D��d�Q��O�g������[N�qG�1��%�e�KES�rg*o�۫���|���g ����H��h{��hݽ��������)�����
m��jÓ	 {�`\��Y
�����?y/����S[;�����`�?.�w�ڂ�)���L���hQZ}��5Bq!?��G��Wm�+�@�7���T�}�vڲ�k׈_:� Sq�.��E��!��]�.���>��m�# �O��rd�nF�a(���5y�Y��6���t#��K޴��g0�ե�R������2���;�e�
�bY��qR�,X��L~_�J�r�&�i�d"L��!?&$O�3�A �Y���	'��$���4���:�#k���K�W�z�C�5ɦ8@��MDYj}��0�RC�i��j_ǲr�a?O�*�j�K�rw���'��R��'�떺��T��"�u.��6�
\�?�O���Ne���X��l����7>��G���댖�4�D=����Q(�����&��]�fE��A�@�C>l*j�f�mjZ��t��<�n�æ��E;�uۧ���`��B=��i�ȿs�;"�7{}9������x��Byvz�ת���tӕ����h�İ�
B��}.��ܝ��Q��5Ɯ�XP���C.��|N��d��>X��0��(��J��B���';O���E�%8xhҺj4���쁽e�8��Q��w�JWNj��pwvv�2m���ނ�[��m4}cO������H�iF��.�?1X{�}�N��XD	ϗKl4���G�p��Xc����9P-\�u�Q�a [��Ws��Tx��霂H^�y���]�4��\��:���u�)^�=�z�q�s���{��x�:����+`C�j?`b�d�%T�6=�E���l�� *#���u�Z�̡�['���?P>�M���jy���o������ց
5��?c����Lm�������\��޸�t�����?�>��%06�m�Mv�婙��C8G*7h��<�lu��W1 ^%�\�,C-٣[ACK��(��Q�$._l��
����lc��o�R���擯]w���!V2jta��%��n��z�.	Pp��*��ɟ�M*K���!��W�]b��I ��:=�7-�e�"��H�#t��ϖ|nA��S���{�G!�� �|K�(6����*<o^h����\��x3�1��^���Ml�;�����Q<���'c59!��L��zp����/�<dr#F�`�'2�/�Fj��,c�%��s��Y��
v0C�`5�e��{��-~e]~�Ո��.�}�MO�v�9^��:��}�ڙ2iU��j'nG'���׿zd�F��a�% C�K
z����S,A,��g�{cFm�&���)s���ZNN ¡��=�L��C��5l�p<bޛ�)I3{﷧��E��qY�����"�L��x�ڂp�H�Z��t��?��c*�`��hJ�� rک��%M�U_Z?���p�b���20
-8��?戇��q:o��f�HKx�5��V������9�r�y��vG�& ���گ�]dN�@�}�B�
��)�s�,�2��g�XF��$(������?\��zE�"��e�%�Z��2*A=j�pL�tP�?D�qL��O��zpu�Z�վ��lr��ܬK2i��O��Π��g5s�6D�lyK��9���q_�)�50��Cypr��!�D���N��TLB+
 ��-Kn{����8"��ŉ2T��`�:=翑1`wjг�7Ki�-��E$���3#� J�.4ї����1 ��oP����6'���Gt� |r�U6\�x��Θ���f쎋F�O���p>F��Mql��K<�6�튕�N)�ׄ2Z#b���t'm*�~��qn�
���9���1��iL�AAo_�O�Ka�J�(�H}�~�Z�� 6�5��\�w�����M�N�ɎbR�����v�ǝU�>	�V���ny�s�vYA8R��^԰���@h|I��G���	��A���D¬�XC}����km�v��<��mK�W!�&�!��d[(�ys�:㱹���f��=��f\�6��dX��� �ӋQ�Ȕ�H-N����aN�r�tH x%EH�ˈ�L��h[��:[!��a�j:��˸D��&���s����eU���gs'kk7/��6���N��r�E����e��s����"�5W�P<��Z��Hū�O����㯻d�����	��f;���%��YD�J�$�*..Y�/s�*��3�;S#Ur�XW�bI?�Vi�/ �ɞe�w���\U�3D?dO��Ax�c�	���e2����m�ȑS CeD���f�h��U}�;^�Њ�Ġe�='��賓|,�d�h�-�|J�)RZ����n�j�<W�1��u���<�l�è�3m)-�L=��8�,��~`�"�bě�� aH�a���Q�j#��a%��;�6��#�rg��)[Y�A[dI ��N'6f�9��! 5�3z>U�IJ+��~~$!�XK}U���?���k<���8����&K|��,S�!��=�۟�k��{b���<rDI�J��b�e�GM.B~���>����g3K�
N��yN����/Ct���w͊(���kK_/�*e? {Y�7�?23���S�X��70��biR����9�Io�{[oq|���cZ�8a���M7�r��׳ -%�S�x�
2q���l�;����V ��]�$��1�Sdp��c����5��{�>V��c�����7�_,uC�s<��%�M��(��>��wA����wSJ�c��y�_ȋc_m��ܛ���,Qz��$��SHSpj%��C��+��!���o#7�rj���<B�;�A�`K�MW��c3�̯���,��?��,dח�!����GZF-R��M������1{�??�ki0�ԄZ;���C���ٻ��g�[Yiq��i%��S�S��هMf �kW��`1o�:0�D�F�KL����G�ZF4����E�8z$4�k�c���B�b�.h�R���9�ՙ+5[�-��O"�v�8La�����]���@�~PN�%=��Tz��%Q"UY1�y[�eL]5���Å,n�v4"s��f8��+�+X�@�E�!�=��_Y�9.�؍~be�w����[yk���(�d�N����"��i2�M6�{��L�q����X�����h��̻�
�w{\0�r�j\��[���?�_EnO�*�%�0�Wc��h�����f+=�Q�;P�l{�4Q.����oa��@�[�&�!�}q̥e�B�UN�sy��[�:��b�Ʃm�t{�\st>�	9��c�(͝�]j��n��V����8l}x����5����iSm���le���?��@ �TP�OT�-�<��ht��Ҿ%[lC%�g5)5�En���*�8���K���f�}C��p�q�ve�����Ʌ���7��C���3(h%az�OLY�.�1�M���΢��};
����C]�\����.��U�i�i����8��}3{zE��a�3�`���w��/�h��dAR�~����q@x:��W{s��5,�q��n��C��򦕲� ]l��qC+����J�:C��g�NOo�' �-dH̋kB鮈ݰ)a�ȱ��Z@(�O�4z��f����u5�3�+�E�vp?ǥ��<�4�j��RQ� �|�U7��?�05�,�iz׮2�g�>9���ܝp`��M�S���|�IA�?2`���˵g��Hx�j;x������bE/��F��"f�]�ah���������)�@��u��=�zk�_I�mǲ���:v��]�a�X׷����G���]-.�P��9���R�G��"C�3G�x!�
Qfˋ�p8BZv�l(�E,6a�6��	P�S)-�dQ�*.�{�d��n.�xW�r��uh����o%bH�o��bY�R�{��B�p�!Õ�8����$����ċ*�ѝ�q�uɄ�Q!i��]Ç����P��	E��#>�`hOb^b�#aB��Ic�XgZ�[��}��L*R�F�N2��Z���e��1'�S_)o��
g�=0���sOQg�ݫY�T�KDZ�Fݝ�t� �\�asT(�y���kJ�m���=łP����6*���V���n�_|����t