��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�i��a
Α1S%� �uj?�L�3��TLei-3^5]E�$����/ԄDa��H4�Q\��s��ʏ\Q����B���x�r\�a�ܜ��L>E4&���L�F�AxR����h�m���W"`���^� �Y�~������B�k{G�=(H&�eM�5z�*|B'iwo��y��&��w����b�B}Ϟ��q���5B�}��ؒ�<ϗ�;��ap��9]�D����ZL=���_'P�R�>4�\eZ%��}
YX٤�ݘ�ᛕ�B�b�����b�8X)���^�}�^ϴ�������_%��/-�{��ɗ�QX�0'�����Ƀ�����"Z��;z],B�=�R�Iirl.���>�6��Bk��0O	�so��r4D�'W���PB�^w#3����j�����~g�X�?M�
ޤ<}�WZn����<�:��cE9�<�7.<X��-���(U�}�\���\�@��5z�Ǆ��:�v�	��4�Dpt?O���*��}0�����p7f�<i|B�r.s�0��"<����$(��o'��(%�]�ջ�nrX<�tz��U{)�f�a�%5ౢ�7y�δ�5���vvA֔�� 
V����R���5,��������+��.�l�2h�~�&Ͱ���s��X���E	��|G��c���Т�q=���.y�ׄ���x/KMn�R|�o�Eo�7��\*t��L#����ºL(�V�ފ�o��_r{�ɂ �=�ʚ�-�^���}!&�������$,L�K#Y����|*B����=��gv�aŤ� U�n��Ȩ_ˏ��Y�ۿ���.]5Wd���6-�X�t�[����I���5�]�.^G�i�D?%���V��^�ZES���=?�A���J`�Mo����9�d6���5_��ya�c�{��"����1,
���bҁ%��X�sVϸ lH�D�o.�m�B�ˢ��r�?�O��"�R��5�7 v����w��fz��!>�w�Oo�Ѝ�[�� ��QǧE�w�q�~�̆(��- ����-�]�E���9ԧ<�2�� �T��J���{(�!*wdV�cdrrP�a����Y���jt6��\&+$���SPN(&"k�@x�'sY�P�j����LD! Oę�y:r�<��m��E'���%�]Bxz���'{�6�F3`0�$;�*$���T:��0�
 ՜�o�Q&뷵!�L(�������b���H:��I�z��G���P-.��/1�a�v�]��l�آ���=�}$��ɠc+)����!y�׬�&;��tMPY� P�6L)T	�L��X[絅��� RC�蓶2��Ƿ}��w9���q~�$t���Ӛ����Y��Gw�>�-.�?��(#�.ށ��`��1�@���ci�cJ����j��8���44:-��r�gcJd��g��-��:�2���R����A���W��d��m�j� ��Lq��mɪɐR��w���g}���U�O+>�a���@�
���_�������*Ѿ+�����%�^���{:Oc-��2N��`�fKl�+���˂3�b���#eu���ׅz��$��3�&"N��5<nu���j`2�lP�q�ݯ�<I��"�����X����W�;,�K?.��,��P��a\+	[�_��J��k�
�vCw'l<��!逭7Y�hq>�d�Q� �p�}ĳQV�
v.6��h3;�A����`�K�!G���h'�k��骣�7_m����҇�Y�����%Pě�tDk����z�/�3���r��oM��gi�N�����?�F(���/�ա#	��.H������m�Z���T�^�G�ftz�M�j%�W+c;���ݝ5|����Ś���9���A�����֭�B�����i#,m1���sR���g�_6$��]?�j�l_o�_cG��̥8㵴�e��zMxQ0X�;��__� G��򄂵�E�����^�NJ��ٮi��]��o�Y��o�m����><�����3*gg%Z1҅��������Rt:�t�!��x�RU�Ѣwŵ�@�E��⶝��p!Y`շ���r��"1�_4S0$D�B<��?�z���t)Y���c`�7�CB���ET$B��3>��������D����b�ォ~i��+)�pg��6��͊6{r��O@Osh�� !/S���n�_�,���#
[�0+Ԯ�����8��-��1�=F�@T%�^<�WƵ y��Oh�
&d��i��&4�i9��T��fc��w��ڶYզ��{��>/R=��ޥ�iėF�#�X>�cocPW�s���a�S̟B�K��^񙠿�m�@rp�^�E�5{f5'��Kwg�4�t����#�B���^����R�?h�+����A�R���� ������5�С;�4����aY�6��d��#K|�|* =-��&�h���2���b�W©~(��lOG~��v�Ox�Ӥ�9�0���8S��1���Y��)+'�BB��1�>�"ȧo[�d�Ŧ�E�H|,3��^�Ҋ#�ج�����"<v����=b�� +���yJԿ!3�tr�tR���ݢ�i�]����'m�c����:����\��$�. ;	xw�qu>��|���m��̈́�0:?�!��*��t��������6���S\�T�����]`�b����^�9�H.f
������sh"�W��	���6K,ݑkhCp|Y�f�A����[�J&���в��ɪb�N�و�S7�x��:m��CVoUQ�m��o��iz��ؒA5
CǶ�)D,�3R?�!�zt5�-A�����	PcST��i�����ڗmp*^L�!Z�K��kE��$���a#�GW�VBLփ���]qT��ƉYK�S�����<e|j�gok�E"�Mz��TVӧ��(����[�/�GO�%���{��{�	����.��$R@��>oVe<a�)/'�6@�o��q��\@%R#�����K���:�M��@2\��_���ݡ:��+�ۃS�S�T)/��{{K��
�6u�:9nQ�*�K�K���̋1���Ti`��~�#�>�����t]�O%;Eu`�FGZ��(�E�	���ڼ����
�}ƺ W�8(��1}`��ev�����z�hN�����Ww8�3O�t/��M�]=�:1�<�K wf��Hܘ� ���R��H���xfq�����x_����&�7A7Gt��W�5	u�����˕+���)��x:�A�N"��0P�hZ�� s.0Fa�YK��.&Z�o�HμhpU��lQ�$L�L��#�C�W�f� ��`��}�����Nk���� �l$���1�^*�X��_���߅�9�3���%���A�y�����+N�k��6��w�Z9`;���Y�x�FQ�e,�dXۂU~���ա���/��D�Ơe1�a�J��v{3�Ć4`b�Xw$���9������[��Ṛg�3f�v�w5��)ti�iJ����o,�`��#��bQx`�~��W��u�%�j�Y��Pm����L��j��[�Fl:�}�o��
=�6�^��U*ܷ��=����*�Agraq�P���яy���
\�&��J�v>H��\X��qi��W�]:��� Pl�Î4�IE���H��,��Y�ϴ�37Ù���<��DP]��8�N.5�,��4f郖d��*U���$sw��٩��I��л��oi���>�]ݔ��!h!Z�mX5z��l��^1�83�pY�J�rg*�q�����\�2Q��*���������[C�t
b�ҏ9�=�wU��2	�R��!�Ҽp<Gh�^��r�L�~�ߛ�2������.7�o{�{mN��S9��V����&�5gz�l@��"��D8��i���t]�F��}��c�1�^�9X������\��̈́khwS�+�6O�s��P p��f�V�=�D��]�6��g��I��6����s�^@�JQo\R�ݠ��� 6�_`���)�?n<!E6B�$PL�ʨ���L�{�w�R��$S� �+bT���>t�>~��%�qx��4GiU�HԸ���ܩŵr~������X0��G�^�lC��CBQ�Dx�D�u$n�d8ج�q;6A�`���s��C}�ܖ�c[_�m{��@L���X�^C�%��<S%��ׁ�)^7���M�S�*�]?�Z7���&���gx�Mj�n�C&[O�0���h���E���(����B�0�����vL#��sA}��!V�J�w(XQnR��� ���W���7sO��1�̟�,��w���6���ՄE���d�U��$
c��eLA���@t{�
S� ��-l��E�͟e
|V��'0��B��oO�%�BEсA�u8�-N���,(#+�{q`�t� ��i���bرY(��2����7p>.C�]��/�u���9}�ٳ�L���b�n�gI~��J?��L����Aܬ]��N���YJ�ҡH^��Ah������T	���?8S�U��)�
��)t�Z��rAt"A{�C����0	�(�)И�
�4��x������O����t�ovA6����>˰�G_��I��(Bom�����^m4��l�Zޕ�89��-I��Y���q����D.��,�����)O��l|���|P7~�x���ͪ�~7苀D�$<<�%/L4��:q��CdC�8����~Aޚ�w�iFG�V�J���G�7i,},�f���}%��D�k0��w�����)5}�7��������c�o&q�a���3l���݄��x�p�'=}�i3R��B �%�ׯ�x��3k������qe�4M4輼و1cT��<�	
u��A��^c�߳ɩ�V��Y��=ճ�r�s����q�jf�]��"�Ek:�6d���W�,�Ǿ�1�9�[F��(���t��fi�v��,"�O�zW,d?Q	Re�;u�n�J�cg:e*ِ�j]8�bK�[�^<�}ـ��5R��2�`��G��RE��-b'�K|9-�*�}���Z�ls��N��ځM�c	kЏ�����h��H(�Z����+�X	nX���s�9�Et$w�7`�z�V���>S��瑎c]���!�8���f��4G���n) �8oP���*��dl�`e��P�S��Ίjr�/&��iɂu�N�d+D<�ٜ�����s������
ͮ�G��"j��wF�X+J���2�:���xW���twd�a�d@�6� r)%̵+ A�ipIQߴ�6��x��8�B�ѭ}�\S�]1#�K^�A�Ý�=�+�nv�a7`KRVB���QOwpt����U胳���b,�Ɍ�e�؏��=�b9�|��@���L�`?B�G��j��꺙�0��`$��k�@���9��_���X�E5S�'ױ�U��lvQ3�꥘چlt�kz���M��\i��,ߏclX�L�8"�E��{ɣK�1�H#Lo��� -�.�u�N�r�~?��K�Swf�`����ʟ}���or��9�;ֳ�����gJ������q���˱ �T����b�;���87�RPw^��:*{��i�� kל{:�0O��D �eXޥ�����R�s��X���5(��G��XWF�'��Ȳ��#�B�n�]��r�e����!ߜ�[{%Uh�S|P�Z�M������%�a���8M��54eJJ[cؠ��<��z8����QS��N�+ �Dkۉ�
S���]�i}�!EI���+�Ql=N�U��=-/l�k�>]:آy\dSO��
�bx����[�e/(YbQ+�#�"A��a*aM�ú���r�5�ˊo����% o�t@=���嶯��q][��6�$�1����o��x$�L�z*�����j�Z����� �6\�j�t�<D9�$ȅ�s��ht#��ɦj0� r���S���òK��R��n��z$�<�B�(O���qz4���RI����{b�$<s���]V`�'mu`��VE���AY�eh;r��0.Ŏn�i�Ķ,{���he= ����ː4���6���}X��䋓�ؓ�}�
h�ܐ��=�'��LL����q�v6�H#��@��ܺ�}�TAˢU�O~8)�>zmO�;a�	;q#��c�g�Z��q�!�9xE1x��x弥�nJ�t	/�б�U=��m+K�L��voT1�ە�E"zfd��/0*�0��F��[�5�����t�	��w�G?��_��r0Hy40�!"O%rȖ�&iD�g3 ��
E���kd]c�cW��h8���5��F��=��;�h	v-��~���&��8�fI!��0�>aZ��l�F,GJϥ˳�y�Z ����	!"$�!�Ϳ]I�����C�{c���)�#,.��3��^�%�1UÊ�ihʩ���6�]���5�ڊ*��N[��$#���`s�"ŀ��<��	�'�	4�a�c�:~���a���(j�
���k�JҚ�H6�HjM��ٷ˕`|�s�k����d�
�s�O��#6S����C�&�L���lo,`��|��}n��8�̏;�3��$� T#�1��r&�o���������:&/V����g�H`;�ə��%3{,Ӭ�f��ˇ&d��`�廝�(��׮f�å7�ĆϷ��C��m������:��j��O��a� 0���Px�݇3���5ׄ�����NL�$���e�~2�+�L�9T7�oY��H����~�Au˧Ǫ^�g�A�zϨ����Ϙ��{]�c��p�)��#{C2~O۞#^)a��R<ޔ����#t��Q�Ik�	��᳿��W����;����vg*�}� Yi�[���QR�Cz_�;>�У�O�܂m��C�;.^�S� �3^T7b5�o���U��:�}mF����e�C~9r�������~\ى������)�� ^��B/�'�k���W
�(��T�$��u�R�Kc�-;��0�7p_���W�*����:3X� ^_8dC�Z.��5�Ȃ`�-�uꍤ� ��l+��Kr?��}L�E]i�G�
JhV5��{���x�������q��\�Y@�!RY^J�܈��X`��6#"�ݳ���X��M���ę������C�������qP�����р��	ª�:8�cK���}�~����7`���G]�R�y	�Y��8����SWS�h�j��Xي�3b�y�V� f���1�S��)E�w�bG_��#�/_ .I���m��LYIG�lB]o0{E$?�#�u4��ݔ�r���h[��QBI6Fz��Ub����V�	$�koh �:�� Xz#l�D�D'`��.8��gLYţ�5��v���z��P�� ��rڍ
�����W�0�r1�(����N�R!�i�ۻݻӸ��2�j	��ƾLo��Mr/��y=֪G:�;����:�刘fO��2�sP�W�����(Ue�w����K6ۊ�Ul�yH�w��mw^e���߳�/� ��+��,+���M<H�
`xE�iΞd_k[������"�����r+��������:��]fT���+͔�&¨���#��	�0�����DV�fs!���M�$��@��m�0Ge��́��L`�_=�C|�
@�m; ӟ*Q�uF�R6�M/���e���2�%p�^�����|�
��*e��Ec-y�CJX��Ӌ2v��h9������nn�_�A�H9�������ț���:|8,li>���5�}��焦�0�����r��Z�T��05�^*�O����؅��W�q���,��<^�,��k��|ﺥ��V�y~s\17�Auah�q���[�؊�xe�Ϗԋ;u�{�L��٭H��*�1�W'�� a?J��x�X�\�8��|*�C4&�װ�㿣M*L��\���4mt�}9�B*�,>�)P�D"���g~�ܥLmXo.�rO� �,V�}�:�H��oY�"ʇ��s��j_���|�Ũ�	�����k��N��R��;\��S���\�8��#R�n�b�[q�>��5֠��r�� �Y���.��4rQufs1̐�����Q�a�(;H �geo~ls��C] �n!5e��qr��4��-;�O�/=|��	ե��#D@H�+�F�ˈǘ�������;���=�D�@J�<�x�
At����"�U������
��_�O�ᾖվK��'n�����Er^�K4,��J���j��׬*�_�^i�[��V֗���numu�P�X����.=�]>s޺X�cP�C�.��T�#O�=է���n�v1\�,q���{�LX�R�.F�GйR�d��u1��Һ�c�	7�h?��j�]'zg� ƽ#Y�FT Q�o>�JEJ���z�ѫ��U� ��� �q~��^@��1C���
�Ab�ۜ�H��f���(%��b�\�ױ��mڥ�3]''O�t0�aK2�p�@�X��~�1	ň6衯o%���S=� �Iul��@j�c4���䏦�Փ�5&I�2~�h����p�\�,�bl�1|0٤�_n�C���A!*�*�7}^xj>d&�)('�0R��������`�����m�^>"�d��F�)���F���x���?k���ol��{�D�И�w<�>d��O>��>�*�ܜ���"op	���l�X	EH�*��t��\.�����e�R��t;���W'���K8�b����s���N�o+9�|������_��9w��Ͷ1�r���0E3آ#����Gf���d�֗$X@�ݭ�r��,���L/��"����X���7��y{_�Wd�6������I�@j�ޮ5��*�k�v�����2󩺙��S>��L�`P4|��20S}'�+i'@�.ި�f��ЎIϛÃ)�K���6o��,���k�y���u��e���9��-�X�To%� *l ���(LE�����gڮa�}�OLǅ�k�D� �%�{jj)}f}Jѽ:
���$��
6�@V�3�*�ŐH�������	�Q���l����:��7��9�^�8��c��K�DQ��ڶ+L���KL��]���;��PP�ޏ�.��.k�a��� �q�|���+Y�����J��� ʇv�Ve�1,m�8�q���l1ـiz֚��(n:3zmo4�O߃?Xk\f
�%&��sY�^+�E>Nؚ�b|t�/�9�a��F����.�����5�0���	���9�!{��=|)�D��Q�匮�5� ����!��]��S���#��H�㆙��}j��,��cI�/���v�@��;�Bv~�[�x�]\��=%����n�<����w�5mi�j��TJ�Md�����%��+T�$N��H"�B!��畨��.u1'�w%_����r��sX}0�Dq.����Q!2e�x�C�����6���m�YK�z�~$��ꏹ<w����]���nG��@lP`��;�&}i	�n۶.���y�g��1��I5�c���]3K\F�|Kq��^�F�H&��VJ�IΝ��'pD�&��4֚��,��ά'���*y(���?(ߒ�5[��<r�,WR���X^)M٪�P�^��,C>��3=Ф��D��C��JFck�IG`ک 貲&k��%�C�`�:��d��R�j#��G�W���{I�V�Ų,�����G�̈�I�г��n��f�5�#3ɢ�Eи���8N;%,("�rW�;�X�	L]C��~U]�� X��v@�������R���u)#B)��v�D0ŃT[����7*���Z�9��ˡ�h�h��z`l��?%�6��UIm)�C(���wL��L�dŁ���5*�y<��n"�Q�R8Z4�����*���ZV�3�j �5���������݅�ѽ_3%AI��LF�E{+ܖ��u+p�A�ﹸ���g4�����_��^e:�Iח)���^�W�Y�"�Ӳ���z��K��&\���5e�x�N>;���1�!����^�cV5y^%m$�-���G2��gӳd���w"{���]���؍��R��J��΢:�i���Cܲf��o]\��ݕ�5$����P �5��Oz�F�CV���v{a���i�}������M���M��٭�#�����'�hNk��O2`$�l:��G����F\.�C�H.9
��րW �`��u;�_E��*�mVt>ݯY��#XΦM[zJHdł��ل����8����M��#�Y�Gh@̅�#��3�V�i���G"�3�t�"c+�������1V��߱�R��� }���_��(�7/<k3{$s�0�?�H��b�]���i`��>��|U]�����9���oU3g��c��P99RN�@3Q��ά4� ̬��Fn���3maQ�,
2��Q�eDw���ڶ����Y4,�QR�}*{�:~PCp�!c���є�n1���Y]�t�ޢ�P
:I��i�C�Bգ(�z`�)���8 7�9��i"ǷMlG�֑�\7����y����Tu�A@V]ϐ�9z��#�`�<PVb�1��� ����C�{^a��,��p�^��ΜL�+��6��4F��^1�AE���BJ���r�e��Eg"���(��'����ԕ��@�8�9�����z,0m��C�w��)s-��wC���8�贳����;?�}Z|������5zڄ�E�U�o�΃Z���o�`�ϙ+�;M�j���g�5;��$cN)�g�����ӂ��߲%���_@b��i���=�D���"I������ۻe�ٛ�P���P�%�)Ku����@A5X〄���L�+̞�#ەH�u1��ׇ���,_@G�G�[E~���QI˛9��P��1���N@�X��_=i��?U�xB�OC��$xNn��NRT�8��Щu�sR{/��9����#��5���b���	�ƲC���x��4ȒG���,w�b˰  f.pA�̙�%	W��Fo��ē�����,���� ��c�>���Os*u�冞�/��n���mb��6eup�Q��� �(s��M��؀�(�^|�ЉK�"���on�q{�Q�����>Y�ŵ���|D���$�Y���lӢi�2�YԢc�U��>u�A,�5�0)�`P�SV�x�@ʓ�O�������	���,�st���V��6Ř7����0�g}�F�[Os��T-�6�]A��~$$�.^�*R��� ?5N�m�C�wī��Il7����	yB�#5��4:#a2N����7������r��.U���_�y;V��;Z��|2��1Er}�.�)]K)s��l��_�Œ[n��pj�	�D�u����Ԋ����BK��cף�0#�L8g+Yb	���Y�.n�T�N>#A-�h�����buY��SB�>O+�rgs��6�^Ġ�˽�fu�r�[U���Lh9��:�cA��|���Mv�qs;]3I�1�m�<���=��\J���A�F:駠A�Q�$���O�	��Y�,{����͒���	�Ο&�- 5յ��ʶ�\/��j�7<QC��y��3�X�� �j�F|.�긏{ch�Ɵ���EK�k����E<�B/*���Ir�u���ЛVX��qV����y\��b��O[�8fz�o�o��r}>�\.�
-38���?�@l�d��8��Q|�+c�"��з&Z�P�ro��%�{�Y���i��ȧd_gP��%�N��=[����&�};Y���Ύ��f�y }���N7=U�oU��fRpk��$o��?w+ׂ_v�>xe�xTw��c�y3C b́��w���{����w��zA��\"�������K\{�=�����r�:�X�C�DpVp=g��9y��� ø�T"�S�����>Z�� �JJf�FGjO�Tl����(N�4�k�g{�ҟg��<_�x�)�.K
��s�:qr�|Kf�nZ��;X�`Z�S����ˮ��u�Y<y+�^<rY)I��P�E}ӕ�P����Y�4b���5�����R���n��M�" �0J�����e0�0)�B(y���7�4�PMxT��'H����q1��J�=X�r�0;��A�	���C4���s����]�:�����*���/��O]�f02�������2����}w�e��:��Ѿ����Wެ9#��z��a�̾�Ax��q��Y�$���w�2�mu��D�QtE,@�[���O٫������l�;Q��,;�ֳow_	˙��~��'m�;��e��`��cB@�UAL`�랠}V��P`�.sq _�%��0��uN>�#S�ʗ{�ֺ5�y��t81K⑮PB�k �����h�C�E���
4���<���֒�XQ�KeLSwb�w��1�l�[椑F��^��kxP�4����:''G�ܫCF�qH��넖�8�<�'��쀓��6w~e�����ĝ{e��z��S8v�p�k����F�OP5U�G6� T	I��ĳZ�,��5�����R��C��.ܵ�%�as���FiP�.U�{�;�V�%㾚�5���%��	�{��k�����5M7NR�t���� ��&g���s�	w@3=��P�a���J��K!��z��4.ޤ�=K��IS"*�:�oG:FpsPk����������Y4�� �ῺΓ�M�_>��o�l�~��5�F��3���=�ޫ̑��܇��b�m���1��HR���N:n���I�B���F��̦�@��%~��q>O��pX���&�6A3
�BZ!�qǕ��)�(��o� �r��yJ�З�L��>d�ɒ����e �8��ߚA[zƁ����1ת��'�ㆥ3h�f}꼡��A�W���C��ͨ�l6�l��U~xLe��C��CGnIy������}A}�^7*Mq��xQ��Q�
E"���Hr�{m_��2{�ҍ��n���P̦5�v2����~��&��^ �y����#B,�T4A{��DA6u�8^�O�5`KçPvU�N�ǐ �}��	Hl��b'G(e������K3��o�+��럘\�.ɣ�����4�=R�TN�.����*[X��z���SL0ҿ>����MhA�I�F��ہ��ЧQ>�FIxlcAC���꩝u	�Y,9wMZ,�<��?~�=�Cpu'�q֔O�^��n?��97��	�4�LZn�*i~&����Eߠ̙3E��_�t��)!�qХ���|Bc,&׉bkA�$��W<S�d���)� ��'�3	f+W=��(���9�%i'Į���z�,0�~��mqi���L��`�4 %�@���R�=��c ��5�`#QX�0���M��"�I�L�4����Ft�^�n-u-�g����bR��L��Iѵ��vƴ1Ce�԰<:e�s8IJd^�h�4��fF�0Z��n�,x�h�����_7���	7[,����%7@g��A�A8�M�T���j��,�Ii^�Σ��%����7zk���؄�'��� �RAH��ÇLH9��HS0�G4�����{mHO�]6q-����ΎT�k:4�|zi�ug_a�:�!� P�n�`!>�������_�&d`d���ct� �O"��/ �����B�{�6�TX�}"��=�9����Z6&G��K�Iɍ���@����>�8�>H��o����G�+�U�\�jn�l^8Ǣi�g=���T_lJ��L��G>ӽy���8U	Uwig�� 3"��h���=�#���h 넠Z��T��4�/i��x���9�GܥL�ޅ0���6�ŭ~qD�t�5���K�����"A�h*.b��{S�s'v���]��	 �_��Ƚa�J|, �X
D�V7��#�.�c��O��K�ǡ~����̲���(ݘO�#
\+(eH�����>�L�6mS�!��z����zn���4*ǔ����w����ٿ�owI߸Ⱦ7ۇ�T2����;@����Ke,A�`�˸�|Nr$�q66O~�q1 �CgP� g����Ӭ���LX�.�<�Ł�"��d�`�Z$}V��ym�j�:}4/��r]�fy3x��>TT������SM�m�e*&����9�5A>���N(�	�'���5Pҳ�bX�c\��ҥn����os��\�_��T#�5[�{���3�)�k>�Pͤ�w�p�c��j�kG�v2s cx�M��'�JT�mP$anjb��A�N�$|�N�swT�#׾<}U�Fd�J���8KWJ��ӄ]��&It�2]�p�#�~�����\5�`������{0pUB�A¿!h�<j5fVb$0 R2�c׈�yj������.Y�����Ӷ�1	W!)E���609L^�T\-��	G�vo�/
-y�"�0��z�J�֫�٧s���`!6dP�R�4S���D��ؤŶɃn�ǒ�9�/�h��'��S�\���N�����(V�7/ޓ�~~����P�h��'e����e����;ro��/ǅ��qޭ��AT(m���cR��]"�ْuHWj�Au��j�hD{��i�,9#Ť���
&C��Hʪ����[Q���YW{�FQ��^�6��&��Ր��e���'lunH]oz�@*]�T����]K"�Ǘ��`�z�:,���bza�=����F�\t���v��B��t�l�B���m�dUm��[�Ƨ;��ݕ�f���ꇭ�}��$���� ��CZ���p�H���	
%�\��}�c�.��1�\&?��ĩ�j���x��d��
�-0�h.{X6"O����k+�o�������O0�P\����I~(u7��,3F�>���+����Dd���Aγf���`�N�ʋc֋�O�j����l���+�{�JRN7���\|�(�
͜�J���_����f\��.SY�=�<�s7u��KF@/X�>���W}c�R�v��0�����C�.���L��K7�Hgs��/}�����~'�>ה�����-��<>b�	Dt�c.�Y�\j�}WXeșސr-���h�	ۃ��s\���^0hp�WT9w
���@q��P��-�n�Q�<Y���Ѓ�䣲��������xȳ�gz���P��lR^��S�ۍ �
lVAI���7[��Y�@�D��ehV� ����=K7>����h�k����L7^�h�$�M� �-����{�*�j�����v��L.&���>�ŗIݦJ�v�;�|��>�UQ��[��e�I�f?`r�����N��d=��֝�N�V-�s�Ҳ{3��W�v�l�!�� ��>-����r&�^�.�Y�-�����7��
F��g3�f��`\(66Nw���,p�X�����N{/�{�����\�0;*)��wAbF�cvBY��h4A���/��}��+r�, ��q*Ü��s�X^Ȩ}��7��O��9�zR&�2��7�H4žeʡ4��f�z�D�/p6>A�V!{�Q� �x����h*&<�m�q�#].���^]@B�DL�KG)ѡ��	$�9��O�F<T���T��V��<vS�Y��~eU�<� �p�U�X�r��<�@�čtt����(q��U���G���E�'��H'���$��Mk�y^�#�Kd՚1O���f�(;�%�8���'��Q 0�&�A��IS*nm�O�s3�:&kW�dGN[t��O�Y�ݸ.�9	X�;m� ��+,ü�,��]��LL�r�M^oߧ�a������?  ��H��r#�3�*�w@������JF�f�?=U�p��/��5K��n*��&6uf�=�6�уX]��nN��	����x���b��q���b�]�<�����7_����bc���j���F���"1���e$��+v���y�#�Pv�Ĝ����\����}�LhB	���J�1�"дdܗ�y2Y��~ds�����jd��0|ef���HGև��f�
�wŕ�?�!t_e y=�Q��ܻ���A ��z�s-M��١JU���A�j����3�4����\�6�YT1Z��s�1����ޮ(�v]��__�T%�]b�����NQ_>���`\�<�?�=\y���rN�wd�C=4���X����mP�e�k#$�+�G���b۔S^:�|���	�|�`^v��>l��(�)��E�Q��0�B˰��y�kM�]$�.��Zl@3���P1'�@�&���Z��^��p9D�1}�,�Є����$�0�˧�2W�h���8B3=����å/�O	c:�u��n!�\0�:=F�O����o��QO[����L������<.KB[$X�q���X�o��q�����Đm��,�K�q�m��Jl�h�_�w#��M��� %��;.d>'0?��D�����?�Z�l��,}~6/�� �k��-�4b����xOd�_w4���օ�/�z���q ����/�7c5��'�d�`Eo��������Dk���42[4�יhmAn�m����S�8l��
^O����}&2`���W�S~�	WY]���]1VTc��v`=>a�G"]��I�Ա�s`��9�	+�P��#$'������ 1�kB�G�ə->A?��S����!Jk��f=9�!\��_�+�!%<���|���cҵ��V�C����b�z?҉H��txYh��U{Mq�^�B5q �Ih�Z�2�`%{�NϘ�E�R¼)����Wy\)���Tl-$9�;�xՖȢ� ���5>�;S�~O����d��f�=�h�!W��Ԁ7)�m[[���H�]Z�S�L�3���S_p�Ws �.)� �k���$烛m?H0+��$ڀ$w��n}�e1�W	7£�*T�#���[njJC\ƍ.��n���6�ӫ	n�y��@�.�&�>/��
�(�<��E�V���d.V^��� �u�@��pf���K���>����؇+�dz�jB�D>���;jr>�0�VG�g��u�o����{���ަ�G������0c��3J͒��G����ΰ�i��=Kk��C �5�_��7_'�U}w����5~NaJ�}����9�1��閜HMS��|���xXV;*C��y�c�q�J��)_QXȫ�Gd%�	�~�6�����j�k�_�̯���]�>����y墜�+�$���z�7_�� CK_�o����Cވc�+�sB��H��}U�!����h�>#T��R��D>	�����G�b����p�"�/�oo�����'����-$aZ���
���������N�����ƞ���JA�I�$���Q�(i�F��KL���v��f�唨h�>����9�+�[l���O���vO��q5q�5��]��y��;Y��`�l��VY�oY���|=F�eX�=�̜[�����õ���7Em�#��B�����Y�
���ݤ'j%�V�SfU@�:׏4$e�jlYA��߃P����"-�/<.����� �0�}��GÚ�+��
�%�^�
sC��4��n �y��UP"X�\�d2������2�o2��f>������Q��Z�Y;�G0�l����F�$?"�qھ��kq"je�~��Q݃�?��ͦ;Nm��\1� KhX����c���e�v�L:):왥�� �����z8ѧYB�V�EK���#M҉�����|tƀ�2��SpL�+#ڱ5*i������N�s��E`f6��
Kɢ�E�H)���3��l.��;I�V���a�i�:sDH[��P���$&t��pq��?�/���,�.;H��ǑKSk}�_�Z��KX[��V2�Q���V�l4���@X����"A�J�_3��n����m���h8�<�N�&az��=8/���r�����	��k�y룏>�s�v�!�w�K�xV7��%ܑKu�>��Aq$�
2������Yh����H��D(���w-�TC2�Ҵ��v�g��0f��I�i�տҌ�F���=~N��6m�����6�:ﾼn\c�����G�x�:��O-���uDE�U!�{1�A@nI��E���VMog�ym�鰝��� U�x)sBW9\��i\RH��Vy���Yd�&���4߂����j?���)4�<!�Cyү1����%����	�gW�UvcV4�V��=�/1�f�ު>�MT�sc�~aI�0rE/��Æ�s
M��/�#>8�����}w�_�cW����T�L�;ܞ�J��#/���uS����)��2f��D[�x�
����D;iN�^{�Ҫ�!�d�gLS��%�ڱ�HU�<�N�5!�����0�.#7��5��H�=A�Vy�Ep�����pL*i �\ݟK}0��A����E������#�WW�(��A��j�B����G'\�kV�]uv@"S&a�h�IN�����5��'�=f}�~�}�6^M�w3�ٸ��ѕ��v�y�x�Et��5x�\z��W�F$R�Vos�i�B���"�r���P0��X���[�8̶�H;
"]p|�&�s}��H���=�9�!��QG8�I��T_�M�6c�	9�Yu�B�P��k��'8�"�<)�9�g��ca�aS!�{���o��,��ƴǑ�f�^��	 ������^JE�����'��0H�o�����_K�<��.=r-�u��.�~|S�9�>Ȓx����O���N{��8���3�3(��"���*o%�	��H�=	��!�}�v!���}��ә��		�k�ń�����i�[�Z�]�Z���,��͝�N�iw��$~�ܡٮ%�'�Q�Vicݺu�P�$D��w�\c�Z�Ŵ�I���$��]�[��w���c�'�Ge�S��m�*�8yDIK3��`�lt���B��|�`%�S�����76�T��:�
:z>TW���/���Sʵ��E�ھd�i��,&�8��̈́�[j*E���9��G���:J{����!h��-1B|�������\��%�?��~�IB�ָ����a�'���f�~k�n`��-Q������N�#��O�d�vb<ޤ�,S�:,���9���� C��C�E�>0��(�i��e����mQ�=���c�^�\1t�,d{F��L�"T�I�����	T���d��P��r�)��,�lD�532�(s!k����J�t������S�R�n�,cHz&lO%Y�Z$:E�Ӌ}OL|��6ِ0�����"�^���%����v����%X�6%��ԝ�R�vi��I�����$��K?�+�m��e�eA�kĲ��m0��9�EN(Zη\�8Գ�@�QB�fI.�S�
`����׏�8�k X�)`�;�58��G>ϝܳ?i�*��(��ji,�2��+?zu>B�W�3U񰨹�U;g���/�I��0&���֑�K��7�˾x��1���߀��w�W����� �eɖ��׆Rⲯ5:�:ڱ�_����aӇ����h��e��XX�wԇ	K���?
����̈�7���� 4�����Y�&��C�|���ФY�5�Z�?��u><{�o�^��+,����?���,�<��-��sڪ��:��M��(���}\��wy�R�gP���Ơ�f(�A���</�Q���Ex�����\	��#(�>�j~���S<0��-�2Rc�m� (ds�|���5�'E��Z�ኞ#�.ُ[vz�z�Y���w�u֬�����qHM=1�{2��'�Ǉ}�p��QK��Y�W�ſ��?�?�$�A�����tZ���Fr��S�N��$TrX#�?'�8���vé����Ѹ�i��$��Y�b�����}5�@�&<���j ��~�z�+QjN�w~ ��j�f�|��9���ք��B2@�O���WB��r��T���64g=�'��>E,,`����"�`*J�B[��ȳ�&� ���o*�"�b�Nߗ��@���G��"���+)%]6��o�Yc]*�hi�&�o���s��!FYh�O�V��W��=k�	��&N�>�g�}ʞBr
ʆ�1������@�u�A�6OD�j	%�>
��*%3��Ϧ�>�m�f��[�<1'*�3ޥ'��Ҕ-�ρ8��$$���v��E3�A�7�ՠQ��_�.�&������$tk�%z}SķȠ���yކ��\K*+�ʳU�K7on���MM�U�<|�ωY����*�$���u��r�q�N��n����8�PҖ_��0"ɬW`�SQ���jl��f>�����0\@g���f@�KB�UE�γ���<�~3Nd��F����7�ƾ��h��k*�p/'Z���b�J�$4��:K����Fm��������xB��fR��j��)����KƳ�/2Ҝ�����nON|3�������7Y�IM#%Q�Wgx�<�4Z%����+,IUV"�a��Ќ?���g��w\�F�kP墌k�nF���V�ިy�4��q���s�b{��+�؍d��9�a�|4zCeEh�l�m~
1��2�qn<��^�˅�N���gZ3	w˵&�?���WI�9hw���,�F�D���J���c`�%�f���׈64��W�'aA5�u�aq�+p�vc[����ke�y�����#Er%�[f�����b�_���V�aG���ǌ��H����V6��%��tѲ�#�[;�;��Bޯ5mJ���:I�$A\v�.�����X0i�s�T��6�c]���x��|���b
ɮxU9k�W�ΐ��?��g�K�M`��]���3��	���H�[(93��s�[�IϘg�_?�R�)0c��]��7,�T-�Maao�72�7+$���A��F���?��&c���Xx���*Y/u���B�䘾G�� H'�lm��z���b<�i�P�i�ejx,�NB=�rY�k9�Y�	����;����ۤ���~,������2r#�4$�z˥rPE*��(T߭q�6���]��{c����	�Ь�c?[�ʹ� ��UÏ��lf��z�L�΋L�<�1j�/�>KKk6n7��Q�"��7$f��w�~��W�o%i.uYӜvTy��/�=Jcn��`a������a���w,��W��]S����?/ڤ���[L�'����e�YV��x0�M�m�bc��w�%`�_v����':NP���qE��+��`V7M��_�a��T��I� bn��H���j�X^?�P�d;j�do��\e^�)�PH��lpѴ����?��=v&"@Zv�L
儶r��)Ӧu���c�p�r�,��IF��{ՓU�/������qW�+�$����"^��[�.��ư��	�t����a%a�����R�S�����n���h3�@c���x�z2Mʴ��\
�>:
@>��F�����N����-ŀ�o�;{>�
�g�ψG�BXso���3��
5�Qir�KTs�K}"�!�;�q����������%H��wdK��WC��f�]�L�����&��A_��7
.�Z��Vϗĝ?��ī���qyGz�����k��=�xe��A �c��=Ae�T:u��f�+�XrC����;`��%���Alz�*TP-I����"�d����E�S8H�����]��E��]6I���մ^�[���*� R្J���8P��}{����E�~�X��./aGф��`���.�ϹI.2�A4�
�����9�U����q�qJ|���휞FARI���j�d˹�XȚi�o�a��~�|V2��#������F�U��H�����U3|�Q�o�L���=�� ��È�cV8+c+P�v����f �K8���6!L��I��S��wĕx�,R��iq��;��ԙ����3���ݦ���U�,5��!�s��j�C��z/�<( ���6�b|�m��-�U��͠R�/��x�]��
�*R�%깵|���Ŕ���_�w֪�)ӈ��RN���ZK� }���8����p�����oH`�=�l��Z\y"P���\��e��+����uM���D��/���
���8���;M�_?3� �t���/���2��f@�L���[pi�[ƿwWڥ��aɖ�d+���,�=��� |A՝�^���2u�ay_n�1���9]%�j�,��ԥ��찖[%X�$y ��k`�ЕwѲ��|=o�	|L�����#���i�8���,V^ÿz�qy�f��e�G��w��$��ܮDt�H����� i�����E�i0.��1NI�.,��+ ',~
��Ek�CB�O)��i؜�rewg��e�#��a_���ע��I�Ĳ�7�L]qkڮ�|��Sz��m�Ʉ�G�80Bf6RS�ٚ�!����~j�a}�y�l,TU_z?PԒ�*vy.���x�L�d=�b
NO?kk\ �Uyo|��f�M@�VM���59l_���A.[��!&q|ԟ/�NL���W�[l�w(�p
 ��$��� ʹɨi��
A�Bu�9x��}D�1`�W{+�DY�����J�	7
E���^�0:�q�3�x&��#Z�;ŏRU羗%wu�S/r�p�64��N+��	7z-�iPzK�`���Xl�ȡa2gb�����ӹ�^�æky$݀6U_BY�TuS�Ր�F�[�w�����%�\`����Hώ�>�9�~���$���ɳ����� ��j�k^$���P���Ќ�#�k	��ѓ�Q��&�􈞸���/���%�@��؇��$�+�F8��PY:���ͨQ��)�f�{7���l��-7�l�oԼMw�[��{� }���n���!+�O���_����Ȫs^�nߐ��)�� _"�qߒl-,4����klw#��*+�,��>����s���F��{m>Ժ��q�L�j�f�<r�hD�t���f4p�����T�-x�`� oD����]��鐞0�Ӕ�ؤ��;g#/{/ �~=h!��n����Pv�._�%����$"N噁M]#� ���i���<�T��s����0({�KP�Zj_#�dw���	��?�^���oÞ��%��>�ݴ.T`g[�R 0fJ?A��Se�W�.{���s�uM���� �a�G>8�L�1t\�X��s���:1E�D ��p} Ӷ����N�ԣ�׸: Ϸv͵�.f�C�E�~˭6��Q��AY��
c��n���U:� J�H,�igݎ��mS��h��S��dĴmE~ma~�[�}l��#�p�Rx�ڐ��-�f}����8q \�яb}�9��.��9+�;W�o�J٤��;WU�	U�N,r�������z�=��Eu��Q�j״�S|�5Yk�1�%�����P������Z%��}�\�Cu���P�:���~����`�����gآ����Ī�Ww~��mif�$ك������I�HME���L߻-
��	���B�z�J�E���KEV��`�x�4~���2�yʗȅ��p�:�Մ��$�)^Fm�r(�"��:�b}�&�򺬂���jyXテ�z z��eOŅNV����'�@�i�:�
����5u뎱<t��JpI��_�x�Ӊ��2+K���u��/���L�����U�md��$f+C�$)�ҙ�������5P��7���\�S�4�בU��lƅ0��y�<�� Xh�tJ�����bՓ+�x. t *�u�!9�����xP��<�����"3�s�;ᅂ�붾�����,��[��s�{_R������hڏ��|1�$O���8'��B-]dS+h�^}�C@��r�i��ꗰ�Mh�}�>��k�,�H�Z"\��p�ف�(�i%���r�ht1�aY�B*�&���'�:f��L�U;q:�0frl��k��]
�qJ~ASP��``}D�#>��9z ��U
����Y�p����W��rݳ�ȗr �
b`�O�ޝ$�i���,�\��&����8��XcNαmVe�4��@*^bسj���g-fW����f��]]e�ѵ 
k�^��Ij�Em�b���v��S7�����0�[��� ���L'���a)��4��?k)��X���X�^�5�"+t��S=��pMT���Cw�`ī�7`���L7����|*NP3?Nɮ8�J���G!s�@#Z��o��1\w�P~d SB��e���J���4�I����Z6��>����v�.�61H�6Ag.ⲄAd�L�:�S��1����A�󀼘�[���&�M���&���!%�f6��<.p~g�롽��D��z�]�)�chs_G���}�0k	�`��b�����$A@�� (��h�����1�6M׈�j������f~0U��[��@���na|Wm`4_�b�i�A����+�$�i8��JNn�m��hZ���{�ה�fU����Y)�.��u���G��L<658����t,����n25u"�K_2!{2�l;��y,
O>��D�6'9i^��k�߬���7�*c���LwHK�ަ�Q�'cn��np��a�Q��0O*	ȅ��UK]DEkKA;
���� 8
�b������/��:��|�i,��rt+�
]n�늪y�[&�=�.4����$ljYS���4���?Zx��HR�}��A�h�~_�2G��sxS�q�����[�*	3��^����EؚvbR=�"iz�e^,�Z��a�^3������ފ(,pjW�Ív:���K>�������*�e��oW�;Zk�`�����s}��$�w<δ� �Z����׽;7ސ��r[H�7^Y�ڣ��LǰP`�҉$�d�$���b_���*4��e(ۀ���OmI�l9?_��=������\����h�*�r�_1�\�;�������jiSh�����^�^-���}��_�"*�*U��Qf[;���oQsb9�}b����������p�2[�G�1+Y��[M��1Nd7��1I��3�B��E���&k}82����,�kx9�+X�q�����^Q�Z�����Ǔ+|u�$6�R��1:S����'�(Z��[�fW���A�D|� �G�Z@��vR�.T�}W�5�Y�i�x���|ߴ���5L4�%�bXvY��_ARw����̅L�,r�1Ի�$)���������%V�=���-[���~Yjr���Ëh���p�"��w� �����,�
�3N4��ƜX�e4��_`�3�X���j�(B�2�n���	��}���C��瑫������\� �5�� ��,��(�S�p���"
Ɂ���Q��P�~�4�y�=��5�C������M�a�r"����<��Ė�b�����/i���*������cW�hlE0],�u�wn���D��j���?<�X_�TuT���"�K�+GT!t�07
9,����Y�%��e^��Q�����f�9ݪ=\��C�~�[B�������Q�i��Nx_M�>�r��, Iyϡ7���#2މ<%�-`Y��j'z�T
./�#Q�i+D����l�;���7/�m]@���/�y��������a���~�v�([���"��U��� �N;�f���$`�3�8�w@Vz]���m��I�e�Ꟊ\+S-Ĝ:$�Jws<�b� = tr Yhw�Ŀ�<	�������Gk�
!i��(���:�U
�! =u��y+�[Ƚ���ݎ�)�K�ף*���"�88z�u����ƲR���/�kǆ�r}[�Й~Jp:&;r8��g�
��%m5�-(M��hm�\a��ԭtD�"��q���$K��|$7�Q$���KzӬ��p!z���~b�W��Kj�q{Vic��|����K����
�%�D��7Jq��h$�,a+aơ3��ڑ��*$�Vc�������]�	6�m�o����HG�=8��&�6f�,ނyuH{9+�=o�$<�^d~�d�)���f,+lnd����O�׏��k�}�����L�A�>�ԶUL���j��7��율���;:�[F^��!�|�<3��>)���9Ԓ�0�uY2������;��i�p1f[���-���Ίv�r]t��5���l!�Y�rj��n�ۻ����e��΃+��-�I��<�s'Q3[��	Y��c�Ӄ�o��)��~ߨ�_��U�j�L��R�x�����9�]9Ds�s���#��a�`�#j��H��YƷvVS�F��ES�P�gV�r�r�F.ɍY�����;։0�B���>���6��o����Ƴ����C��~k������=%�=�XD}�Q�E]^Ɯ8��V���\N����2��.�9R��˱/A�>?Y&�N�O��xt��7�#�mm�9ּ�U:�N�,ֱ��2'~���dZ��&Wv� G9�0+��@mw8#<:Nu7����E�kע�	�6�Q�622#`�H���7~s��I��8S�:�?!�@���
1��`�0�R:�d����:��DAa�Vv�
�B��Yӏ$�ZCOa�}��.
��/P�f:5L;�����W�^P+�o��(n�#�'���V�1>c[ٰ��7{Bv�Q�-�WC�/�}�_�IWT���\&�w�Yw���ԒLS�'��m���=���e�󃗃�7�׹������^����
�w�/�)��6�j�B�����q��2�S�v!�O$ ~M:��Ů!��1���*����zSQz���Cɜ�_�B������u;�4HW��M�wh�6��q�V`B8k�ZҾ��?S�t#�����{��𱕬��*M>(eG�>���6�v�ve]2�>Ҿ��+�Aɳ�����������|��D𿯨����hRg�Z�����Y��x��������7�ϧ-��\��5@�W4$u$�t �	�#G���F�L���(z�9z�bs4���nA���q~�qq%��/�:�~�c�N5��^��o��=�K�o��_��)Z����e!n���`$�/a�Ίb���]=I<�?p�q����b{(۲�5��ָ�$.�W"�s��UZ!��*��b&��K�n�ʪ2�@cTܦ�Ԃ�{=.���I�jޒk�0��`�V/�G��R%�w��'z��1&qi٨YE�[m&���j�ݚg�ʦO3����Ђ�s�zD�Ɓ^�����Ni.h�Ç�/JԞg��X�~۳-��Ϯ	�*���ץؔ��*,2�^ٳ��U\���)H���#C�<g��h��,��(!�]w�k*<$m��&$P�d�H"�Rhe��y4p�ܐ2���2s��e�� T�ä	@蘵9�Kd�����'AX4�� ^��-�L�aoM4���Rc���'�al�?�o	�rYM�7Sd�L�8�ma\|OIY���D����2�E�nw!�L}+�GT4Y�3�_�4��X9�?�!��N�zD)��'%�>�|�:�_��|U��%��
���<s�[H�*���fM��`U���:v��ۣ�1�߼2%��!��� �� �{F�F�=o+���y�)n�
*�)N�����4�Ƶ�.
�]�}$�^���=	�>��R`##J��j\��J��<ξ��Y�7�ą����ג�+�w�~��%������AK0roXo����8�X�s��#�6�ڴ�id?�
���F���A� �c9��AEj���/G�!IZn��R��U�p��Ȏ�4��,A�ByL[�!�pN���6�b*5�D��1���c<*�������	䚢�I	p������i�>��.y��EU+y{���G�4��ڢ��%�}y�E���^�O�n���H�M[��4d2�*?t���յNe6�L�FC��t9��Dq8�ۢ֑ɆFo ���
/!�I������6\2�.��@�{� ]�i�����}��3olU��^��J���|���4���idv���Y[���~$�w��"o�B�u.�%�?������$�4Rv�گ6�6UC\�nj��ok�b�P�'fʷ�������8̰%n�%�� w�w���7�Ό�`Fi6&=d�;��
Ӭ/չA�����Q�Ub&wC�೗�LnX�Dq�P�dr�6�.�NF��%ib�Ͱ>0X��K��Kp�`��5��v]�֌S����6��ay0�Boh~�<΢�5�*ӓ�$ d��P�͗��� ��{�Edb٘Ka�#�ț�6���z_}6�(��`��#�ض}�^��wH�^8���͈}ѫ�1������:���?�}��:��Q�U�A0��%��~�1�V8���j��:[;��ҧ����3���܏~b�{n e�G���$�C�̃n���赕ܼ�ȍ���MBD�Y�J�̾�N!s�����#�l�� jOH�g	�ZOnU�Kp{���_YkC�=`y�u5:��w7iz�I��ƅ��[�A�;��U��}�V�V�ykg[7	�1��ȗs}Q��s�6� ��H�����/��?(,V��Y���Uك_��)8H�ax~��%6�n�K�o���-=2�K�Y�l>-v�j;+�����>�1�J]�yn/������[5L
vyr���������x��(!B���j�a�����~j+�"���'�{$��#��葨�6�����?���>xy��E�j��	id4ygH���a��6�1����b�|����IU�4�z���*F.����\�Q�^g��CΦ��]���8�_%�D�K��J��-;qw������#h)F��[���t�WS����o՗��Z9ۛ}�"�߆A�>�g{��c$Oj鱩s�����	v��>=�5An �`�u�v�8'��o)!�����Y��Il��aa�]"�)�m�65li�|���1e {�[�7�� X8�>�}���2)�a�&�Y�%V�a&�s^,^&64�~��Nn:�#;y��L�>��?����F���vYHr�֓�,Ϗm�y�D>D�2 ��+����'.�{Nx���F������ ��Ρ�7�T�v�6gZ�S��r��`�/<)�W땏��$�y�U���#Ct� m�(�Dez��q ��D��iN�BFk�jHG� ������Px��V��Ϣ^��/I��؊@���70%�n'���,auv?�Y��K�B������0��u���;�bǳ�ι��[�Q�f$F��d�	z~�Fa�ؓa@�c�	s��P�{];y����������˃�U�a@W��e0����à�y4և��\�h�e����͜5���F�gj�,1����2����c���u+7�oH�U��%rpQ����������u�Z��~�3o������@��2k-��ш� ��t �?@�̫n询5[lԚ+;��C-P� ��М}֠�1y;��1��ic�{sv�`NH'`��~qQ0���14�sC��|��T�/���S�X{݄ȝG.���qȌ�3ږlE,�A;.����<�vԶ3�v^U;�'��K:^w�٫�h�N:ǩ�Xfxp�l32itdo3R*�<��U~�Ǘ��p��1B���SD��ַ����VU�?��§f�y��4v���v ��NUg��Z�¶�n�X�\T�ě2qȝ$�/_������� ��M��حy�p���|J��]���]��|^zd��J>��n;�WaO9�m&%���{��|Z��\�E�/��}�/M�(��WT��.>�~��I�菟�|�MD m�-6&�B2���7L�ȑ��mv6��]���O{Z�����4�ґyȅ�;	1�p�b�����c�����!�W��֢P��"~�<�}mv�Eq������>�(�r����o]D$jjM�i��8#���/]�W=�}�K�'t
�Iy������m%(��ƯZ����H���]u �B�����u��\�L��^O�r��E\����y�ū �)y�Y���6�6�Zy
���֑������Ľ-˂U.82	���%y0@v�vK]����~�S�F��gj=�����@�u���I[U�6���@.��GDMl�3�,'vU��T��eP��Y�� ���`ؠ�z�J����5ñ!8��kE)!`�7�� �f��O�F���:�Ծ�<��|��Ve,�ɰt�v����g]���7Z�i]�`:e�Qo��;��=Me��e�g��:Pڣ�S�J�UҡG�sΦ�ddN�\��L��94K෌�)�U]�����@"~��}k_���Z.;�C����5��9N�|�-͒��`>}Q�Q��~l�AD����I����`�A�J{�u�h8I/Z;��5�0%">Y�3P��ca���+e᭐F�f(���uڷ6���w3u(��Y�&E�l`����t�z�
x�M覝����P�,���U�oa-@���7�w�h�&���Ne�&�ò�iw?�қ�>t�FE����j�M�aƮ���y
`MQ�vyhp��K.�eU�CdP-��9�x`�6�9	������ε��Vh0����@*�~��͜Cz��~�G���*šb͆"�"γ�J��2�0�e�FP��S�J
8#M�j!��i[�ȳu��m�良�~�x�Q%8]=���dvA����zlvN�|�-�}	�����w�o&�/ŅMj|i����	J�0d?��
�F�P�\:9�t�ٿ�x�;oY`�����Lш��ޠF��Lt�_E��(LR�����|�'���;��*��4��-8�i�#a��̛�]�R�h�ޒU��zD/:��j����6O&|.��f�L�s���:��fgr�QpA:T5ʩ��]�C��NpqW�50��).�K?Ňث|D�q�0$>n'��t�S��7M5B��D�X%�7B@Mﾧ��F�9������w�Z��l̓r� ������f�k�?t�]�� 9/<BdOf�Qhψ�"�^�I�3r1��u�V��#$��КB|a0���;�:w���}�����0tF�IW=s�?�{�mv(�j���GoN���2Q���ǡ�Խ��'S�#63/Oi��P�A${KD7	��#��h�rM��*|R�-�W�,�m�y�N�!���\����#�@�^?႖,�F��Tސ�e���Z5D�t�}�_��m�نP��P��1"]��k����3�\I?��rݞ�f���{i�9T�\�,x{!���ih�M�����ob����c����r-�$�����8(��� ��y��IX�|5�tIWS�	U�2��h�tZ�_���e�Г���!�V Ƣ���\����:��k���m�!>YrQ��6~���qVB�C�`�N��w�zok���/@�Od�K�XL.,%(���dVE�c���2o�g5�\�r�w���R�ɟYj���S��m�86pXz��G^x��QG>�0�I`x����Sd��{�=�B9��ltr����c��k2V�}��[�?�>�r	<F���ZQ�Id�C� ��������=�gnD����sې�����b���Rbg�;j@QӉ]K��	���^��l���u��׵!�+jgf�5�X5���ݩU�����;;VM��+�?N�=��7�T�pK�`z6nމ��z���@���HX�D)I��w>��L�_uf7���jxZj�����g��C�~���a
�<|fª���c�5��W��l�d07?��(XP�^�'�+DX
xO�Q�۫^QQdG~!&Fjš|��b��'H�ñ=��ĉ��)�*|�	@S��$|�Ku�����)'�7
2����OZ*ia��u��ԥ��@J`�c|�"I{@�Fj��_vB� >�{�!N�Y�� ��v��dL�R,�Ů&��@��H��9H�'�F%���{�V�"�����9��%�E�-�^��As��8��\$H�hZy�B����m7���s�4�M���ց�)�)SXm���4#�;`#9�-���	��Q�on��,�貀�����8^�[����q/���>��B���#���9p"��a{��sKD��������+�(*1������D\��Ȕ\�Q�2�	@v����s���m��Kn���B˅��޾�1+;*�;�����V��z2o�����6����3�XC�h.w8n��:&l�o���D�R�bh���b�^���8�L�?�^%�kt�ҳ��q��WD;,<�{*�uYWj�;T�\�B��E��+g�Tdr׌y�4�W<K^�d�r^�g:���v�h�����I��6�Ҋ�J�D>��Z ��(��.��el���n����������E-��K9�n.���`�a�K�Iݲ÷��>u��a�3��I���%9�|���\�Ó�)&d3bA��)�p��W�I����ґFo�%���vA�����#~�J{�fF�s"<��%#hH���0i���jo�p	�57_��M�|��ɐ��.L0w�꤭�;�"s�i�-�.�܌�����ͬ�RF�����
Y]����X����3�(A@k�	�T~�e�´گFΤ=_������D�;FG��^��H�|ڳ��SZUm7�5!US�y�|���em�0��41�Y�=�J$z�mǢ%"ղ_棥�.u�u=��������)Y��f����([Q{��4���`�F�K-���"��@��I���e"6���G̦=�jS��zE��w� r��IE�8����蔍:��ٻ �mt4�BE2�w͖bm�i�Q�I��	�|m�bؚ&�.z^�����h��g=�)HV�8���uU����ۊ���t�4=<o�.5��ptq���~�Fe
i�a������|�u�q�Cg2����s�È�2}��R6Z"�Mj)}n �f�7c�D�~�4�p��E���¸�� F����7�t�i�)t1:�k���%�Ea��$�p�;�:�lփ��gz�Rq��؂�0�,q*��W�/Tɂ��&d�'A��x?M�$�}�[��J0��cB����\l�=OS	/��Q��pĄk�E累��ι��W$� �I�t'}�z�;S��b�����5��P�͑��v�H�����Sa!tC#W3zTo�ߔ�xu��#���e�f��� ��f�0�i.�O�9'�:�y:��Ry(nq��Ǆi�	�5�9Q�0Ԇ��z�j> [+�qL�6V��������հוP�/g�ʪ����7�Tw���D.�C��-c��*��M]0Ak3V)j}��Dڐ
GC�vo�b-�6�&�����_Iv�X��˷C���\��M��/J2��qw*�����tuᷓrɫ�|�܋wFE�u{_k�����Gr�c��۝*j�$�ڪ<��Z��~�]���̶/�Al#� z֕�?ӂ:}l!$�h���ti��, 5ܩ���L�ϙ�O;�uo�X��d��`=z�D_��శ;[�$���d�δ��jD*C
���E�g pu3n�	( B#�N�QJ�Z�m�����{�7��m<H
̒D�(i,hV�C,�o���;�5����|S%��܃?NR��@��_/�2�(7����YP
f�W5�C��Ds����][-�9�񱝄�8	��"����PCb�a(���& e�C9*�cH���y"eN�z)��Wt�h�7#�F�bIv�$K��Wd�XQ��������d���Z,��*m�Ą�I&7�P=@���8�ZF��/j��̒����PhW�������4hU���"7B�
j�ʍ���`�d���Н�	`�ؼZ� Y�O����Q���OAlT���4��߬��5 �� �d ��8
[1�p�׍�E�sR��l}�uR�I�&R%c��57�������y���[�']Q4�	���
P�HEPt��9��}�A���C�9�����p)$���҄��q4�k>�*	�t�9�i޳6������r���Sl�S���ڥ����>=���x��'k�]����`c���lf�߹i�u|���=(
��������t!G�Z�JF�в�T\f&׋OZND7pG>Q��xI�S,��Q�4��q�6v�-w��CBx��f�T��D����	 v���x��Y��ү#}#��l�Y�h�D:�= ��_2�U�k�|p�V��5�t���m�W�����=��Nm�k�l,�9�#����A��BP������C|S3̎$m!��m��=���z����H�K\1��뎙"��4� �IjOx����b�ΡI<���v�r��H>jw���ʻ!��������C�v�J���;�ޅ\*�������J=>����-��BP��OД������\\֫������8����(��|����%����+;+��$Q(!���hS�gk���1,�ͬQ��Q�3�wW|��s+��"J�$d)����7�0���Fhik��zM����p�}N�	z)]wG\�JU�O��y��}�-�����
��0�y��h��Y��L'\Tt�1���5�s���з���b�N@cPؖ�y��-���]I�Ǆ��`Jw/�f8o�A�����6gI�O���j�1�"0d�M��QĞrL1�g�$�,G�X�X@�I�5���7�@��z�?�� g�1c�A��n��[��]�ӈ4ub���m��[�,!�dN8~��D:�ѷ��5�+3��P:.
�2ܡ�&�@XO�O�lP�(��Z�^������ھ0�q�Ğ /�A���{�%'�닜�;F�0[-;�#�g(z�T<�jذ���U]�A�Q5]��� �h�������1Hc`�����v����ɶ�Ӆ�@�Uy;��pM[����5����