��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|8���e5�I��d8<���ۿfk��B�8G�&�υ�V�>�]9�c��a/�
�b��r����(ڤ�$m�3�D�+�.�������9wa��"��0�+v��Zq�������V�4n?>��/Eܦ]�)h`��)���qB���-���MV��#�:����ǜ��1EC�y�Χ��Y�w鱉)4���Xǲr�-"��=Ⓩ��Q��&�0U��_�Ϣ߽�2\�!n_�� �I�I�ͪ��O�2徯��F'=�
ڿ��y��9�}��ѴAI�\(qx���C@~��4[��R��Ŗ=�R���iF
����D�Ff|�v�TY9��~�>1�ߢ.�f�{�8|�3"�j�: ��"�r��.��AC�S�#ͅ���.�w��]���F��(�Vcs�)W�B�����N�TБ���T*��TI����=L݂�bB|C�s*�Oޠ��d7t�����1oݼ,t/3��D�s�7��ߵ���ˬ�#�^��G
p�t>4ar���^U� zDL�X�?�*,�=�����{�0�l|���������qq?��+�-!h�um*���9�*jq���R\�ց��e�ҽ�d)��D�^q�b?���d^P^�2��:�/�ьɉ�,w��a�%|$�!慊	��"����:̊AM���l�F�73O�M2���sQ���+X���W|�X#�q��g;9^*��7C��"�3��@�ԯ�{4�N_��]�G��ӈ) �L;1�YLܱɡ�-�>�Qʬ�芎?,���..f�b�U�ʻq�)�	�;
�s��L-SPy䧍!`��K�^t�P�[���)<�"(����^H�u���̴�z��&A�>
�΀ȇ H�뺢@�;"(�S@c��:9�4�c�R<\�����_=�����g��@�rȀ��9��X~���5:��^���.�g�2<���g%cKi0Sb�&5!L)_�t��f���������^�67�n-����C��t���h]��!6g���-�j]��o����	��DMU��6M� ��bkSX+��0G�$.-Vh�y;C���
�ET������#
���ο2f�>��Ys+o�D�Z���бnaęW��,�MJ7<������F)!8���Vc�|���pY��Y��9�^�?Y���|N��ִ��u�j�G��
�X4��T4�'�+U:�Vg�����]�Q�={{6<����(dXz���K}l�'Iz���t�d� �̼t����c<V���A�ۧS>�I�u��]$bݕP5W�W�o�Q!�a�u[����;�s�n��^�
���y�J�Մ�q�$
�3��3C�s��E��H0�s�Q-��`*��c�=ey��eg���*�ǯ��X�#޹�bc�����t��0��j��bd���~���%��sSs�{�W��3���}�b �1^�����G]ט�v�k
���7S�#�K��{������g��9�����wn�_f��g�,��ll�d���t�峬k�hד~�^&����`�ε�l���%u�Ɛ����nA�%@�M�'Z±�>�����G@���:f�ApB�.�Y�2we��
;��l��0���nMS0F�^u%���<yL�������J�QN�*ܷ����"����y���ĔdU}gyH����5�ydb�#6GQ"T/����
���#�qat�C_Շ�w�(�c�2����Չ��tk[&�L�۝w�-�å�N�+g�L���|�����s9��F/���3�m犺�i�.}�d@�]�X��aO��m�B%O�����dy����MRd2!c�P��X_��:��ʹ4s
i�!ICf sL�l��]�����W ��P�6��!7v��$�іe�	X/u#�D��ӎ�q̴ۂ���Cγ�F��UF�5��d١�j��Z���j3�UX�#Q@� �����pݾ�O$L[�u�If�ù燫�$���o�P�O��[P�wr���O��ck���i�T�g#rYŀd�Z��l�5R������-�}{ՎR�iV�}Zݭ555$�0�cN��L��T��>�!����~9�>����ݿ��t��(�mzET�C���WW(�ۋ�_�T���F�?�}�9�>z�����&��4h\ �9ׄ����_��;�c�[ƴ[<<;��l(���'�H����)F;h9�J�<99kw���A]�ھ�7_�{��T]�n�|G���������ة�es�J&��s����,�����}�����v�X����f擆�qs>(y�ν$�����X�'d+�@�Wj�y<�O��+Ԃ�O�水N�����r�[2NJ��ӬY��o=�0���Uh���ex
]��%wM�����|����=� p�O�pl�����ZX��e�:ϚMT~�,J���<c4.�^��R�>���\���B���Gߔ���]�Zʞ����Q`#�&�H���Rw� d>okX�W�H�+p��[��첽��+����A�w��"(=2��D�����NRF��H^
^���Zr�����)�t×���� �����Px���/�\�Db���5J�8��s�miqA���x�%��	''|�
�$����'�ᨗ&w)���j�qT�"}��������/�oe��Q���m�n�/ /������|o0@=$V�?�H10�/+ouU�͞�$s`~�)���ux� �Ѡr6$α��J
Q��I��4�@l5B�	/�C	l*̂"ֺ���鼄ʣ[���܁�"��j�o+gT��[B�Ï�~�LX�R�J�:s͕�2�	8I9�ܷL ��E�֙��vl����gC�%/1�q�[I�_��5K�f��C�S���,7$��(�?<9-�/�cl�L�����V��h#��S	�Tי9P������zJr&8	�6���b�(�-��K}���:�+�ޱ?��Jy�����4��[nl�k\�L3T[I��a����{�u�\C�ޟ�{I��(\%�8S�|F9C��Z����cf�WL�宋h8-pn-��Ɇ''n�2�A���11o[�z���.L��*k�2b@�����c-�)&'�(��uڿ���:6�nv77��q�v=z>M��H�'R�[>Ǩm��f�܏� �/9�"�[�!j�Е�y|"i���6�eRhk�i��ᔼů[j��PW>f�TG����VR~�����۞�1%�c��}y�x�f/8A'�i"�w'M�۝;��� 
��$MW�wz������ML��8srVԵ�-d���(���ꛊ/S_,N񸍧u���s�Fj�i^�#�݉��!�HLZ�>M�&�
a��0�2�T�>j�zz7�R�OYO*��7"�㽻�O���ƪ%Fh��p�"�=v�Q�.�?�hkJP�r�a"��)%�΍��)J��w��R��Z5���90Hh	�n�8x3嬰�x���Y����n�܄�旓-'��;r$�#
������e��"SZ���l4 �F.���G^�����
��j�P���iƆ	��=�}c��m�S�%���&$��b}�0�C��6�V��&CX��71��hIA���ټ8�{.fF�D6T��5�R~�[������1g�:�|�҈��;s�w"w�O!O!Vﴱ@�w�Q��;���֍8�c&��X�=a"��T��d�I����	iL��4��4V��_?ΎB:jt��Ke¡�����]�٦a�f���C�8y�����"b1Dyh952y��k��/#�4Q����rlRs/5ɾs�e&��>a����s$�-�^����B��3��s��p���S?bY���sYn#��1y�5�uB�cO�z!���&lf�}�2�q��f�=�SY����|\d�䐆��		8Y��u���J�R�V�y]��ٯ��%�%��NO�Y]�+5ڹ��!*I͓chB�p��`L^��h�vҭ�I�)�~%�S�9�?%h��I<vZ�Y�^�u�y���	;�����	�?t+�����&�����I�P�H2�P�s�|6P
���!�s�[�H�AϦFV�,��p�Ԯ>�.�t��r�C��`ILZ&V�����QzpEV���g��o���{�M���+Xؿ���'@L=���f��"͕�~&��ހљ�T��;Ʒ�y��A�*�qF:5��k�	I���Lf�� ��.��ՙ�qIux�̀�Ƚ��-�,�.y .Xظ�/�A#I���@�d����놱�`�OQ��(s9�	'��P������Z]�<����SYE��tt�-�_�-�}�Ό�(��	�F��B�kM_�~�X���0͡Κ���Y7\߅���ܮ��Db;�$��s� ��n0��eA���N�7r�$�1[��<P]��a)H�m�
Exz���J40Ꝯ�ŝ�{v�3�Ks�$))�Mj�0u����Mr�� f��N-�Y�[#|�v�n6[ۻ4��ֽ��D�v��d� Y4*e��[�s�T��U4�t@,����MNjm
  �p��f���z?�ࠎS�;� ���.Ϯ�U�>���l�N�,�6M���M�[�ڳؠܼ���9��mS�ϯ�%������TFNM&�@4銑�eM�-�;�[��Z�l'�+�842������p�@5$Βp�%
l7�9>��͆hV�5A�'�6���y�(��N�>d��|��(6��8;	��a��4ݶ��Uo�.\���s"v�'�>�2#C�b��j�u��@�"�?���ǷPE�Frk������n �p#�=N����~1�ԎV��y�l �r�㨒*����Z�� ���^@���Ufς]t[���s�+��"����!)�]{���H���^!q�²\Y�K��?q:�� 1�*٠U����" �Ů�em�uL}�;
S����me����lt	Q���>��� v�g�έb�-�� 3U�t+vre�)�z�*f�&4U���q3bg�|IWN�m'��JmE���	��@C��(����~��!�|�ke7�`O�_ՙ�}&��LYSOBꎘ�=(��[�G)s�~M"ui��o�3Q��rQǚ�Q�9�K'0k�u5ݟqG�'7�pc!�)m5�(�mpO��A؁t��)0��i q����zd�jf��(*.���`c��6��G���ΰ����~�t%^�
$�����h5]z�n��hBC��S�vg/�a i�R���HuޅP��8�P�����op�A��Z�9lJ;
�ȁ��<�&Y�ߥ�Ṿ
V�%eHx�h�_�u�m��+��q�%ϲ3#GG�אg#��1�G��'�%\�߄l�~��k0ɋ�_-͛���'�!IK��葌���9]���dǵc�Y��,"h1G�0.e����-Lu0$xr|mK2Gܓ	qߟ��\���A�s�ƶU�������o���E�,(�,~\���0*�������G��k&�\vqh�'�a�ZCK�Ñ��Y��ڡ��TF���R�p�?�P��?��>4���Lk�6�[zra�h�S��P�ܿԁ�T�PN-�3�zv�8*:��/�ٖ3�R��k�v�HV��&W&�Y:�g�8>�v�Z����	?����՛�|O!d�s�6�{��n�*v��M�XDb�KC�4.Ťs#��3q	h��zf�-�ae�t��rty��y��j�xO2��Fa��s��������M�6o����4���r@o�h��#-�+���!�P0�ɻ�;(�Aj��g�e�d9�WjS����	�P^�R�b��m���0�֎�^F@��E�Cg�Mێ�F����z�ղ�Sp�q� `1M|�x<���n�y���$(?��gR�!Ft5�Z�#v�i��Y�#EC�1�V9��#�N5��=S�Ş)6	����Z�ޗ��$��5�X��ܭ�u����&�Taa�'�Nko$y̱����5V�����>�<�q��?�OM�o����mʏ��r�|J�����8���~�*�׾Z��~/�O�[Y�z��W�A>�����[ٍP�awB����D�S�-ޢ�p�|��w{�u ld7�wj�e��z� YN�b�I��I��6�
T��S�Z�{�X��������_�7A]������	�4I�^C��T��rO���5�\���P�ǫ��/���S����luL�����0
�j��Aއ�i��D�r�J?��vӪ�f���Ŝv�Yɞ?,ˁ!*�|��`���<[�?Z1�4��<Я`��W�~v�n����DO֙��:�nV��\�Բ�ʕn�)��-����݌>罁�~����γ��e�22��f������fi g]%�X4����}Z�<T��ɥ8�E-����{����x�m��9�<�#b�F����^���m8�l����8���o�0V���;o��
�/�Ũvŕ^ʅ\���[<�nDO80̓��"����^l7/�w��\����O�+�𯔙m��X�Y�5Q�Y��3�Hw�6���O�c�k�G���W��'|����# K_�1\!�,`�9�7���<�l�(j0��Ϯ�ҳ�wh�4�dϵ���65�~]��*�����T ���g�L{ṵ�}�_�s�h*��?�<82��( w��j+��x>��kq�.7j9���JƷ�Wk=[�w�@�����*{��_��ϫ�裩��%�ˤ�ܣ�8��ݣn_�m���3�I�O6�B���mos��^A�o�@M�?��m����	���(�� (��ia�!֯�����Y#!��B^np��T���L��2Nl�0�{I�ߦ�;{n�JƖ������1V�J��	­��[����Sy�{>���i_#a����~�#�A�x�d:��ۆꖊA 7bd�h)2-��<��fW�j�"��_F�B/�E���Ih�oas�7u��kA����K���V�T :.+ Y�g��Z���K��F�Ca.e�\c��[�q��7��f��	���ݣ�V�2v�AB��ϱ����/V�X��2�wÌ��羒��������\=��k�	q,�E4=����BR��y|�Y%� 9$��Z���Vޮw歫�W8)�i��W���A���\r#:7p��NT�c�!��m�W	᝛�$����$U}~��{��s%��A�9�Cr���+�Ώ���z��u_�N��b�_�y��7; �|i;,tpa�q��f��z��p�fM+��>%sFѬrh�T�pNʉ������/��udZ|�2�#ԯ��<8$s�"��GR�� Q����3L���a��9!!Լ��D���G	4X��H3'_���?C�Iv��ݭ���@|j�J�b��$aQ�6�,MȬ��АStwǉ�S�pp,n~V�9�x)H0g�^(���tQ1�w�t�hȪc��6=��(~����GĊ����K�\��S'u�����������H'd�N�wYyҌ��U/��Ƈ�8~����;�ؤ�Q�`�g9�|�g=^3(��+`�&$�V���d�cP6�Kg��-��J�d���y�$�͚#��{
�.o)Jd�N���?8�����p��}Y�I�Rl��)gH���ƚ��B�]��n�|R��6�<�����$b>E��Û��~���"O�'%XQ9��4y�D��B��is��XUfz�O�u��ʞ����cM���I6�êl�x�;mb�uu(&݈#��-f�M�"%�S��N]ThF;��b�{����`m��G��I��>�>�[��W]� IAt�T����*;�}�(��@.���� ���ןtZ;��s�B�T��{�o��U�������"d�=��5`L�� ��)���ouTe�¢28��Q��\~/�r�gyK���46�OwT���:E��������du��ڕ��>wW��X�%�S��>��E�"H������s뭝yf|�*���G���q�[�u�>!f���+�jG���;�u�5a�5�T�i�M��M����J�/�o��S���sX��佶��OP�	j�1�����v�D�� ;9�nK�U�����#�!H~v48S��(G�.*}1������4*��x�H0GmP�̃�d���?�#E��j,2a���/e63m�x�� ����G���OV�����&��ѻ�s2�L��R�!`:� OJ��S�0ю��*�p�qJ�w�~��b���~�Kɑ,ml3�4�2�MS�w:T� ?�e������49�+)�QC����=o�����`z�u *�������&Yӗb\�+	��h��'P,����N�7n9���,20.� -����Y|�1��Pe�����aX�aM(V�e�8�x>�!�3m� ��-�?�ԬK�G�K/�>:d��<����U~�`�0��P�o&zV�v�t҅F��t��ׅ8ʏ
�z��-~��aF'p����w�ί>ĝ8�a��Ɔ-��gd��=I�S^��2�A����]l�ږr����4�+JbE��?��A2(��yشW`H�G�rh[�U-����8>�Q)��5�E�9L�U�S=\��x��Z�N��;�%}WTP���e�@�*U=��LjA��
����j�t;5/�`�E4�1�x�e��﫦�����4�9qK���u�Ww���lc��k��5���O<c�BFb������"g8�q˔��{Ņ
��CB�.jV�H��Ht理��V4>��P�C�N������b�Mw�V�b�#��n������j�Ȥ ���ʓ�x��^z?8HV#�z�Ȓ���Y��F%S;�mPm�C���"V���{�w����M;٦�^�C髛3#y���E����o��\O26������S��y�ΚR���ñ�l>2@yڛ�
4�I��B]���y�@z�,�ڤ8�4}9z`��R�Ȫ��O�&���p��4*���J"�
���	)� �W�����`�)9SaQ�/��8:ST\�?7��p�8$�%�L&��	���l����鳵?�8��.r�Ac�Iֲ!�Ĳ������圎�5���̦ԯr7�����䯳 �(�aL����ZK���C���O+�/6�*1�@��v澼^k���3�$��eOkJ�.L��Ô��f�����-���B��֞r.)����>֓��̣XN;8�C������X�J@�yv����s�9e�h����2#��y�J�F����� U>#V>�������p�����W��]�T�Z5�0�� �1{KShg��9�(��CB`I�-�̦�#��m?ߣ<v�U�|�Y��0*d�8�.YtB�I�� Oiw2b��nz�d�/	J���r�C���e��3bdM���H���n�����d��5ntJ�7�:��7��Vv�gS�Iw�#��@?�Ul�[g���ۿ��k���#������jp���iqO��S.)�A-�J�e-��[ܺ���TO!*���)��DJ��A0х}VC��Ba`<t[�������
P�\]7�q8�,�v�n�&0^�[0��p��zT/��Ύ�#���g-�^�=�6o\����MSD��'���x��\����ؼn�qv�^f�=����xd�>�8r� N*�J����;�7��7��ȓhN��+�$���M�.�:����"��������Ω?�}��'Uo7ń3��S��&q^&)�د~ܹW��V��S��|�q�הwz�qp�J�2!�>t�G�'G,�}h�C�P�44L�G����}�ѻ �eF�&�.�T��A����9lS�����\��G2�6��O�߯t��)kK�Cc�| ��U���#��3����Q;I9^�����r$�i5=�`���}x�+Ц��|uH@Y^�w��\^�k�,�����"�C=��=5�6$����7\P���Wa���f	�Q�Ѽ��l��o �Sx+���*6��9["٤L�7;ڞK�7;�����|�_r�#�v-�~���+w����'�&$	����S�_�.�E������/��0�@��[�@QG}�u�a�ԭTDQ�&�/1c%YrE�G��`��_�(����0��֟�܅�������ױM�zD9����[1	lsw�5dS��D�w�/�BM�D9��	t�]����xS���As��F���W�5LP��_�RܢK�w{�l���K��X���<30c��^�:��Z��dt\���u�)$�6f��o51�+h���f3+E�V]��ݯ�Fḗ,*GZ�JM�������j:���
0�avWpǑ�=�b*�e)v��+ڋU}l�nU�D������MG1�h�܂��'\H�MH��n �W0������p��华h����Q�U��Ж1l�4��#�⿅	��~�G�B���A�`oi,��G��o�E�2�t7�J�}\:�UX����4:��f���2xc�A&N����I=2)�qe��	P�����C�����8C�	vC2��ؐȔL��[4,�K��~�Bʸ#ǎ/�c�A� �f��ӭk����.�ˢC!��)�J�@����Pn �����ׅ�[����wO�Th�#���sR���A�S�)|�<e��c���&>�?(A>�J%Ѕ�=z��Xt;�����}$ �if��u��q�d4�yѢ<�p��S�e��z�gq�d��|}��_�������bzZ����9SB;I��AP��ܞAuŝ�=�p;:;�y�Z�}Ү��+�V�&9�h0��a2��v�Y�����Y��D��JN���Z\נIv� ��z|���c�9��F�W��>� �2t�qϟ����1��Qh�VqlZn5�cO����ѝ���}�����N�6� c�D��0U�IR�	�fz��w�>8̌ie�� ��c#���W��:�
���%�:���к�e��"�����!��Nݛ�uv�U��rO��a�Y Ӊ�F�ݖ����0-(�����@;lMe�|��{������$�)�xdr�}�EGR��U#���֘���7���bSM�G��f���KVG��������Ϳ��:�D�^J'��|�m�z�i�m�m11���#b*�"1QS�a�kD����̐(�X 	�B*��D}K��A�]�R�9O�'�w��КLK��>p?���P��Z�6ǡ��;h�Ma�{b��xEfօ$}o���Q
��i�/�tG�*؃!��w�Z��u�3��(��fzWi�7��m�6�O��4�� dŔ���*2���e~��Aeor�����<S���@�j&�8<٤��[Y�LAǥ�+Q�l���Gϕ4�M�	8Q1z{[\#8��)�����u�/��ji�y#�Xb�%X8<0q�{<H�햡h�m�^�?m�+)�O�R�xU�*�Ӛ�0;6����������#Ct��`7�����V��?��D.�;���Y<`B���uFW�z��@-BJkj��\ۗ�j����
ͨ���DT�ʗ}n>u����b��>4����ƙ%��N��������Y��F�R�F��O*�Z5�j� %�I�v�3yzDT�����+#J�L7\U��X�'(�*�T4����7�A[z.�rV��L��M<�e}3���E�C	$ �	*��iA&��YE�R�2j�*Pb�Ah��r3q\�s/"s<�������Fh �� /)�h��CALP�$E/�jg1���o����	�����_�	�|��=��� I8W���L��F��&l�qΞ#g����m�DG��p��!���D��;�)�=����~�d��|D��E	�Jmo��KE��}�TA�N�ei��",����y�x�'�)-	GREL�en
%�/�Lpy���O6�g���p��bT�3��"��Ɂ��`����ר*���n�³�,�߾�|5�ޕ�q"_�d�	@N�.����7Dg�F9��YA�M�O���� e���T�r���hp%��&�a%pX���O�*��ݺ���0("軠|Q����*�S��]�c��#`M^i���j<�L�ΑPӶ�m�$�V��Z�Yu8#$���1D2����i�.��ǅ��v����k��:N�N��;�y�b���7,�4#O�7�K�v��?������������_d ��B�����C�S:}8���J����ڔc�ⓦB��y�R�?�����C���'T$�=�,�e`k�l��f�ċ;��	�n|	+�B���@R,��KX�����?{�0\�jT���lD,@�)�e��
˭G�=B&!�n>�>�)ab�-�I�f���m���Q�g�.�!њ�]��Δ���>e	Z��qC�Vr
f1��/�qR��@��։?��nn�%@�h(��a#e���9Z���Xͺ6=+x���Sm,.�wr�����z�<@N8����z?bXuX�X�bync^	Zp�c@l���n��3�Y5u�ԫX�s���	�4M1ɖ}��bb����/ B~lQ��!9�!։�	o�������Gڰ=���B1�Նy] �v�L�vo�ƥ&3u0L@jq��_�Y9��Y$�{#/d��N
�2f�fL�N�5��Ksfb�D��;�wqj�f<�#<<�����s��D�ԭ2�����]۩!W��=o"�	�c�LA�_E�Ըx���F��[�Qh�%z�9M�uHv�ݍ� �#41�_�6�C����
��`���"���S��I}�D �L@�vӟ�8��ޣb"˅x�,��*WS��J]�!tB;
O-�mf�j�יŎW�@e����eW����K3"f �9����(*+ꎥ���<�D;}��!��"���r`�B5�|�>�#|Sv3>/��V\RςR+��<�n�z`���UրY�X_D�v�o���OPr§����YC���YRY�J|�qJ �jv�g��Q���I_��Œ�BO�VC<�K5�B1��I���v'�L<Ґ{�viSԮ��6�n�4ݟ����6ǀJ	�10��a$Sf�@�9)��:��Y�����A�R��G�io�=����~^��$����	Y �즪���h+��̩�6F[r�;U�S�H_�3q_��$�ޥ�΁�B���SY�2�~��rK-15����ԸY
���[�rnG��=���v<􉐢Lk�վ*����7|ݠ�N���	H۽�sw�E�LRB��q,K:V�����N7��˒�0u�~�v�޹Z���v��r:<?�w<�	�E
t_������o"-�_`H8���4��V6�t����6���*�!�-]I�'����0��`�r�����4ͷȦ�v�jW���Ѕ[?J�9�X�V�^vhZa��d��"\aG��#���Ϟ[;9}RG��Uypj�Z��^�
g1�]�nR':�b"��iL��WϙQ���a�����r����Y}���2D��n�bC�,h28v�G����D�����͒ɐY�=�Ҡ�����P��8'�/�C-M����S�#)�5�atnl��wH�|����҃�Au"O�u�����ޔ�n�5pF��E�֏���w�y���.���x��Ts�П��9�0����V���<[�H��[��oe;��z���:��v����"vJ���8�Ue���q�J�>늟�2C�/J�Z?��
��v��P��m�v;$۽X�b�¬�̓8����g&�:��̛&��	{kX%��]�ڑ$sj`���ҍU-�Z�Ǹ��ц���P0F�P�ǯ �C���TR��K���B�#��0��.}��c8[�/rgk���5l�ޜ���Q��MDo`�;���U0{�(��]d�0���P�j��w�v��h����;}Ns�ˣNkzR���R�[D>zr���d	v���7[ ���#����Or�6���Ѩ�����>���tD�,��s'�D�V(�z�=�D]DK�u�]gDp�/j��T�q�O�T5��j��{���Y.�ؐp`�l��E�n+o����M�l\����s�_sf(bB]3?�(W�^��͸��^7�0��.GÑ�o�W�Qf��z�M6���TG7ڝ�l�����7�������.P�h���:�T���Y�m�����(��{5���b4R��Y�I]�(��z����v���t�ƅBA�1~�G�W[��w(�R	[�$���TEKtނ)���!�G�k�9�8���oF��׃��(ޟ�^����q*`�,�����g\��K$)_�dUuk'�e��ܚu�Ya	<z���(r�&��|����
0�YH��`R���db��ۙ_��9�
���г�F�bv�J�bS���0G���L�V>z�����{��%��p�#�[�j�,�L�)��{?��1د$��Ȯ~�E�?�<	��-d!}����(��6�d��
���U@�v��f �D�Ƒ�;n!�#����7�bz�W��[�r+���
��Y��3��v5�p�On,(Cړy)��bQy}',�3�T�AA�PT�`���P���^zD��5+ſ�:��w% ټ܊��-ػ10^&˓�J̨��W<�ZҎ��/#�mB-`��67>]�z��9Ә2n=$l���d6�5�M}
qI^���V�x��D�!Ĕ�"EBR2�W7��1�$ٲ�����w�2p��;��;[�l�n�3<��M7xH�C��{l��f������`B����)��ɾ�4�;u{�_Ʀ��^ةe��_G�X����}�!_���hXK��A'�BIbE�J;���@9��X(6CX/Z�t��A�Bѽ�֎��	��i������������t��_/�&x�M!�`��N�Zҟa��*�T��8�y�s����`�F�2U\q-g��D�R*��=_�Υ bt�I�6�PI��@Q�.��uY��[?��N?N���Y5��艻D.��
�mc�ڈ�>ӏ��8��Ku�ŹB� >��?�I��o������Cl)Bi��7X��4l��U(}�d>]$��8T�G�BҔ�[v�Rv��_���X�y�WXR���PV̕B�_���J�X�c�x:l�-c~_r�
+H$7��~�-�&�P"��>�m�jm�+�`�\��!w�N�{��s�gb#�]�\�fjiͬ�F�|��a�i��B!<�ҬOu�V�;9<~W��	��P$�g���Y���I�n��Ԭ�jD��P��y�+�����$Vhg������1K��t)o��[��J�w.�����6������]4ԫ� ,GX��Er�i&�q(�-��f~�F�a��T��gK�i���$%K�1Q3҈� ?�����5C̦���������(�D���`����8���s��l��V���$����Ϸ�^K�28�����/D�������#�:���P��$_~խѾt��*�^!h�k¥�8>�ֳ>y0���^CW��/��9����H��=R����ݛ#I�>ې(�Y=���aW4�4Ƣc�F+�?��{&��h㎒�Ԋ7&�� 
��eU������?�%�
�Ľ�L�H��aa��-��1˺���A�	�#���/[x��V,�n>'��LR�Ձ�i�
�ή�ѧ��?9dO���&��ddƉX����[-<�w�}`F ����i��:���K�ց#�y��5���D�+����|�霌����Ci`-~t���n�#hh;��/�ůiy� b��l$;B7f�L���m��~j����<�6o����3�6p��}�T-�{2�j��0e
�x�n����/�ro��21!\���[�* x �-��X��}�B~$� ���.�?A�Wi�xqSCfd�DY�p^��f������J9uZ_|H���<��9X{���~Wd �RX��[Dx�}LP~�����X;�mi�c&t9>�x E�V���ђa8k���,S�р���
���17������/	�=˃G�	����B���m��O'*���Y�}XrMB�"�g�6�WY}�-��g�8�e�  ��ܺ�Q��n�4�c��޶���c�ie[xZp/⽫M��a4u���H�Z�tb���랴��vs-���jm�@/9�V{f0�f�M�l������E��|ɒ��-��]�q�7�R�{�h�F���$�6��0y��\�ջe�G��Ǒ_pTj����R��q@�)��NWe4-d@�Ӽ�'vp��a���?�I��QFLwX5���Л���[*
��W�!C�y�q�L��i�w n*X�Hp�Sf�*
{}P��Fj�����>�$􋟄�NWc���D��)�u&�J۰��@�Q�����Ϲ�.r#������s��-�R+�u���d�&��� ��x�ْ��Ci���o\nR2�,����v#�>�W��`�ٝzQ�!�(;���+LZ�ݑ��S���`�Dȣ��]����|�#9{*�,pI���trN,d�e�2����v �4�	5>���	Ȕ߲�^��Pv�ۖ���G�w<�㗬�(����bo��6}��^����nw)�38N�˴Ir���~@	^���Ev]`��5�L�þB|eQJFqv���L��V\W��d��v+� T�w��PTJ[�O�H�J�[�˗���&��6���c�'*�LO@5uڛ����"�wWSM�o8�7�������ãA��0��o�tF�����v���=��e7�P��K0����U �Ki9���d�@�Y�E8fѣ� ����5%�v/W�=qYD1�����;�<��Llf_W?k\S��v;�3�]�Q���F�M㑷&G���#�>�)��T�dBǾٱ2s���4n1��l�M?/�1�˚2��賵�������-#��-�xAEi�nF0�R��}�O!�3� �>��-�c:���>]�d1�H�a��PwG����X$�dh�&� �w�����b������eT�\������i4���?]�yR�t
@�MO�7�֩~��n�9a��,��>��\���CFKEʔ�А?^�0�ݲ�d�inѺZQi�b���Xdw�'���/����Fk~q�靖�?Ds.��L*(��|����FGÞP�Zl��r�|ނ/!�W������H��@}�`n�{_*�g��2(�����`v���eM�$�1��Y wC�Y�2E���X�&��-��t�y,�B�^O �EC`Ӷ� �F{y��si_�Hs�qO%�>�g��Z%��&�5�8o�;�k@�q�y�ȥ[-������E\l������y�j��Zwg���r������������%oǓ�2wm��%9��GC�{�f����D�tc��2��>���d�C�m~���q%��Bo�fy�
"�(z��b��4����8��s��x��,_E�)��J��`�ga%�yeF�8Y �z�me6�����޷(�l��L*yeR�fO<Q����5H;�ܳ]u�d����BH1�3{>M�)t�&?�`��4� /�
�\0���,_<(k�
��8�dm��<�cS������Uo��M�!�hG���;�2sZّ4eR5���p侮�TnĮ�W�6���c���>a6W�ԓa�U69�R�~�����ݼ3.�S�WaEm�f����Ob�pU�<O��(���4���1C�zF�R��!c%�ܵi����O�k*�*[W���"��z,�Ø�^>S咙z��r���M�V%�	;e�y�K�h(����tG�k�-���pk���c��B��+D��ձ*v�0h�=������͖��|�<����>��rFe�8�k8T� &�n���/y�yf�J9�-!զ�lޓZ��m�3��ť(F]h/�����<�v���j-R�I�u'1�?ˉmp�t����l�zXS���[ʵt,j�W��2d��
� U�պ��b碮��\?b����RW��b�?;��$.Q���]�O���7���,�$����/q |>/���ߧW�����+P�:G5��'{Ê�b�MX�=*��_$�N7
С"�sEk��l5A2��a^�!����ki��PnM]�.��҂�M��8a?��~�Ź�g[�q��A5��& �-!�n�{�G7�cyF���Eh���r��'���g�05��#��T�b䍃�T�-�|<�+v�����o:-�i�xC���W1�V��N��Ҫ�YmO�s���
����)��Q�<Q������_��=�<jO*t��xɕ�y�!��:n�n8܂��,�Oh�A&�@��$��r��'zm����>�߆%��T
��[_��y�Ϯ�~eZ\ޖ"�lU �������>ՓL�腖l���A�Ф���8,��k����ai1ѿ$��8������
�g��9Y�|��f����[.��?��v/n���M�7�EW���Y@�_6��ʈ�+P ����OW�,l8�Pf�)�&�l���tf+� c��CK��Df��D!"��������4���֘�#�'�,�?�P����^��r�
�_ј�ܜ��(���V�@�o��x�H�g 
����5��C���� T�q�35�q&�Tq1����8(j�}"�$Z�hE�̆��8�'?U0k&GQFV�J�z���:l����Y��*Ńw`:q!b����p���9�RPЬ�$:I�6|���l����m�Z����3��?���=������zsE,t�<���\eOAg�P��W$c�5��eSr��QeU1���w����$yY��� ��)��p4�AI�1��j�ǚ���=��ƪ	bq�<����(�U+�\$�	�&GNF�m�����ݷV~�DY�eÑ��} ��D���}��m�2�ċ�jH�|FJ;�鎰���F7b�kH%%D_{��~�{Ԇ�& $��a:7�Z}|�r��M��4��Gᐇ@���n�Aw����s12ŷ�x'�ɟ�Dwh<k���������Y��˷t��ࡦE3��M_��xu�pT4`��@}\PvU?�pi�0�j� �����>��g�}ȎR��vY��QA�<B��td��ru0�u��BӔа�7Ē"A�������@6�i���%�������|#oϞ~��C����SՈ#8E���Z�ۜ�&+�Ҫ��k���4��38����{�k	�r��Z^�`uAq�~6�o�,�>���V���ϛG7tqwCdv�T(��j�}P�~2F/I),�����ŀ@o�ks-��L\���8�s�Xwx.���P�΍�w�p����aC�#w���e�f��^1W�I��9~�A�vԇ�T��fz}d-����MuC�#��K�\OX_9��/�]����7s��sӛ�I��Ď��٤��F���X��@�k��k�&ޅ����������3m�)�P}!�)���w�mW�k�+�\4 ���c�UQ3'M��mH��g��8��7�4΋Ͳvz\�zʱ@"�j���+P�X����C�p�A�;ė�_�J���<���bS��� ��}I�8W�?��L�ֳ�mZ������43G�P����S{ž�^� v�|�#2�4R:�d�1��Ά�/�5�?<��e�)xI�G��$ϵ�E����Č���PCs�Z��[��C��\ԞP���⧏��y��"�4_!�{P�/�����Q�����c�(8��^��jt+Y�_dX�	�l��G��,�)�^�gH�8�n:?��ڇ�7(EP���t�9�	R����[g;�&�Ư��u�˖���ͽ�:�~�EL��ʸ�gB�.aV�ٝ>�v)��np��T^ )����Z�u��|�~V�Ye�%@���:���/ҙ#�	`!�(TxG�ʕ����.�Pm��!�ư����>��n�Oen`<	#�00�d�S�C��(�sz/�������^bP�c%��2�:����:8D1L�V� -$�d��F�\c�� �r�Y	)��}V�It�o�)����t���]D�x%}{�N���0�Y�_�,�G��e}��j��s"�V�
>%�x|�@�Ċ���YF�#��h��'K14@cЄXu����@�:Z�t/��v)*l���B�Z����R	�/oH}��U�V槯��%A�eZ(ŋ��L��H��u+�ؽ-��Mv8-Z��r�ڎ�n�@�9�g����r���ōi����6v��
�.���FK�� �O��e��T`�z��>�ZV����ҧ1���Zϴ6��WT,����"��&���"*M�NVe�l�㥘�J�pA*�rq:7��)O��%�dq[e�t�{yE�%C5��C���x:Av�ji��3����:��C(�5 ��?�xj����]Dj��։�I�]L{\\A���DɿV1��r��0f�i��w`�0��N�$!>�	��/~y�o�l���9�����`��{i3��qcani���2��`�v�z=��3�'�����W8�SK��=���j'���;G��8I�(^�������%��G�*iG`�8ۅ#W����uxL)1�L���UÁ�Į�#�F�!��̇�� �fI*Ls�@*�ͫLp��*�Z�	G��~��t��57�rSB�5��y��n�ć��e��ul�	KݹS�.�c/�!f{~��u';♤'�P �4�M����:�5���v��9���
�C�h�r����p�c(a@�p�|3JJ+�֬۷9B9G�|8K�UA\�G����N����w��P'�P����Q)���J�F��ʷ����L/i����q����A������l��c�FWA_B�+��I�2ˈ��3�QǶ{��a���������?�a��7]���l$@�T'Nc_'����mIG�1�i��J%�i��XM�+�n��[c�I`Wl�8��9� @mE�����0;^~��_j[0Zֹ�u��5w�k�0�wMg�2���߄�K8�?���2������T<�Y���Fgt	3��e�C�0�~m8��;᧤����"�Z���n�*�;�ZGwHA����G=B�����hô�;���,�\˓��1N� �S%{&7�
��5�ݬ�#���9���Ǉ�bJ.�9�k��j��-z	F�%(�f���"G�8��{��zf<����Ũ$�2;���.��t(��"aj�D�֗2 +"�r!:[�(Awʋ�Һ��.��lш\���	��oR�d������)h�]�L7����
�)���T�!n�(.伭U���%X	�}a|��ן��z"��X�M�[��HBmC���ϝQ���)\^
�.�}h�������Kg��p��Zr|��qpf��$�r�E4+[�j����/�dBb�+>�5[ݠ�m��o��\󷳑N��/8a��f
��ս�����v� c8�M�u�lh�������v�I�.7���}WA�]����Ф���u�/}_����\����w��>q�1KA��������+��Ϣ�'�j34�尰 .��V�yQ��Ճ0)s|S���YՐ��F�E�:@.R�zKd��SڭR����Q�`9�0�C�MkL����/*|ϑo�T���
�W'k8RJ�,�� ��Π�Z|0���/
Sg���|�*�K,���#M
ܖ��z��Ȃ#b�ۋ=3F%���vT�k�]`�����Аr� �J4�	���f1Z���2%і��$�ǣ�Pp�l]������?�01c��#��ʟZo'��:�q;���G����w>^O�>I%����c���d<n��"	��?&Y��.�#�n����#�M��p�a�o�e��\��|,m�2��ho��"���r�+��ed�2^��K�/r�i\qTHGߐ����>�d��X�˶��h�Q��V���F1����E)���8E����틇�5�Ed�"U�g�6��iC�^�~�%�*���u3hV�O!- ���|���P�i�	~f ֬,�]s�H��S�  �1aP�_��K����ZY ط��e�?J��fV�x�W�� yB��q$Q�������|�^��u$^���c�3V��>{?���r
L*AE���^�U�M"� ��jtI{"�iir�A�yp�ژ`�%�3՝��K΄kB�PD�*w�Vu����uu�h����ư�5�M��8��^�O���H^kZ/r�*������̌�Vl�E�ڶ�~��D��&4"vD����u���_���{ގ���ש�\��Nu $�ʜ��5J�7���hǄ��m��hl�^AzlCcr�BD�OW]��88+�#3(7" ��Z(n�nǮ(1<,(�e��}r�����I�VX�k7�z���?<5���`b��)���zӧ �{��6 Y�\�Z\Ɣ{ϗ���V�Ӱ������m�d9�faGjў�bM�zo�lpQ���hf��g����3?��{{&��ɑ�)����*V]���5���eKN�#í�>�p��E?#�6t�m��`{vr�!�5���)�q�b
�&X��Y��?��� ���UЪ	J�a�)!.��Ӟ��.gog�t+4�_`����svy�#�B�s��Fz��k�H����{�ߝL�Gw���Y0���0�0�r;�ҩ�\ܵM_J&�N�_�̀J�pz��$����h���%�ا�� �m�}��&ci���zA��>z������6��z}�=ӧ�z��L;9��K��j%�F��52Ni��Ap�XY�+�~�'�z*̂Jl�FK��Mu��;�L7 �n��e�n�
�`͍jK]�.�]��B"�����ʫ�6*��ijڞ��P/u;���{9���ߋ巽)��\"f���!����pa6"��2�A3 �����G@��D��T���~�)$T���(u��e�,��� C��{�,��f����x�F��ioް�`�`��ĸƹz��Ns������z� �p���&��DD�'��+D���>|<�y_���<T���?�i�elٚ:&R���$�?g���Q��6N-�����K��0k�����a[5�P��>a�(҂�'4�����߁c�b��>�2	F#h)�����|AL;���X�sevRc��8E����Y}N��h��qK[.���A,S}���������,�nR�IE��%�%"v�_��X2�������J�Ͳ��u�S��Ë�������M�<�FK��E|����D��-��g��	c�;V�$����W=����$��nr��V���{P�N�K&��-�	�5����/��:�$l{��J&n3ښ����\^��>�h8@M���͋\7�� ��&��8����w�u���`6��V��%�m�p|��%l0�ॺ���GZIg<�ӈu���y�v�R�g���D����]�$2�&M|v���t�zj	�ڝ�����xA^�!)4v���X������v~)wJ�Zz��[�=+��, �Mnihk��b�7�x�>oa����˵t���5g�!c
s�T�K.WW-�b�.��O���p����b�K1�� �et�
��ݘ�4�Q=�܇J��!���l~޸��L��d�|�Y�����R�Qh��WA�����ܺo��mKv����V�O�骲�HQ���&EF�􅱥�����@����i�76���O��%eF:���"R��i�Dtn� X�]+||�zA����}[�^?CK~r $�a|������[ӭ������kRmF(�e�1[[B���*�qUJ/�Qr,ݾ[2�j=���@N��Lo�+	*0D�W������mM��)]r��� gv��AQa��gwg�I؊��`%����Qg��9�
�#q1�i�=�*Y�2�v�?�ub�9�n@��f�㌩�4n9RO:��8���0��>g�0�`{,� �0�e�.�'[������f�����qT�N�}<	�XbZ�ּx���.�'�A_ޓ]�jcM�+$E'3�QT3��DHL_G�L�$>3��vh3VOq	�֧��hf��ZA.؊��"�.|�e� �"��3Ǐ�i��t���w�*b��(Tc��B�~�uyg���m+h�&&A��3rw�RgC��m1�C�8BSa��g���3��?Ջ�: �V*;igB��2��V?E�M~�#v�=�cQ�dDX<I\ݨn#�Z,O���˪V_�y�5<ǵ�j���XQ�gUh!��s��\�⹺���@r�
�\���&pe���b�K*=���m�'���$@ھiسq��/��`Wn�b ��.�;������7�ZB&oR�����LW���U(�m|�3q-O��Ɗ~N��~b	����T��!�!�'���ʌ��Q�)H�?�.	N�bd�p�^z"/{��ii���А�s9���%��s3�y�pz�`a�l��*W���,�T1_�-B� ֋�hX9�}X�����"\�5;�j8|�Gr�[�>�MA�KP՟�vg16��LgJ�X<�3�Ob�Y�ZU �̾&��'�z_'�c��M���1H	2��"�Y�L�A҅F;�ύ�M�ji�:� �5��_W�Gy��<������Ke�2�W	9�r�3|	�|�3|��Wz�$^�+�Z8=c�l��jآ����^��w�d�mI���)��ێ�?��E�S�j���8Ё����W����u��;r�d�O�u�,�v�ߪX�?�Ԍ G�0�F��E(�w��q��դ5��	E�ctژ�=c�0��ŭ �/�<��d�|�Hg��	�q�b{:`�,H�J�	�Pd�=�?K��-<�2>��L�5���U��������&f��z�-�$�/���'�TE�f��	���d�E�68�re&����H�+E^����6e9���0�[�pƈ1h)]T�ўWWG�:,yƹ�7�-�&�(C��:�*.��?�0�nn;�h���0���_�BQz����b^,��C8sʛ�v\E;=3�7�Ƶ3��L9����|���!M�����z�M�<�1j�#���V�K��ΜZB Sgl4�������"�
�Q���#&��,9g��3���9
��t3�&m�$��4拼?I
O�p���WZ污y��p�]%}���	�<��>ya�AF�DRrF��A�7շ��aHQ���*��"�´��nF��z��ĉ^�~�I�ղ��j1�I�x�C����2�~K��D��y��1b�����J'��IF���iE��?n�h��"Hlߵ~�>����_9����a�K��{�ӻ���Eֱ�8�Gn����5��u��*]�YC�I{�)�I2��o=��Bl_�! �� M,3@�Uu}����� �Iڢ]M�0�Z�� �e9 F�d�1���O
E��DAG ��So:_\.Jw��!�-H�֗ĭ��d�{���� ��l�/s�U鋖m�5�b��f�C�Ns�ʏ�ZH5}�zĀݺN!0���,tp�l��[R�[7�a����9����A��=�n��&<jn�qv��5��z�@:�b��sW��Pf\2*�&:v֪�pon:Wr^��&s��T��)��b��k6���<q"t}k4W���'�϶��Ws� �q�I�n��N!�=�y�X���0:u��[k�in�^*�����9P$�U�2�].P��?%���#z���B�5G�����@�kR�l�qZ{;��p��x�ք�i=�O��Ƞ\ul8���eqhip����>��a�=r f���	�m��.�<C�.�?�{Ɂ5����FL��b���W�J]�Dq�61���g�~>����)L�۸jz�b����G\L�)/���fA3�g.���vײ�:�{�r4|u�D#��*���ɞ�n�62��#.�� �F}c��K]n��E22�iҸ=�F^��Q�C������<˸])�#t�����˷]q��A��J�2m�̠҃�6#�eri�S�n�g�7�6W��$L淩��\ X�Jc��;�GW����@}�Y3qy���B����yNUD_�lNm�ES��#Ž�wȥ�_6�0��飇?���٭+����+8�	�wNzҿa>��E�Oo~��--ʅ�!oS�C����<ҏ�!5��w!hv�?zy�un�3W�H�k���5+�n�%�!n¤ �C1�#����9ʸX�Yb�)m��V�z�X�Y�MQe��Ӟq���ν�T<Lqy��ns��%��Q:dr����N�w�NXhx�9�d$��=�����N�yٚ]�m��6����do��LwI�C9\�]ҙ$�7�]�<��`��8�K8x�'�̙�=F��6����WF��d"���D������0X�_=%���"��Za/Ǡ<��t��� ������&d��y�-���.u	?cf��,������~���tC�����/�B���4)[Emr�CK�Ag���<�B���	F���0V�|T3��2б����٘��cO.�"��<�&����vW�j!b��}�T��I�=�Ʀ6Z�#���>۾�����H�r:ʞ�w;�������n��
D���@���)�]�{���33tJ���`I|��>O����ˇ��1T ���lnBzkt#��"��]F@։D�w��G����D�
3�!
��2� ��S�wץ�Q�S )^|�`f׷<tp�_�F��j΄������j�L_�=2���H~p�vQ�F��,�>ތ=�]���svK���)�P� ,K>�����,&-� D