��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjfm~���*ש�?PMOAC@���c|s�vR�c P�)۰j��\+Qvt ��L�����s��*�U�Ѫeڰf�G����ܓAKܾf��/m:r&w�`0��{��M��=�bz�y�[1(�Xl|�%��ٌ��� �� @�'���E0�-�����ޕ�a
���R�g��n eP��� �6���>�)�*��^�%J׾����l,��zMy4E��/��&=L��a�m4��N⳵�C5�8�	��z���EWT,G�.�c>�c\�����u�D�n�K���������|+�3"���P�zI��Au�E7��/�e˻��6�Ą_���I�AF����^�faV�ϵhxPM���_���J]���G���J���U�F�Q=ID��JOT�P��{%�0ӿ�KA\X����˶��@�+�4x`AIu��qĢ�1d��K]V�ڋ���*4L.?O��7[�G$��r��k&]G�G�j~��S�`��u<��K���rn�OJ٤!t�"�(3G���
��<�Hn�������fӥL%�gp@3�1QSoӂ���2�m�XVJIH��a��A�*
�dnW"nl�O�W�������+�n�k�{�I��Gn��:A��}8qw�K��Nr50�j}�j��	%U_��Xm�
DFO���ww�Ql=ݩol��'
��g�&�Jm5��F��h(]g���ζ{��m�9/����;��>U��	+��C3�$)óu���`Vm�߉��.P��T�r�]O��۳y��'�n�Ȧ�),`��G�]�G�֩�%����~A�6K�� 2���oc<]�iz1�~ϞNRu�3Y���HL̲A�h�A�l�%9cX��9���dl7��6���ֲ��{��H��C4�d�c��7�(ts[R��uEDp*��)�p���f(N/�*��/v`u�P�� �^���<�V)\Ldps#WX	��y��� �𾪫����ر���.J;��8���ڽ3I�׷Ï����C$b�e²3[EW;�)����5WK���Z,�g
������o���%{�!|�a��(���h��*w]����S���ٸ�O;ĠY4øh��ʴc�^��ğq���I�����W�Um)��v��{�����7;�Q�ɭX�m�ѐ�n��d41�|�7D�5�^S��d�5��R�-2���ȭK��/k�,"V|��q���k[�����Te����ef��f;�P9�Pdq���m�W��K|�u�|L�h��R�и����S�_W��7�������R[;�A�o�Z�7f���#���%n?���_���$�PB�@����l�m\�A� ����-�ak���X=�l��<�zdo���w�Dl��s��`(g��ׇ1Ra&O-T���ˋ�.�z�j�ܱo�Q �dæqwr�,a�����v��Ùҝ�`@����p]��;i�v��A�`]F%��U͉6:Ɨ{I�;��O���t� 0��a8��@��:���Ǎg�unO]����~)w�,��M��O�/Y�Qv���U��j��k��/0��m=ج�~����Z�B�����d������rE�e��x]z7v#�%u��m��<3T6� L��!&���{�N�f���V������G�P������ؘe���ݗa�z�м��,LX0�_r(s���u	Q��|J��>�/'����0��^�#���%�O�9쁋i$e�M�ʉ�K�"��md�#l�,l0 �ȧ�s��wc�k���R��@^i���1T����P�Ce����`�Y�z�^I��`X��)�)4��'�I��p���`�b��*\�$�Au�>�&8���˯�vJx�漑c< ���K��+B�1j�6X:߱���+{�y�s8d���F�����)�>]oS�X1�Y�ar'Cu�(<3~�ׂ�ћ��eib�b.�&�]�f��JU�r8m��jQ����4e���Y��d���$��,�������wq��(��z�.�Q��=�Ƴ�v �Z!8WM�W����-��A�1ۄ"�C������-`�{f��/,�>Kuʎ}��-�wyKy�D��#�q��vϐ�y��}��1�o�c�<�7N�>��c�PV�x����Ƚ:�FSX��>�=�`?���\ȴ� U�Di�-��er���x��7��$�JZ�0S����U���^eK�0�����9G�YA��yK����=<�C��.����!$�Ò���a���nʹt��E�|�~���
G�~FI����R�x��I�� \� ��֡�^���/�E�*��:�Α}����~�Z�Rl���p��{��e#�b�؏�9��v��f�?=R �I4n;���_��]�'�t:o���L�3��D��q�2'����6tR|��*���3�HA�jJ�~�@��7) � I��y��tF�m!	��v����X$(_�<y?|�b z;�%������>���~�b�l�j�>)!�����&+���7'��:�Y��p<��Z7.H"�d��:=*V�Y��r�t��[�]�h���^�>��7tb���v�!���8e��".����th���0'-jc0p�&�#���}p�y�smu�{P�Y����p���V�}Y���̪�k���ԎA+zĘ;ȸP�J��J�&+����.ú��}1����Bt�d���Q�`��QY�0���ڰ���bº$��~�99͛8���u_���,�X�:�FC��B=�@��	�9B���_��+���8n�[%Kuـ]�H�f�,Z�2pU|n�o/r��͌9).ި-�� N��an� ή��cg(R^����u�]E���_���Y]ࣈ���6?��P��o���ׄ��#\��.22�1�	�V�g���{�shp�i���oH[֢�%)�s�o�E��4���D�������V'�~�z�D��94���
��p��hխ\�z��Ż�j����p�����BZ�*;,I���Ӣ�E-J���5�X�q�r�$o��yOv0V�:a�lk+�R�W���b���졠n�R�%/x6�A�xB�X��)���ǆ�w��E����7��2�g�=��2ʁ{U��`W��!¥HB�T�*�aSi7b��@�q�S�����=J�/s�\#�3�$��|�}�7I�9�醳r����fG��r,�)G �X�u
]lOqNW��<��%xw� gK��_rd��f���Ĩ���?�~�<���N��[܃{�Q�H�0���yB�b�Q���X��a���z+��s8�	�=�����eR���� D�T團m��ɗ�5]��Q�_�ަO�m����sjUt��Z�.4ձa�p����{X�	?g�raHC��CY���jC� ����
r%B���@��+�y�:�s����{w�52}�@Q]���4TWԄԫ�x�'�u0��Ap��MȺ��U��L$3�t�갚*"��oh��m21i)��y ��â��Ȝ�KJ��Ė�>p�)2��漆:�Y����
?���w5+��*���b��A�Ui���m���i �@Vd'x$���o��翳�C`L&�>�%m��7M{*���K���3�$g0��=� 'Є�qk�n�:�uɁ7u�(go��k�M�ց�me�i��5-��{����0TӰ�b�Vߖ��v�}G��CPQ�џ�/_؞,�Ĳ�o޴�GNN����:�WQ��6�����Ȁ�)���Ex��*X.��:���8�G�|�ͻ�_!��Lw,��� G4+�ĲV���%{��s�\K�_G�L�)��z�=4}Aq�"�I+C��y3��m���r6�ߠ������/��d�A���,��FC�*���)�0@P�)��3]I��*y: I�Q�Ƈf`�H��b��ġ1}ތ�.���*
���m�>�wHdK��B�Y�iή�m�W��rw~*)�Z�X�i�˼�2�F@J+�v]�~r?Ͳ!�H���$��u��������r��$ؐ�0�\C�ƍ��# �7>jo��#���<������\�!}J��9l��}j(u�,���E8��q����T0�(�.Q8;N��أ�߮��,q!1EA���.��빹�����V�Wls	[T�?�=Y�^���K��Q<jl��ە^��H���-��������
�u����z�u���D����w���i��ڑsk�RGL+���y�ĉ��J\U���f���X���-A��(�z����ɤ�j�=3m����GnI��ů�� E=QU��n] eѣ���|&���2⁅�ygD�����p᫖r�����-���t���F���&��չ���s�3f��+p��9Ct�Y��5���{�%��9Cɋ��_�1��d���/X�`��!<�L�zA��a{~ HȜd+��޳�P�GN����#��.�AS�.?s��F.���EH͝:1��W� �*D�]��S?���ظ�!��S�)��&��n�(9��*گ%���M���7P��1�����?$ݞ���a��u�#�K�^�P�5��>'���r�a����~��3����8���':�]=I�K�]s.�9L�X���:[�8�fU�|���\�c��]�t�/���E��!ɱ��y��>F�c�r=�.9���>C��� ߜzYf��߱��+�\5��5�as�����;5��;�)^!���:�Ǘ/{m��*�*�<Q� ��W��w�]�Ct�4�Y'�ȭ�C�s|}���`͟;���j>*�	�F��x�~S�'�5�Á&��2г�Lz�xy1���HQ����֥�B��4��(JS|IQ��E�x�֏�u�7sv;[Ov�����2�������]��[�B����1�-��f�0�;�H=�_ڗ�}�Z���SkYж�a�����d�� ��Ñ�����8ֳ&�Zc���<�L������q䆬�*i)���X��{�����$��:�7afm��}A�L%H�=�]1�r��d��� �T���_�y�,X�"[ȭ�嶖����d���x�
SX�MN�i���٫�qy��W����v�s�n�`%̔[vH�3ʻ� Q꾞at�"nR�-�	�5�}�H�Q��YF�I;��.�!�
y�|��t.O+(�R�X�x{���
[��e�D��݃YQBė�q�vtʿ��O$��I%�F�.�o�A4�C\9�hO?�����hٔ�IV��q�Q8	��� �s��=�=x������M��ێ������@�F��(�h�w��"W=���I*��6��}�d�lBӯ~H�#���f�GÖ9����*�6z�
�K�ر�������~��J�a�!��3d��^���?f�1��N��^���d;rc�q�s�B��"�e�ޒ�\Hi���y�3�Vy�Y���9Lx�JEB�����W���/mO�#U+��z��4���g8��Zh���s����,�pfU��5�am��F�����X�t���%9b/���٦�F��(��:E*�W�?xydf����%'~����X⊧`乫���t�;�<§�'�d����cMk�s>��\�qҒ���j���p����b-�֞����A�-�sP%��@
p�a����&���3���z_��3��=̲x�66;d"14���%��ʲ���rV	����4��WF����G�EӒ?]�O�f�r�i�d
eĜ��-�(f�K����x�C��m��� ��z��!; ����zu����b���l�o�d�Ő���#_& �� *�Vݓ8���2���o��t�S��XNg�n�LQ^mo#PY5��%�ל�鹱=Ѩ^�� ��0s�25@��F��
'��+?(�-��o3wy)�O��`�_���ؒ�I�g�v��W+�$��A�i3ՙHB�����\�1����aDj�X�4�Y:fEZ��a?�誗�R�11�)���:ѕ��V�-��BW�H�6?l-�ٝ��R;����5'~�(��O�q�mN��re6�脙.~'����� ru�g��#֨c.$��N��^5�ZǬ�&�f��eV�<᧕��\�;y�]�y"���^B-��CQc�Ĕ� �� _or���~!�À�/h�W�,T�&.d�L{�xΜ�C�;Ih���"c)A������F΀���x�T�\*q�OLc���:<hYi=��'i4l?�!�B�1�$)�!?�Տ���)��=�������m��y�Պ�Y[GM�^��i�3��1�.=���}�JR�D��I�$G73���!�]���Z��fݤP�* KE�5�7,���7�PE�[���a`�o�o��sFh�\��)2D�ؕf��C� �)���Ճ��x�a���X�X-�"�"K�/��� dd�R���k��\J�^�A�GM��M,V�r�S��lb�! #hsF~�3����d�����=����cN䚖�8 ��i��}��4��4���7��/�C �~�����v�K�H�"�����sӽ����Ȭf��gJ ��ˌ��M��zS��.��N�8~�5���y��=�,��7�
��2�:�}9��.�;8�	KlJ*eQ�Bd���#�0�V���P����6���7�=��x�4���@F�.��$�OX/�j�A,Lk��bC1�8@��T9����i���ىx^:�z�W�:G�z^5`����.d�%FD����1���iD<�5 ��^EϽU^��/���ޓ&�_�:����S㖻T��6�I���ns2E��3�q	�Me�����z]n{슡��^��߿��7>��˩�,Uq9I%�~���0{�'�.441L�.y���;�M);���&)c[���Zf���z?���!�z��N԰g�5j.�y�OFRn��+zɜ�MB�H��APu3] �n���ůGp�3�R!O܇�4:����p߽�@�zب,3��U$��M�\?�4�OZ��#/2soYwX�_��?�;���tV
�/6��3�E��~��5�I){��T���D��O"�9̝:Y��C1��� �"������Z;�M]yc��5f��s�G$�P��}A� v�>fߤ�����4���[�OWg�u��u��b�U�tv��X�P��v3�/�M�6���}a�i���oU'���-y�& 	*Kv���'fZ�4=��#�,�������^|���~�p	�H6���kd%�k׷�ЂW>�=C(VE5���6x�F���ٯ���z�w��#s����I֙RH��A��b��ݐ����ج�Vl�u�6���
�� \�kH���e�SE{؍7͔��	�Oc�&��$k]�H�����ݕ���c�ե�����1�$�@�i�I	#^43],��p�Hef�nf'�s����-�WkD(����������N��LĖ���t�5�3CʋC ���e��]D���!X�u�=4�7�d�8؇�Z����f��7Sd��+�#�(�F�M��3+�h��ۧX�D�?*�,E�B�J�E�e�ndu9��<�aN��e���R��0��� C�@d#���s�JW?��wGr�sQ�ﮏe�L+��3[s���?���:;��tb�)�@mmj�WaL�\�!��O�bM�˾��u�:�Lݝ�������>0���Rt2ͤ|^�&���dٞ�� �9h��)�.�l�GU��p"Z���$�Y&�*��$�S�/����Ǎ����@��*�cM��Uqk�6��_]��ghѿ��Q`(�������	Z]�7���׸[�t�rK>�S.�+4�J�G_!i8�g_�1�Q��a�����1�vĔF��h��Zf4�nK l�e	z�:%(6�R�]��G�X�d`�'���!����1Vr��p�����"R��_Pkq�`D?����i�Ŭ�谫���G�^�r<��K<��fx'0�?ۣR\��p� �2"f��+A�\����Y@6 {V�Z�7�h�:�֛�&��&^�&N*��Φ��o=� ��o�~Cȴ/2V�$^�RN�d^����@!1��O��Q�P:0,�Eq�/`�"�B�\7����б\�[��v,�qs<�S7�U�q��<���6@O-M;K�m�{�55J}�=1�tj����q�eC��Z���Xs���ºuw�2�룹w`��>7�%N>��A�q5o��٨Ў��P�
��W��]�[Es�n��8�Z��L��}Nb�N+v�O�Ey6L~\�Vi������D8���* E�d�SU� ޜ���=gJ-�q�񓚱��U6_]T�n)�wq$���-�ϧ=m'ĝcWH�%7�����LI��ݡ1�G�=2���ϼ`�� �hg�S��Lds�\8��뱫9=x������lFZ�V�#{�Ŷ�����#�e�y�6^���1Cs�����������r@�����NӅ���b�C�]6G��}|WM��P�X6�4Q4!� <$��o}:�С�f��I���0
�H'��XN���g�(�]uD�ȍ�O�dU�e������OS�}��Ӷ���߲��FqLy�>����a��U+_@KѬ�|�gLI��Ҁ��U3Y��3��r��"r�uw��ǧ��߶R�"Ag��L��Q^�Ym� �2E�_�us��{��/���[�jo��~'q��ⅸ�t�b��u�s�h''��RWG�2
�
�L:����=�m���J{+o�� ,'�����k̘|����)I���+��O�~����d0%f9�F�ω��)&(�@w��p[LO�{/���;�<:���.%\��`Z���9��A��,U:B�3��߅����z�
��$J�%Y� 0Z�!ࣦe.b/"�:P����G���˓��ʵ����?��G� ��-\AJ�fO����l�ǃ#�v�E.+�H TkW��)���^�㉨����<�8N��ca�S=��p����Xmt����2���,�;`�1�f�{�M8?��)^�C�`5�V�1��u�KXá|���WWxA�$��%�b�o��_���ꟴ��m���,:�f�/�ї�G3m�].�9�Q���s�.�a����зNP�/��9��3ԙ"s�
3�=��h�֮�2?�������v]��E}M\A��$7��ȁ�D.+�X�!��ڢ$ڱ�xI���|����T�w0�Q�)H@�h�i ��ik��E��.r�X��<��\ec��֯�d��6�4J�V��T�V	���:_�;����k8���ۗQ9�K��֫�¥U@�|�s�ܼ�v_;Nc0J�B�~�p���ް-3��Q3,#���G`���h�#/HY�:�<=��3F��촚��n:	�As>q��q2m�C�X��̣Dor����·<�	a*�`�u�d��%���_�{��[m͐D�ˬ1��6-3���6���ې(hW�~��R��Z����/ݑ-�c7�_(i��� �]�y��8Q��_e�>�m�J.�5/�^�^�2$�:�򱂛�z�Vq�BP���Jp��s��@��'D�X���\a��/l(=-[��:�I�9+<t~�����r��2��[��iq���ȑ<̍�߰�)�c�D|+�6q �b���1 y|�"Z��j0������O�Ϩ�����Sd��A������Q���z.�j�Q�uJ�ߑ�rPx�Uj$���6BU�gV�������2By̶,[����FY���;,Vp�tUi����4I"�d��3�,L��ԯ�u�RС��12y)/jA����|���Hⓤ���C�!B����~��+���	N��@���R׏�;ey�q� 6���+1���4q�)�^�����yG�>ĕ1X�7>ɇz�����9��Rc�I�z���ͩ�/���3��c�9EXG��9�e^�6�x���1�G�胵I�1@~�^��"�n ���/����OR䷒'���}��	3�s��|���#!���.&�Îz�Cr4�r߭s�S�<1!;�~���^M��Z�l��o7�xE]e�j~Fg��9��)C��TN���6�M�ֻ�i�Ղ�]�zgl�Ҫ"6��3g�Y�K�N�,�烑�F_���A%��K�����:���y���ENw��^����m���kAPx���Z1<�.g&����ª���d���&	����)��|^��vʨ���'���4�f}��<n�$tv�H�zkS�vc>R�덨����v��'<|\	�����pP���G�H8�l�1��q,}�K���b�fe��`x���T>s��-����j�����8ƹʹ��J��r]�|T`�Q�Q�&�pW�H�{����j-3���_	X��x門������)E���/��Ċ9\�����5���y���%��&��Z�{�8�f7�ƫ�~��y$���4��� ��`�P.��*"T�y�4bK(R���a٪����C��2:��>,��y�y��s`�S䂱�3F�ד3���ӱ�����u�����'9��# �]U��	�5�8=:�zU�����)�[ʠ�,�p�j~@OFl/��z����źK ���e��[B���!��ӯ;���p��%�eJ@W�(�t%��e��k�E'�!t��8��e�-��D$wX�����T�FB��(��݅�q�ܲ������ڎ�zVd^�i�c��J/t�Q�m�2Ѐ�����m����f���+�A��S=лH����=ԊT�"|��_�I `8/8�cd|�uԳ�M��~���J27�U��}8	#@y��N3�1�s�ۜU��z���e�{�/�����z����n��M��Q�Fh^.�@f���݌���o9F?�۬��J�;�J���I�d�TWb�̺�i��Y���t��Z�[M�]w	���"�ɍ,�r�!��F7����Q+�����ī�5��RO�J4n���ά�Wp/[S���=+�v�Έ]Dw�}�ϒǇ�lV�JS�n�W8
ߚ��V�+�
���ak�!� 2Y�9��O�K���#Alj��\*�v�J�O:�������Gj�l��|�%�-�h�k�:	�'B	{�;�9��Ϫ�����O)N˺mJdR�d�T��E&MO��qK�����	�8�}�P~�As�&�|��߷�5�%?��Ҟ�T��lC���(]Itw� v_��9O��B���tʀ��:t���,^Ѓ^2��du-�6�����Ч����W�`��2�����������:�T�<<}|�b���n�<�vq�� ����{�~��Ԯ����9dz����yA��J�Z�U��!��\�7H�&T��)�k �)�KO;C|2��~��1�2{�h�s\%w���T��gTœ�
.�Rq���ic�k�[h�WXb��F
>�j���"�)/��z/ſiF;�`�u���0�M�5�F՛��F��RMH�@�"����(�"������j�|�u����F�c����vb�qS���ǡ�<cS�,1x�h?i��ٰ1�m�Va�UҬ9 e.$2ֲ�o~�i�͍2�^	%��Xma-�r �U�\���Tn�ڊ�/����F�pK;��ͦ�ɝ�1�S��9��0�#�v[��zXb'F���>	�Y�)�W�\+�Ĩ�y0�9��@0���4闲���e�Y��pi~���2L����r����cs��3=���i8�uIG�m����U�y�f1r/vvS_�I�s�QY�Ɛi�G������jˎz��;-@U�v�s��gH^=�E&R�}�v�*��~!�IG��q���0�R���b��AO� ���j�O2&e�ʒWұBѰ �\�0v`��: �����E�ܧ��`���T��x�冺��N�lk�=�W�87�[��&a��y�I�~@�߯���J)e�j�U4�?܂�m�@��ۇf��5�d�lt|X��[;k��l�S���5����t�콩y�%�wE�)K����V]w|]�3'md�+��������׾�T��:H�<b��ى8~����h�"��������P�z# xE�u�{�l��]��g�ǇE�+�/��#H��+:��aG�pp�lrbD0,`��%e���QR�K���W���̮����
BN�6���t��DWC�����Q�Qn�/w�H��;�aೡ���R��dm�Q LA{��H�G��f��yks�D(�߆���(mG��5�c�o�ZY����[�5��b���H� n�&�KWצ��~���1�4n���̟�����)���:Q<�}��&��l�&|[���$�b�ߍAXL>�ʠ���|K�a�O��Ȭ�}iA�X�ɨO��#�ɝ/�mSe�%ġl�����d�D�R���8�<�m��y�f<t��>̋M��a��]aA��
��f��>���U+)���(��.�+j(�	�������/���Rx&�b!l�ɫDVI�u��x�����˅���Nϼg�kذ8�tM�S0�.��Ӷ���º_9D�y�ږ����;��<�q�����L�*��_R�ϋ%�b>禕�W�)C�]�.�>���R�q	��g��p?���6�sM���q��U1p��#JE���{�0fB?0-�����\�[�֊��MNc���;���	��W0+���[Nߐ�	G�j� 8�丌ݍ�C�6��/�-�T�t�Ƥ��A���F=����bWA�c����Z�r+�"BD�3v����x�~��~��f�]hsU9�)O��uY�k��=�h��Q�Ml�-�KUk0'O��o�E�!!/�L�6!{���(��}�p��o]ͳ(��  ��k$��V��O=�=��+�Xn���oDJ��te��l�P��MY�ҷ`3���K�1��U>�*��2l����~�b꫐�xϱ.��WEf>���\��R�%����kk:�؄�x�<۷߰���TضY����)��m�>v��lmk�C��q�;���N9+���(�N�p�*JX�,��2��cK2yw��'q.��m/[��y!��f>�z��/�|&�8\{���0�9�()>n�v�3����e���w�=4E�%Èk�����<5�K�O;�Ҫ�i�q7�)��됃w,���ʭ67��7�ӿJ�������n���B���/�O��8�q�:� �uVm`:��Ɗ�U�ggyQ�_;V�; �~*�us��d�[���b-��PDxrґS���շ���*ag��06_+ ��e� �*�d��(��m�D �Ό"�������/�����{B}�塗�3Yk���P���	|��� �����|���3H�p�s�W�-��%���O��5b"����U�������n�y�˺�`���e{�Ŧ�M��@��?pb��p�+����Ü� �0���K�C&f�C:�_crj�ڒ�+f���(��Y� �u�M8���F�	�9�p�s�0x݉�h����c5�2��~��P�f���`[g �-2�4t(��"��JR|��e="d��O��H�!��[ϲ�gE�-M3�N�FO�9J�P@۲�4!�m5,PF���8,z٥&�c��%�����|y#�|²��ض��p�7_3N��<�A�/�����BAp��Э�	2�7"��)�Z?s���X�J���[%l3l���wa������E����e`a���:uh�����{mM>
៳��[�q���y/ѳ�4W�ޮ��u�a
 VР૎���0,"��S�Ҝ3-7�`�ZG���Mڏwk(l���aj�U�A=,�uQp־:$��f�n؉f�C��A}�a�� ��U��5ϧ� n��� V������ʬ��E�/&T�g�}�mɉ2pʪ�>�\u{�6��n���Zb����5�;���v@"s�	kv�ZV��o��
8)���ZfUǩ} �
�ġFf�HC����7Y�C���g[�Z���XJH�4�8`�(�߽�#_�3`���i�ϒ{�L��%x`���	��nZЉ��{s�ͫgY�ϝ�����-��e̘s� ��@����s� �R�(��"X�Sc #��P2ƀK�5��ʉ&�-z{Vg����Lի����L��;� /�<F	�;ϲ�K=�|7o~;l܋����*Ig���-�'!�Z�'����%\\�g��/B6�[A�f5�q�`��׫*�<~��}MF�@`�{l~���j;��s'A�p�(C���SD���7AU�C��!���j(6Ԅ��c]� X��J~�@f7�̓8	�f5���[^����^��	���>E�V�~Q$�t�,J�����Yb�W><h�NI�b�x��~{"����@��V��
�������ٳu���g��8Q�n#�����*�NnW�c�Ω�޶/��
)��ݙ��i�� ��lś����p^4`�XsG�_*W8f*���O�{;��P���o���o(�ǆ�K+:��E�M���nx���*��fs�}�Nza��;^qp[m@�����}�rN<EQP�jKE~��D����ePB�]Ha"ᴅ[�$��)ꥯ���/V|:вe�(g衅iY��Q5(-���x�Y#o��s���yb(0R��Q�(�PtZ��~��ŧ�zU�o'C��S������}�|�ĉh�z��0~r�뉞�*���PVݬK���f���:?`���� h���T�]���(��֔Y,�8z����*A���z��X�S�;R+;8O�*#4vU�}ð���sl�%1��i�^�i~�Bd�Rp���rG��_*~�a%�b��'0�� ��l�1�\S-,ߔl��
�F�앗8I��X,S�19�Q1���iX�׎����C���C/���Ҕ����M63����Aڞ��Wb�Oٻ�x�zVW�o�f[`�Ɩr¼�3���l�8&,�)f���@Zv��e�&�d3\�o*��	���Z��27L�#��
����s�����	�(jd^r����I6��� �.++I��z�<�:|�Ϋ�b�*	.���tӷO��[����8S����B�a%��w������5Gv��T�V���y%K��$ԭ�H�>���#S�[����g�,� x�ʲ��� �1/&����	���v9�G .���W;���a�oċn�8�qW!�1[���E8�x�I�C�aTM��t��ۘ`���5-�׼@
�**��[���߃����.��zь��\m�������s��'����A�bp��m��ƀ��a+��0'�y��^��!�	-�È����+rW'w'��mB�;z��o똆L4���fq��]ki��^�r~��z��[^v��=�i��N�5�2���Y]Ơ�/���&J�r7�rh�M%��xoR��sX����\�'غw��żL�T��pZ�k������&	��h��	�l�_Z"����p���Ǽk���j�f9-łF�,5������p�/\��(Q0�vϷ�o�SPKK��D���=QWE@TLͅ۴�����b�>�>N�%@��m\�}�o��b+h����9�:|�#`��U��]6ǍR��2H�Og�a��,0փ>�g[f��{yh���3C����MQ��i�'ǯ��W�.�tpz����!��
A<�O���f�+*P�%&���M+FUr�!݀{��W�
�WC4�GKlPfLM��7�ؐ�����̪}q*������޸�;H���WhK׾�����FGz���vxG�PV"H��P��q]���ԟa�D}d.֣�,��Z�i�̞L�38t�w����4���W��`��4�P�tkpc?��¡	*���x`Ws�+�_�	*�1�S����F�.�o��T�d�D
2���nW��zb�n��b�����k����bI|-Di�2ƈ�ײ��O=��!D_&��1\ￒ[�����?�S#��L��l�D�����+������?���O�~�8H녵��Xi44����a1�����h��ۃ��G3�&���?�(��R��Dh�6��)<
��E��,�'6��R߲�]D�d��o���M��@�.v�G�OF����Yԩ����I~t�u0b&>�����+�kGY������$��*~u��"���e��T�'��s�	U�6y��
�(ˮ|������׮Ͻ'�F-�E�|�;���n�>���F�� �P$��~�g�77ʅ���7r���BWѾg����[e�b�ݼ�(ѿеy��a�~�DGbٓ6ap��v��:�=^U2�������l
��!���f��BQ��gY�u�G?�
8��*�x�{�t�L�}v��o�5ʵB�3�y��H��]��,-�=�W>d)�R�ʑ*��=d5����<��(��t��J���E3ب����֦~?,m?��yBw�D�J9��?���7��Ea�-����
��fߧ���&*�͍��Rx��u3œ�;����C8 �D���U�z�$"Ek��c�J�����cǻ�*���ߟ��է�F�5_I�܋�9�� �=�0��k��ʤ;gu������19����f�@�B�*��qU @U�:���!�%AN��P�7����Zjv�� �X��wܪO�h�&�^R�i�R�{�p���K��-]}�xӭ�>���r[�F�`�* J?��]sO�D�U��^�<$�ۗ�L#�2v�������b��G�#�<�fx���gp}L��~n�s�Bs���~hu7�J�A:��U�Hwo����k?C"��)�,��J2��D���֨ld.9;�N�������n�uqc������_ҽ�[��wt��^�B�L���.�����sa�f��^n&�d��ip�G�E��ӱ����8�s���3���C{ֲsZ�_4��.�M9I��rՍRo��:�F<9mO:�R
Z9�h{�IC�M���nӒM�y�Xd=�1�Ɠ���V;ι�		�:�Ӯa�G��Od�c��c��%��Ec�,�Z��\y4g./���2R�6{��A�@��ܯ�pD�y���6�^�G�Q�2ܕ!㲛�$�o���@�E�)4À��n�jc�xD�c��V�� M��s�%�F[o��?4�����S|^�gT���$����0OF��f�����������U�F/�4��FEh���}K����S[� �܈N,�V�i�T���J}�	Ú\<��9G�rd ��GE���yvv��u]x1�~�cz"LɹH}�ٓ�G��J]U�>�6��?H�*��������\�!���G��hj��!��Xxz�P��j֞Dc��j)�E���"��E�[��-�~�p�p��qp���Vgf�������<��i�;��B��v2��w7�2ZM��G��ˡ��r���)�Hn�z�*�������`H(�dJ���f��[�dJ̄E}��\V#�����|��ibK�6�<��w3(x���j��y���-��v&q�Tl��K��dg���a\�nhC������oD���U�� '���P� �#TprN_����P���o/\k�6T��T.���Y��~rY9�h?�B��>4�'cabmV3��:8JpP��ʼ��K��f�����W��)���:��$a*�D�S����?"���O��]�lWM�[UEA���0�i�3^�.��������]������V|@�Ʈ��OH%Y�7���.v�Ư���LK$��B�)�ՙ�ζb�_6{���w%W�pp ��X�ް�܆���'a�z�(�$#�lx��7��GQ��wit�3$�AF���]�䣎���قUdS>\!6�Vyy  ?O!�ᕱ�=���py�3��W9W�n�T�2�bG@f:`�w���,��be�u�Y�d��N���*��#!,���=^E�J0�4&����ү�;F�Bh�t���u��z3y�U��//]̯&������'�D��@����C��>v��$�|�#�|��
{��Zc�ߧ�Gd3�T�Z���ٳ�����̰/l3Y�d��+!Rt�p��T!��������L�R�p���A2N�p�!�Exl�W�R�g��@i4�bdL8-N�W��3�?��N�r1w~fgBR�����ܪ��ZڟaN-�u���{ow;#+��N���d�8�%|�{��f;�vr����0�������x%��!�ß��L���u9�Q��r�����'�C�3��
ZSZ�
ܫ�����䟉ݭC��k�=�r-��`�@<�4��������h��B� �u�^��g'iE2K��L�D	��rXc��	�C��Q�N�����|�y29-l;q�諡�N�B����ʤ����_@+ۂ�W";�x���1�D�߁&�@�4ٹI\>9m��#κ�
�`2lfd���U��C���H�G(x�A��d��ߒ/H{u�qg!m�R��UX}�k�L{��*��6 
� ��0��Vc�A�ajl(�B�{e�J<N�^I�L�#�u���G��M7���5������G+�W&��%���|�
y�I�K��8����ꇸ��8~g������"�w���V�(�h�?7�VO����f��E��w��2f�?͐ڨT�N�s�E-<W,+��%Է��Z��ߡÄ�v���L��9tG;�W���&��mPD�v��&⫢C��.��͎3%��c����;xyB���!Oa�ԲI�� ��ɬ�4�@��ȋ;#Kq��h�'P���ltS����k)$�V����'���K�t�0@R�~_S~3F�x���X)	��
N��$؞�B����d8�Է�y�d�]��)���]���ס3	8$6�hJ �ʥ�o�G��!+Я���D#�>��Ȩx���9�
aL�a���b���`��7s���3���GةZ�t6��ވ��Un�'��MeL�5����L �:C����V��� �VC���Ե�޽:A�"Q��w#��ղ�g�U��0���*���t�a��˙����H�%��|H;�[����0���U��_���T�L�93N������^�x�Dƥ���u��+�6�������co��%Js�n�{��R���6e�*yI?%�hV�l���h���Xy+BU�N6��p��@�i�j��,A�3P�W͋��;z��>%�Ǝ�	7��J�N�y����l)� 
3��zTl�*D�\�6��zt��qQ4"��;5sX�؊G�d�=����d/E�H ,A�@�`�N�R���3]G>i0��6�-��v�,� `a�g�B^�x�A��>Gd
��̑+�uC�l�_�ݥD��/�a��p�L6�=�ڒ�X@�WT̕6�'�x�'��v0߽0s��̺|��4�e%�h�hJ}�т?_i��kBV&���F��#mN���+��7���*�W�.l�o�-u�כ��)�n O��6!�ܫ��)��chNw�b�b��{a�x�&�ea-k���d1*@��B� �D~c�|���P�`��v�D>:W��V~���XLr����BE/~�&ƍB�s��X�헿X�J��X����X�Я�'��SX"{w�M���sY�av�^�T(�Q�Mq\�K��\y���_�ܫ�c&U*\phq6mz�Gɍ�5����-sN���/�b�T���dn3�D�u�N��[����]봢V>10ܩb��t��p�������-H��:���h�?n��u���g�O2#Ċ��F�/����;�A�������s,�sEM�n�oO�����agT�l>�´K�E<�N 	���s��%��dl�z�d�?٤3��ϩ�W��P�<92dR+"E�����=��r� ���|V�Ú	��_F�·��
��z�S����y���nk�a��E�艩�`6�m#I>u���4���sYջ*����a$����� `�8X��j_���)�|ه��0�+��3X���*��6lu�L�-�ב�]q��;c}Qft�ox�����3�"�6�ٷ4�GV�yu�S�R� j�R�ն�w!4C�B\|`"���V䷍Y9ŏ�U}��͍}��e�M)[t�����Dy�H�3K��ɽ�p�����5 +��E�s�0�� ���"õ�A�K
�� �~��{�,e��0u�(�o�ZB@�o*0Ϫ�ԾE�bϹ��_7�ś� v���l�6ֹ��D�x4�Qw������3�}MQ.H���r&$�"����f��Vц� �\�i�+��!z����2+d���8��i| 
E�0�k�g��E՘�Ɋ���>>�]�"�OKlDR�Ӑ5ҩ��A��R��|WV�0�*� ܐ� ��Ht��1>Dܠ�B�L�dğ8��"�$�nI�LY
؛$��	�� S�$��c)�g黜��%�@^��D��[^��uS8j��fEL*�����
N9�qӟ���E��_�
KN]���k%Q{���R�+��G�F � (����J��w����V�LP8}���/�sJM��`r�^�#���("m����78>ojcP�b���_����.�y��s�C6���Y�����<-���)�q�7�3��Ŝ$�>��Uz�S=O��ޭ�����t���	9�u�i�	�ga������+��y�x1��d��#�Q������ R�"�s�ٙ�yơ�S[��)�(d�1<��V��A��%�l@�H��~�ׂQ���$�W�Nڷ���FS-�� ���$�C�xw�D�^�F}5�����м����+�� `�70��g�bxV81���h3~� >��ʴ�1q�i9}��a`�WC�����˽.��x�C������n�t������*2�M�-tQ���#R?�k�MJ�KO�n��/��|����	���ڝ�gi���#)g>[Uճ΀L��S`� ��D�>��0�wa�j@g�n���W�Z�~�H�F֟�@@���+�؈�W����@�nI�+�X,�H�]J������ʌ%����u�A9m�ff��1�|��R�􏁥Z��>,d}���ԉ[��ʛ.��&ۘ<M9_�'�c�d�=��O�ވ�����p\x��;ڮ2}�
M)	�O�Fʐ í�h��M�Y�����j$\e��\�=]�3ngT��l�s�^�A�yv��Mg!�Z0��W��C��.O�!A�(����y�E�z��+p�5z:ݩ��g	�=*�:Y��bU� J�Ԫ�Y�8����J���HV2�3ͻHS���@���(�۷#���XE�5+a�	���H`a��㰨��*���D��׻$_sKu�+��>���yL�T��YkK|���ti*5�7�+�j	�f6�d�}ٙZGE�K��i�U�AۛQR�;�\%
��_���X�ُ�t��C���/�e����H�\���~�n-��Ú_���vS�����DX������/쏶��V!�<�݄��r���?M�@����D���������,�s	�������S��*�>����+�1��i��1��@�y�N.�����m��w�� �oQ`���d�����J��=�� �����'�j�>r�C�6�tZ Hӂ�k�3� yZ�/�ﰨV�5Y-�5�����7~J�XbF?��l��Q��H(�{�F�e���ɳ�N�3'�]�O̔t���\�J=�K�w��Ð�'����Fȉ�d�����o"�m��<���P���`T�d���q����z?�����դ}#���d�r�̊v��|B�"���24't�7jx�;��6By���v��<���3�1F��j��+En�S���d����u��/����,��>Ơ�f��̽v�K�W�b��å�ɳ �H�"�d�?ir���}~V�0�w vba�\_�R��-i4�y�fǗ�R��56����T׍�!B���dyVN�Ո˦��'3�����y��]�$qg"��M>�� �w���,I�ݻlPl� o�V�y�)1�kd��i�������c^�����Ouɾ�TaLU2��R�_��:�U�?"�7�@�NJa�G�C�BRh�Ty���H6[1=�c�\����tꠈ���.�l����NW���WI�}���ه�!b�G���d��7g��}Y�g��K_oq�sFb�laӻ}�tF�y���S��-���_��z��3�~:����7�yۚ�\��G-�@�#ɱ~YL�;�e��o�1�_�������E]��Y=�A�E���`9���~�zK���ކ�0�y]���J
��oLh�Q0J,���y�b����t�c#NT��%_Ʉ��i�pP�O��a0�D���$�����=������/�8����`{� Z4{}�M���^ؿ��4�[��r�2H��Z�+����d s䍞~�����K�t���y*���=ȳ��a�iF� +�2+�4�}���^5%�mܠ��$-������v!8����������I�C����
9X�x܀��o{�s�!è��_[x���* �&O���_
ja������B��yqVA�
�p�
�B	D�:��[I�|C�� ���օ,�賎X��ĺҋ�CG�����k�C�Js�2歼� 
ʒ�r��:�ȗ�#X[��O#���]��[�9���)+Me�����	� Ϛh5�ɇ�z`{2_[����r�g^�Q����3P�[��� mG��ըF�Ө�iA+���5�X�C���*�u�~�v�Y�i�4d�� �]��R��UY�Q#�����߇;" Δ�h,��e[�Ķ�'���F����.�g�ل{�O��9�S/@S�M����܍�C���$4��g*�^!�����7(V��B>\W��4n(� �8e3�t����E�Y��N���TK`�-�5d�Vr6Hh�8�D�T� =��E>������p���Z�qI/��w���Wym>�����y�;Op���,�@�M��J1��FҢ�3�3a���l;�H^}�V��L�)����=��댬��,	������ ���R ����Pd=�;;_�=�"[�o!�F�9��}����W�xB�&��Pb�!��I8��C����	ʈ0����0�;����5��h�����T����*f�e~%M�!N��1�U�T=u<7��]?�D�e'i�?�~{JU�k'����,�<*|,gQN�p��~\L�u1(�O���-y�(C�x�.�H�E�4F,�.�-&�7����E�;�纇yME����<i�'��	�#TT9ʔ{��X�)u���c)e�@%rpZ��GOs� P}��u!m�Ln��B�Ӑ������a��������]hJ>Q��Z"���.ua[���|�&"O{�>����f��J�))5noY(��0��E>}���p��e�5L�:�{k��#�e�j�T�^}�7�#=�Я���+�E�S��M5�.��Ɉ�5ɕ�#���O/��A,�	0��5�,yά�N�D#����_���U�Q�����Oް�a�}�|d��>P8H���}j�1c^�f�^�_u��u��W�g��me��,&P;�{��e���d�򯾝��ٱ �\{ԗ��b�Iȏ0gs�uڧ�\ V�â�)�X���8*D���y�Mň!�_��h)(Y�^A��ȳ�-�|k�a{�>S���n�'À���̎M�cXTW-9�9�;:)p.���y��47���γ?|��ZB�k�U]_����F��S-��ގ��2v�\Ee@(����]� �$2�6�o�4Ba{�Ǣ�5�6�/=�����Bð.��t�sr{�^��*����R��F�j廢�y�?@`w�e(��@��2`���w�*��,zO`����@�K��ݴ���HZ���'��y7������5kT���-s]~��9�U�4'򸒓�Q�+��G6Q�"g�a Z
��q�@bm��l��0��W����T���b+�x��qg5=��շ1��(�~�>��9d��DǠ|gW���|�R��E�Cr��r�w4��������/+�v�������������;���E�ɤ��9�+,��}�o�1�`<?�DfM�"���h.lVom�y���w�Y��{�����t��[��E�F��AhW��'?���v��n?�BV���󲿘,�?�K�#�(��k�����V�nAw��#?�e�F�Ё�DjA�5�w]��{9���b86X��+j���b��r�K�ţ��U�cH�0��I�V�8�֌��o��wIM�ʛb��	b�����t�T�e��/#��Ֆ����L׫1^��S��=IK2��]X�
�!/�ϩ���Y�h�����N�%����P�;���	~
�P��t��V.a���;���}��=���w�����j5�MJr�C���4�x��d��1�'�2�ҕHC���Ne�@�@�(|�C�؅�l�W�g�񿲹�=�i+��.~z�n���&<�QS�`Q]�JE��R�%f��|F8�Ӄ��1�J��T,�&3܁G���?�:S�2U,]fN@���K��BT���ϯ��Rj�/U���w���1��ڍ��Z�m�/�7�C��l6^|-,���oz
���۫���}[��lg�}�4p�ҰϿ�-T�}B�ӈ�V'�����K�R�"���;T������6{����3>>�o��94J�3�#6��~�zܹ���B���g`�o<�e����g���Xb�!����x�����ZnZA�<�{� z齜�3�=�
�6�)<)�J���"~�r������c}��N[b�P�L�-����7���z�Ϟ1����4��3a��4Q�;�J(�qv� �V̭^!�^H;���?�����!d����&�|ɼ�� �6;�����^�_sq���"�t� N����}B�(�-87�4��Z���>>!�$�ً����,��;iǻG&u8 ٦�ql�qI�
�s��{�?�ء�ESt]�e�6zʙ����s�[�ul���1:�k�E�F�آ}b��4a�|'�Rl�p:��6-4��갦����R�ӫW�f�N�t,4Ҕ]���=)��I��^��+u� �'W�sK���ۏ�☩^��<�D�
�!9� |��4����
�D��+��;����9�NLr����Y���0������EI�89��>������PjM����G��v;7��Q3���5�Q>�>��'8<��6��ڶ�T�f}χ�ȑ��1���,`i>���z�P��]���z r�x���j�0�[��	ٷ���Il /��+f�7Yr �δ1G�9�U��.�`i�fN@/��*�Aj�:�����$�m�"����ı�!����=]�'ŀ���=?����^mFQ��, ���%&r���Pj�}�Xq{	p9��TFn���q�[���{��'�c�#^�)�ra�-�o!���M���A��B��)_����RF�z��"�(����X��õ
�fha�0F��w 4��.%'o�ix#�HUqk�$�oB\�ȜQ�s+<�B���k/���'t�Lw�M�g�5����nF+��l��o$S<S���������`��A'���&\8Dn�t]y�*D�ؙ�(�uE��
�(A�.�C�&w(��G
�!�����@T[�U�ӈ��,i`�rLrU !��8Y�~e�&H�L��"�7c�}��S�h+�_HR`�4�������:�ϧ@i���U�M�9�8��3�	���?sLl0�	�j�#�3�ˠ��|��JMJ$	B���sl�s?�1�wxº��f��j����	��v�nu���蘠����y��UZ����]�<�n8"�8����}k�[1�.�)>�᲎WMY3�S�辵�n&Y�(�<`��m$�y��l^<0����O�m\�o�.cܦ�g�ֽE��	���k��T��%�!":��n��bz�9>�|��cg�'� HL�VQB	&0)��T8]�k&nň����ԝ`�>ۆ�Io�����
��VuRC�ߩK�89�>�8��mPd�?3�klL[qM�ImW�k�S�Ul��ЍK���r	A��K&*����wd�w'o��W,�0��b����}dN�dQC�ͼn�Y!��9s{�T���
�.�F��P��k�ei�{\�NOA��w��ر��>]�� �0�њ\n0x�G��uEQS�|�j���N�c���;��nS!z��ԣW���j#��ƒǱPA �^����8-�i���җ�4Q����,wIE ��
�S�<���V%^H�2��|C~����*���G^R,A���N ����>v6�V�u/gu�٦f��$M=y����M��S����V>�Z� ��B����%�����&H��P��ZN�0h�2��p^��HЊwɑ)We�c�:%��Z	SUK����?����.�W4	��2���:Z��U� �a"G��z�"��~��m��X�:N�	�6�l�zTDr��=�t�L�9���0랂�K����*j%-�.w��}(C5��(�՟��-��@�����W��A_��$�s��	m3��2T1kO_�Rn�V��o�WN��Cz��"�LY��H ����!X�:F�@V��х��=|1
=Q�ԡ
�k� s�c�6���G�g�}i�\��%�bŧ�Ui��~g�]%��b�=��q�M���S_�����Fҥ���`L�	���H���>��X���n����Zތ��L�L��\x٬#d�h���y�$U�l7yp��e��u|f2��&��Oڻ5_Pm@�B�XYʣ��q�I_16�� }�XŅ����e�sD
�OS����C�G��핪�>Z?�z!��T��K�͇?Z9Sy/�3�r*��禮5�x �spPM����0~��aM�\.N��	���(uʮ���L�l�fLo�ǁJ��$�E(����-p�cS����k�נ��������͉��p��
|-�����Ȩ�ä��s(V$��G��Ԋ���Y�z�x(�C,P����`��jN^N�c��~��?�[<ZtS��q�y<`7�	.�m��D:~;���' ظ�*CߢN�LXl���o�R�Ⱥ�hn^xH�8�-=S��$�6y���Lܐ8{�5�������٣�>܈���ƴa�qxp�#���g���1ߕ�y�!�'׫5�T����O;��^R�p�ʲP߭��J���]j����7T������:�U�}��>���0�_� �V.�����/ϖ0�G�>)>�n�	�\�(���nEI�*E�VcTN����^U�!�^7*/d�����TI&v���K�W	?vOIЅ�<+b7P�����OQ�X�y B�hf[d�Z\	"<Ů�eI���U�w����.�o-������'G ���.{�'zc��d�J���v�