��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�i��a
Α1S%� �uj?�L�3��TLei-3^5]E�$�����~�J|�<����Gy9�������Y�W`쯄��`��jA�]��EL�X "W�)�R���dF�4��1�����l��n0!1(��Bқ��'��������Ͷ��7�s���I�ެxr�t�Iu����v��D�3�<I�&���t"�q��~��b/P�<E��Kb��4�gV��Q+mǉK�.��
CЊ�d,�O;����+� Ok�m��"#�����.R�)D�jiv�ֻ+�; �N�1*�������,�g+�Wp3h��Rۢz8�W eł)����-����]_���_	�`�n��Ť�w���WN�YA�,�[��RX�"
{����3��l�C2������'��0�w�?�ɬ�5��R?�ȁ�L��Ł�η�~�Z#qX"5�W��\`n�X�[uq7�����xHx�DȒ�6�'�.�e��~>�a���*u��gL��h|�p���ߎJ��%���u�2ֻ��MIX��FNL:�r���߶DA@�X3��?^���j9R(�g�v*;��.~Q���X(jR�֯�r�4Y�z�Rùd��Ϙ�^W,X��g��=�I��&߰�oP�w��`B�A�Q��S�ݜǃ�U��
q���l��Wg�P�ߑG1�]��p} �iB�Lz/t���0ë7���.�a�:�&K�~P��&iav������)���΅A[VcȀ��^�t-"��2��&�	�,7���:5!�
K��h?���*��>̌��sh%��C[����E��4�Y�*�r4�R��)w�M���9Fe��cF�jG� 788ebƫ�OJ_m���,�r0Ս3��<=�%om2P��$A;a{�Ḷ��`3���Q��kr�cj��d�V��~S��RB�ĕ�$�%� ���a�BJZ���+���G�s�:�5o�\Waa,H��U4��'�wE��%�Wl ��K�݄�Q�YX��M�_r�ߵ��&D�r����z�	�JK�DwHWe��͡!�9-j<���A9�#�jVa�^�L�w���1]-�ť��X�U7<�_'`��4.$)��R�<� t���JH��D�ey���H��Nī�nTM�A�00� �N�ʹ�f(97G�VW�s�@L����OR$dpٔO�|����J���#)(|��޹p�PX =�\�9�%j��<�3�V�O��:ޕ�e9�Ǧ��r֣�b�D�m����݌��k�k\����G?X��u$M������=�`����Xu܅ǥ����G��o�Yد�-������\hr=L 	�@&�����I;={���������#?י=����v�1�rp��!��cY.\w��L��s
A�<�F�;4Z�!��c�z��X�(M �cL�ï���ϗ�n�tgmY�@�}�WQ|������5j@:��*��Ɩ���(8��x�JYC2"y�	Ȋ�&�� ɪ�@ J����pʷ���o����͹�ya�_Qby���5B��=>��qS�{�B(:��BZ�?iK���6R,��:.kn�a�`�'��c�a�w�%���:�����B3yp�vK�~��q��ʯ�����'�(�G%�6��#�n�TB,E���VzKl��}�yz�#%�L���c@�;Ӟ���j���q��
�u��@�����܃ft�a�Y�K١}�{�n���������f\���#O-�X�v1=Ek�9�MH�i0�k�B��ޕ�n�����Ⱕqi����tq��n�t1A�à>�8.�4�,|s|aϦ'���M�;*6�U�Sl.m���E㻆g���\��#�!RWDi��x�c��ByUU(��C�o33��}��O�+�k:�Y�~>��kx��ôQ�X�!~�D���u�R��m��*J*-�vˎ{�̜c|��x�sp�w��tb�(��{Į�#�03�@r��`-3�Ԭ�ˬcG����w����"tW�_��ԇ����,��|�J?C���BuȬ.�_;ZG����א�<s�ٿ��"�[���H�O�$��vN��Y)$!�{��xq�LotK��&vA>X�j�I���P���� �kn&�7�]Ʒ�{E�^*s*.!�q�jY̖�7DM�)��,�':ֶ8�үt�t��� ǻObp3J�����3L�IE���lW�k��7�~�F�����k�֔lъ�w���%��y$�T�b�F�A�LXc��>Qnr� ;M�ƒG������N.���J{)2T&�M#�M~g�o�<rXJ���*��3W������f�3N T[f�n�.L;�������I��_��g.����nڒG��٘��,)��
w�qJ��p�6��&(��Vm73z�S��Ĕ!F/Z�w_�oh��C��g(��2B�o�jw4���Zb�#�Y3O>�ԟ.u^ٓ����Ⱦ�Wt���l%&U��aN�Ka�(�ޘ�5iĭQM�� �<�I���=���b1a�Vl-K������bԈ'��$iy��p$�|ޔGYe�%��n���2����YM��έJk�i��Qo��wV���i~�.��p���O��G�L�Ч�ݾ��'rh!1�C��ɴ|U�C���>��V�5K �(��ߎʝk��CX��h�Uw���7r��S����C�� 3�I���8_C��Iz�F��}E�)aM�`��)�E�0���X�lX�܍��C�����K{���BO�o��~A�f �����P�p�qс=� 墨����N��5�����!nw1S�����j5xh�#��������ak嫝��~��Ϲ��e�6j�W�r%��^��P`-֖@���@���J���c6�(Y��˝�)�x��u����v��Nz�*.$�zJ8y��/�8��	h(5L�xc�W��(eol��xe��9�i��!�T���1�"�_�ԅ�˧�}���'��V�j��z�򟅨�!�'<:\��Ś%V�����b�ӗ��J v���"�.��`πl^��prCrYi=6���"�p�yi�#���_�o!׼�>���;����о����EZ)�cp�!��D2yH�g��S$ѣI�(�I�ɗC��Gx� 41U��S��T_�nNϝZW��@����d��Rrݼ̳�����n:�h=�ݮ:�|t�7����e��\ޗ��o#"�7ƫ���uQ.�5�	HѶ�Cc���l���j|È�M'���@�-�w��y��>�(ˣ��ݍ5Pj��Tеx�*_���w��2ҏ&�[�Rtw^�[n��n&����(��J�m�n[N�W����v-�@)8�] +�������՚-�l#8���6��;��#��A3#��}� �i�c�c����Y�{l���b�8bdъ��w��Nʗ&#ߙ�eO-�8�ټ*z��G��E�����8��_��Y�~�g��DF֯�w&C�#�C5��xR�j R�H4��̆%Ka�7Ŵtx�ĥ�}��ʐ�m�{�+e���oe'�� h]KR��ɾ�zeBÑ��3����B
v��!ʢ�%�I�vB_�� Y�d��P��0�α���+H�xϘ\���1��."l\���O(��/���B7(��5�I��0�Θ8z�P��^U��Z�-r�9�T�
������3�ѵG&��L��$]�=�#��a�8�� 7�I
\��?xDG��OD�� |��W5�\��?�"[Y�L�Ҟ9cr+:�����}�������E9��Gԕ!�,�i�:���>[�wEN#Y�Ƽ�h�$7�@��{����0��n��(o0��ձ��t���[������!�P���� @:��v����r�3XJE�6Ι��F{2����t�
��Z�Iif�1�(\��I�7�Q3�F�_�M�D7��U8�*�����`LH��Gl�=����q%���7Q��R@���G�f�*�S������>�W�҆�a�B�M|� ��{���i�"���w���|�Svv~��2�p����n�c��?�X%���l�ղ��u�,7���U��o*s���*�D�+}�#�?C�Y�~�CcÄ�g���j�p�:gFq��o���X	n����W�n�+=E$�uw7��{��5C��ck�S��n�A��0��5A7i�q�fv����k�>T$��BlTzP�xP�ߴ��&*ۃu,z�����-�[{G�m'>DɅ?t�v'kZ�Z�3���5вh����1|o�(&�:'f��SK:7Z��jb	��/���i�zV��|��\	{�p����΄&�u&�A��e���|�F�}G��Vg*W�a�"�����\V	���i˾6�h����,h��]?��y�}�Ѝ��������˛�	��FZ�!��Vl*I���Ԅ0��[����_y�#�~���7�z���8��z�2}mX2NLF�n��??��
�� �MMN�ޭ����86�����7q"��i{PI
�=��{بg�.Jt����Sݫ�	��Z������T�q.� X�|,��Nvl�X`�2�Lj�ǶQ�0��ftf4O������=R��Q�"�Y'��>r63�Ēd/����G�h��Wy�9R�K�p�4���7c���rU@*���t�O�����2Nm��ɂ�i�����"�I#��0j���(��f�C6>,~�>#�%�����bHe����w�D�5�Tu��,<�F���r�3AZPF%�u+Q���uʿ���Q��*,�n�Ч�|�d�qHE
Ur��È�cS����[��f�+t�_8*�~�<�x���X��$�v�$%m��#�.6�,X��R���:����)5w�_�&i�F������.�:7x��X�~�k^�>��C��X�G�H�z�����x5V>
fALP��m�:T��}
�H��/�����u.'��`;Nx�%���K�X�R|�f~��jˍ:�۾f�ϗ�{�;Y�P�l�%9�1�T�ӝ& ��:�ׁ�AaJ���ou�ؗep����Jg�(��`�oŒf�ȍ��y��*�#��]Ꮄ�.\��~�l�v��d���B�.��#��
�����ɗʟA���������v$��?��T�sx��� *��sf��nq�BۈS�^�Cewh@#�*1�o���ùxcj������A�Όg�*�U�	�~��CYi8CkaY��3"^y>���Řg�՗�´�fd=�B2�F�4K|���.���A(�ؘ���3�i:�i�_��Dr�g�&|_X�gkw��COM���x�N��&汯�[�65��Ga��N$�Z�/��2JX`��
#�`����Ar� ��p#�C�
�Jk�����EL����|,�w:��\k��ޏrN�g;T��]��S5���0�'�� �e��"gX��C���>r�9v=d\u��d�=t�����BC7�MǱ�pm��5����`��y�-�kR�����H��t����z'�7���j�5���A��"=�2ʲ�Aƚ�� ��ڃ�;�_�7�29ϔ���nT]��T�+�鑑�u�Jg\w�����ёգ-�*5�f��`��R�=Q5����k�g�5oq�}B�췃c�F�E ���u�W14�n��p�ǔ��}U��8fB���L�Aft������1�q����3ox|VHZ��
#��Y�@�m�X��}ai}�p>a!�]�v�X��&� o~8�䫦3x�W���`앞��V0�k�iX4Fw�Dkz��fQ�>�S�Ƶ��/O��]����&v~��w��7 �[E�k��cWU��@�r<���r�I�竇	�����޼T��ǭ��cK�u�3�ғ�-�$H������X����V5i=RmZ����Z�,�[A>�2���}�~��Z\M�4�|�<�	��BZ`��)�?`S8BE0���Ѳ����7�0���%I`0�����S���A��NۦS6�?Z{�Ɋ�[���2#Jn�y=�����Y*4�aR��O/���|l�B�ч�+�H+�)jx��A����}M<(�xN�]�/
Ð`���Uhݡ8}�$@����Z���HJ9���@*������&	���筰�ĩr_�B���2���s/@��5'� ��T|�x-5��	E���=�?#�BY;`Tc�Q6� +�83,Z��=8̸��i�o����z`�-���Dҭ�XH���L�p�j��5};�J���(�~�6�pV�/��u~&��o�h������4|���5��A�15��
�ύ���k�쬂�vi��H(�5����b�v"��3� �[��� O3C�r�,��w�W�i����pN��	�@�M|���mH�ABb��)�P�����kǄ����$��� �Rʅ(��G�1L�����~H�Q���ɷ'
��z�K/�YY��@�[��Ҧ�O��8˱�_w�n��t˚�Ǘ �e#'���;$�A�\�VM�٣v��$��]Δ���ɟ����⏤xQ�,��������#��4�b�O�_.�#�c� ��D���O
(��n�`��8�M�-e40qR-҄��pmAS�T΄	�̳7�]{�{���U?U����wvޅ��8�����aR����/r�!1>��{�G�Mp����xX���������k�_�c,$����u>�l^�X
yB*�L����͚�ݺ�Jݤ��. ����>cu��a��JO�MS?��4�!;�Zn�Q<d4��U��xk@�Z����;�{�L:ǳxὧ�����;t����%l��i�J������p3F��p#%+%lR���
Y�	 *R6���kI�Xb�۔
o.��YӋ�ŕ� ��p�р�9���)��ȕ5+�yZ.j��;o`o%�7nt�Aҷh�k��֬	 �&�iv�Q>��݌E)�<�sa�uiD�6�1%���Nh�Լ#���:�QaH�N��=�hR6�('����VU�J���Gț��I1��3���0ׁGo�����e;-B�,��$�����R&���ŭ��ߎ^��fxD�p=�+R��������v/Y�Ʀu,��Ô�S��ý�u
Q�X8,�}����/@���>=�%P=e/n��5���'���s��䡴=P��Q@��s;~9�'��H	���e���d{_�n\����!�Rؓ��O��iƚ�����FS��y�$��B��Ϧ�6P�#�J
#Q�>�����	 �pPΟZ-q~��t-OP�^�v���}:��X����)�BW���bx��L;�#SZaV�D��U�^�۝� -�!�玊��H��X��������O�>
��.�$��ⷩ+rα�<�5�{u� �m�`:�Q>��8�ƹI�¤&r�H�����Y|�vv�������]���Y�-���+L��xN5?��-��'��N兀f~���d��`�=�H�x��"I���q�-ᖭ�H�>X�J����dz�@�{�*��Vȗ\�VbbC�,2��!���BM��]	�/'���{��)lhx�&g��=<�����	[�zȣ��)�]zMW[r^Y�Y�\e.s����H1*�ӤЭ(i�;erܰ�17�ܦ� ��F��]��?���"p 7��p]E! �چ�T�=r����2?���ek��d�I���i�����G	⒒�oW�G^����,��g���0����ͤ[�n��?=4��g�v����t�CkFpX#��1�նv��d��!�as��Y���
��x��5V�� ��~��]��{U�6�m���dw-8��갦�>����CMb����r�+��/$1C�n=�W��81��r�8b�v���3ש󅱾��PL���!>�x/�,K�����Kɇ�a
���gs�Qv���2�J/	�1E���� ��-���$H�(�@9"�}��Y~N�> ,��-���As|%�gRnFG%�&q�v��F�WZ��a&�3�o�(�>e�
�7�CVW�}��r��x��E���K�뱐�G�VV%��s�#�+#�xT�ae�Ռ�ֈd�Mk^���]M�m���B�ƥ8;xwQ_|jЯ�,�AJ4�smG!��ab��X�q��JF��>K�/����e��lqjdM.�?�PCn5��>�%�*��
���r�נ�\�SX��,�o�B_ ܹO��o�,��9���-��P۶�@&M�D��e��{`/F�!E�):���]�h\ �=+h�h�j�F��9�91�"S��Q��� ��\��m͵g�K���i�K��=ؼs{������궧�/�(� �&=O��EZyj�xGv"T�og�������m]ĞMk����h��G����-��P�L��Zg����Ixl��:x�͙P�|m
B���[���G�/����ed���z-W���5,'�x�+��9L%��;�ܦ\F�Ո@��&{�P=�l��GD�/"���x'���6���r^1�<d��j��w����P���z�p˥�]��2����2]��7�O�W��_�J�F��i�� �Y�akks�q��b%�X嚈��hw����甚�nڦɍ�����%N�<�Y���a��hjK:�9Zrl��l}�V�B?�V��W���n�1=�)��?��I�E6 ���#Te�F'�������o��H�B�LY�M�4�Qh�1�n�#b_��l��������X4��Y~�x��mCKsO��N�]Y`�s��;-�!��U!m.�o6��0�5��}~�<�Ԟ��MC������>,G1DH����eB�q�H$�(*�Q׳��P!=̠5K��m.<�������Ytt���GWw���#!%LxFbK�@P'�p5k�饁7�D$�%k4�.�C����]����ĩ	�d�^�z�ˢ1c��ׯ���{�n�5(���z�E��Db}UB����������w�.��崅�
����	���_Rw������*���4]Ms�L�ķJ�]��Ɂ�j��W]=`x@[x�� �"�^N~���J��_���!��h�2��Ve��L�K[�9/+d�$ �4;�E���[GO�߈�5.85��`\ph�6]��2��L��J���h���{7��L��f��O�⁊~��EVn	S�ʽp2>���'II'J��a�w��Z��'j�g�X����6�P-uU�ؑB`��n͕���aZ"��ѣ���03}b<�x�m���|��z1�ʋ���#eK�&��ؤ��
}s�I T����ͺ(#�f���ڎ���ZZ|�R߼0����;��iG;/��b�*�_�#V�ϋT`����ލx�Bruޮa�2�8y�b�FQ�(^UI�$I�g>a�c"���a�8��>�����r��V��:�^w	.�%�}��	*��Y~��G�Q�P�S��d���c����K2x��~�$!�R��J��X��z�Z�\Lg@(���ώ-W�rT"t)�J�O�` '���T�5��µ��ۛ�/c
ث�/Bl�S����v�$Z4g���t�༻y�u�<��o�LrN�]�T����6Eu߰w��1�H�*/���b�������fv*���i��yH�D����(�!	��R�N���'�%��Os�m&WXI�K�)
A���Og񾐉R�㶪��콤p�D�l�R�J�!���U��b)�2a�*�(bǾ��#+L�|O�����q�;f��Qd�ɧS�f�hʢ����:y�)���F��X�� ���wz}�{��'D�CU��bKI�5-�5��㏕Z�$X�\�V����>J��ruY4�	A�m�.����VZ���;E����L�T&�@i�5D�+>�7q]Vð<��rl?�h��/z����E�ͼ|�a�эPMf]�ɤJ�8l5�e�<�TJ~�PTD��֜��
*v�u9cIv;��)�����۱]*`����I�Vfv!�3�����r�h�ҩ&C����%{H0@��D�n�7.���<�H�������n�M��c"�C����8�k!��ɳ)䆰�VKU�xD��{��u��l[�,\�5_����O�z�o�ھ�=wb�&R�~����?^�d�j1�ywWmm�DP�)��Ǉ$�+��bk����P9|� wZv�ѮV+�_V ���N����a����y�E�X�J(p̈́iJ#*��=Ǖ���1u�g�hl9䓖�3����}������������ �u7[�{�$����x�>`�,�u���v5J�"HaI�<p:����M
�ӳM�w��5H���R�#�%���H�3��=&�^�cw�n ݱ�o���-�?��3;�Ƨ���BM��Oh�R�4\LpX �0:����6=UFA'��{�^<�&��n��ݘ�2�8��&E~�s{O���)KD�����iS� ���Z���VJ�]��(3�Rw�H�I�S|����q9a����z�7$�֎�H��v9��7�/qr�]8g��戤
r��*K��F:����3N�,Ŀ})��TWvN���_���ژ�"i�:F�I�sۢ��Q��Lk�2Z��"q�M3"8�'zhD�&\7���������:{Lx]�C7Wc�
��B��{!�vw��LU�p�3�a�r�&EB���#�u���x�+�t嫧�nQæxn��/���nb��.�n�s?��$䀨R��.��`�Q�D�\��Z#�G�}���z��x��n���#����N�Р˷� ����Φ�������%A�#4�ߍ�?mKez�p���+��п�ę��3d���v�h!�ا��;�\(�c�D�N��R����B�}���2u1o7��i}$���8���sF뱌�=0�w�t�����&8��m�����%�}%��|�eIz\���_}�����ĤB�H��3ɛK��u�Y��qљ
�DG����y<	 ����loz{�+� �o�^�lmM~ڌi'�J'[���,��C+�*0u<9XV��~�$�p �B�@?`:��!n*�c��Zo��C$*���	^g��m���t���~¹��s�������c�]��YU O���z�|� d�\ �V�ъ�2�(�8���pkc��l�;X���W�hA*8q���(f���4n��S%�W��Et�%������v����}{U����&�������e��,>�ً���t�-$e8����ڭ3M�B 2̜B�^RO[>�T$�_
 ��3�.�]�s���|B�If�y��H�K�-l������6���c�S���-�VP�6�S�%J`Mbdv��o�{��ܿ9M��]l��ZZ�_����#��̊�`�=�3���E�o��m������)W�)]��=��ȤN�4���gY���8T�E���Eb{��_B���Ж7����u0�]��;�!"�D�^gլ�@�O��,�j:4�LP�[xP���;���H'VT�����3��������(�8��~J� t���
P��J�D55�I����8��!J_50l>NMF���%<���-�
Sb���I>4�I���լ{�b1�z���N0��az����)�}�M�&�,�<2��d=n��SMn�8�p#��͌ߗ��	"$��h��]Ú�O���Sr���O�:�;������5M��|�"_�l�Q�R	h�GDcdJ������O{�[�||�.G
4��z���Zn㳄�~��aV_ݵ��jM�����[Q5�S\N-T�Y��u���h>]�-{ܖ�c��"踚 �Fn�<�R�9��!��V��Ng���[*��:A�ӑ��ӻTW�ہBjΏ>��Ӽ�u��aV}����>W��w�'k}��tf��=����0�G|���A�8x-�����i2W<�4�o]i�(�p;(�`LPY�sX��<��&���Q������i�湧�t�A���2��#;44/+�'����zu2,d�b�ޑ�X]�g8��4O�	oR��4�=���������0���C�߰]1Q��0Vp�K�SP�(ʨ�|��⭏~d����}�5�*V� Iˢ��8������ա��	
����t��!�{��W��5?X$��2���!�C68��t��JK�q���_�A�YC�{l�T�(jD��]����A4�(w���Y�c]?�bU����O@�i���BI�v�\ߟʳ&��״1�����#�K�f����vh6�L5�{7֛M���k�x|������	��0V���ѸN���;qZ ���/m��Z��{+�YIo���.#y�#mP���=Z��ծ�=a^��ehg�O��
z	h��al~4��T�R�B������{�m#�o`�]�N�$�� �d!|��٣����DǮ;������[v�����o�>j�c��?���8���1��>��"8�x+$y�MRWTv��$w>p���p���LupTG�:RO������w��Q�/pH�.`�ӎ%J��7,e���?tK����\�y"���MB҃S��Vڥf�o��_=��}�;ժ��7y����N�Ll\o���	8���Q��Uօ-:����p1n-A�,�O}��ɫj��\���ְ?���6�:�-���|��\}�s͇���ݖ���9Y���N�@�^��C��|n)��[o���-��g�����ק�
�L�k�Y�I�}�}��꧅��C�9��.�#���*�pp�,;�L����te�jY�o�گJ	,i%2��:oq�G���EK���w�w��Rs$�E�����``x���r��{<�b!h��z��`.Xl�%�z���c���V�?�:�c��D�����7/��}�Jf�	�G�#:�}嵾:(�F������-�eCU���|1 ��r��]%PR�� #2L�}�T��_G�L��S
<h�\a�)l� AQg��� �{)��C�nrl�.%W~p����x=���0��a�n�����_n) �c2�V8ʕ?4
��w�l�ݒe��K��� �N�رi�����o5Kd��-�Q�G�0�A|���ݍ�*ڦ����܈���+��l ���@8�l�hĎ-"��?�|�*�� �������k���u��qI�M;n41-M=Ǒ��_�)/�����q��_���Xd�N�jj�58#w%�w�4�D��.:mЇ�Ӝ�-~NJ�\��F1�N�VP�����UսQ�R>H���	(H�Ʊ_���p��(�8���g���.�%��
0�Լ�$`�1���b����K=�F�?�ՎvM3%�?����=̰�x[��v�*�H��}c�lOJ�sF�ׯ�a&�Y��V7��ن ���
��2�/����$8>���I���5���+���;R�@}���t��9D_�гCX�<�%�G��iU��.���Ɍ�[���#�<23��2'��נ{j>2�J.���36l%�ĳ��{?�sN"�	`� �2�6y�a�d�H��T����Ms��񎈫�-�5F��nI8��e!��ph����BNO���D��kzu���e��H��p�Ɍ4��m�+,��kU�_�M���.�ZH����^�V+�=�W�h�xOgM�K�RH��G`?�$��(n-9�-���z��<�� �<�	ƪ!eT�F ������#�#��16��L�z/W���g�]*\�n?�VG'uqF�a����%!3�Ҏ�����pt)����!=Z�$��ҹL��;T�Wc�2�g[���0Ko{�8�\�x����0m�(A��߷J骜̬R.�\�0��7�GPL��d���5f���W�J�zM!v�Y�/V�^1o���!�3n�F�ϳ�F&-GO����J��j�;����姰�q�ٲg ^lXs֬y����g�!�1�����%�����-�r�Sӽ\g���a�F��g���Mg�Y,:Џ���Q��:g"3��x2I 
q��M�������@��c'��L�C�~L��L�A����N�u�����%�,6L��7$%2	�*Y���fT�F&���<F�G��r�y���C�E)�RllO�69��f(�;?��T'@SɏܞZ��H���]®�)y�W<���{�5lXyMO� �g&�����t����E?��ܴ��&��>[�0^�5{�x��b0׏�9o�KPɻL�G"*�-�8דӱEVh>V� =!�4����8p)�>υ&`҇�[jCQ�L��&��̪�q[dx�&�y%e�N�d�TB�R����>�yw����<�+�ɹ�sD�����z��A�S�ʂ	
�q�V|�W���	g�o�C9̦�%����Gi,��j���rC����L�V����R��@y%_`S�r/��|���&U"�W��
2�U#��=�`���\�*@g��UnB"J.ۈ�>�h9伱��G]B��g�Q�Y��)�8�������Wuu����XVR�liS/ś�+�]��S�Bl�ߦ��鞾��J��vZ��b���L�r&�QP(v��-f�
j�OI��z���A FD:�����w���_}?��+�U�L;� 2����`~S�B��!`���B���	L@H�C�,侤�2Y���N���8z>� �-Kp4<̲]1yB�)��&��H�@�S�i��50RZ����(�c��Am�����ȼ��e�
@䰯q��!��8�#��lV^�f�m�M0#�Gw�,[���-��9{^eş3D����s�f�Gm��1|���x�i�YQ�~X�����>LmE㉕�D�6b�c�r���$ݮ��U��PG�'�j�~�?����Q1c�}4������|�_6i�'��� Z1z��iQt�n�&*�K�ԙg�M�\�w��b4E�b��Tg7CU�D;��� K����.�%	6�_P$�K�c=ItA>2enRu͗mN�����@���X?���$}� ٫�!w�ʿ'jz\�	%�l
/ڞ�N���4�~w˴�7�?.JAL��2���!i�S�,���:^	e�7���1���U���F���.
#��r��.��M���]N���3N���@�Ar�>;�; �T��-P�D2�Th�M�V/�[�>�����x��П���qY�0���L���\.EĀ)>I?��G/����˳�U��� 7`4e�cD�='�:8XfSX��e�M~=G��'���EF;R�;�L< f��y��c�_L��qpЌ�����J���\N�����K�[�:��~�Η헒�B�{�!��:��XL�ѐ�e;��7����U/���np�6j���-P<�&��۔�x�(�c�k;����eV௽�q93�{�]�\��ᝈ�7x�5��?.���z?GK��_�?pm�˜b���YYY}�	+�ٛ�˻~C��A��$NVI2+�CI��ʮ ���Q%�$߃����8�X8L�AwYϻ�_�Ah��/�v�m��D�yx�z��?��m��16L#�|+�;{ Y՘G���C�4^�i�I5��H�j��
Ew�.���u�\�K���+��[ii8K1��1��;�ᙒ �Ӎ��apW�l��ד޴�>䌒�/����F�(kܝ�m<�0s\��:ud���t�r�54VA-����X�Y^ou'�IB��dW�)/sϧi����DI�8��4WD4:��jN�!y,�O E��5x��k���gX��=��xl��&�U���}��O��xE��0W_2�o��\�>yg^�J��sZ�g���
��o+M��9�U�`V��`=*M��י�j$-���F	��O��~�^8�7���Y�vӜ�]*� ����#�T8Q�::�(=�t�j���`;-%��(����W>�Vj���d�?�np���������&�4�h2������V�B�\���d����x���daߏn�ʫ�������~�ݾK���Zͤd����`֪_}�� ��<�V<���#3�7���2�"ˆ�c����j���c�V-s����W<'xD���G�"�^Tݧz ��f>y�' 1uw��
x�[��#�9����{(��ց�}��� �[R���IY�2��5
u�	9HŜBx�ٽ!�[+��h�*R��a̧cT���0vs5�q�hR� Mh�+�>�����i�y+��m��E��D�)�X���q�i��?���F�/�x����\s�8w� ��{���]�[K��c"�C�4x��%�/�x�-����N����P��tz�r������X�N�>@s
ٺSs��SjChFV	ic|��;�,�͎�]�
 Mڀ�R�#2���&��"��(�JX����0�@uu�-�R��HN��'I�N���b��4ZY�]�sn�(���D�q�W��3��J�A��?�
w� '��l.opx!oY{��H`����`�������RdDv\��}e,�`��tu��b�Xq}D�*Z4��G��>�@,@��>ֵef_Å��b��RQ��1�ӫ��	�O��YRQ��}0��4�l�D�M<rq��&�FѷpJ �]�hԭ
�d�a���q�@��=XUjd*I�1�;�,��B�ط�腽kH7��ĥUu.�x`o!Eu��8��Sp�W�UkC+�H㰷+1�}�SIQ����#|_c�|{���d��\���>�T���q�g�/^gP��9���%|Jy��W]�<Uךca�7��z��w
/�\g����H6Z��h0��
]�Z�RA�%[ (zn��a�pؿłp蒐 R]�ˑd���5r����m��·,/66.��t:�7�����JE��Wv�i��=��T3�3%%�n��0KƦ2��b!-+
�����"��0������ec��;�X�%����5�t$��:�����9=X�`����K�)�IWz�����$�D�ke4�j[2���V�jƾ�h���ֵ�!]�7 �Oo���:��Wk���$ǵ��*�N.Qr5��<p�}���~Ӎ�GY��~�@x9�j�����#DlL�n�	�PI�Fm*�H�M>����-�$��K����[�C����Z׋ڱŁ�������p/�I�M󗅿��Y��Y8N����Eǳ��e*̗��:3d��y�����'ݑ:˭G�$�V{>?@�eژ�����B�רG-�����N5���dޖ�4���b�hq��&oOAp\���&�~�NB��۾�4��wn`���<h5�Sb[+$��к���Lx0�P9�����k�����^���0�[�q���b�c'��uc@	{�Y�����v��>A�������5�p؄�z�O�h�;��Ź�%�S^����=e�/*� �3�KŽ��._���L�W���'$��1P��E�z����Oڶ�_�Ҡ^!g��ɣ|�\Cב�ݙ�s�p�\��k[�I1�uֹ� n�94����zTi}�l2����^�@��	�����`̌��߸*he?X&�P�r����
O.�V����-�8��$���A�Ns3ą.�G��/��|��t��hA$Rհ6N�T��E��f���x�^B='��7e���dZǼ/���'.'L+n��c>����{�]	��C<\��:�H1O/fYƃ&>��$4G��N��Pҏ�� Yx�i2��'���։�k�}��<���}|�� �{(��^_=�	<���Ȩ�5�4W=�X艴��\�_�C.��/�8��_���lg��s�
�ޚ��)���������ߝp�~$%YtrP��lC�E��ɳ�� %4��R0]Z!x��lXSg�<N�A�V%�� "�M:
�j�!�m��{b n�+܂1z��ب6���.��-r�KRBP/�����J�����S�ا�n,�������|��K�B��=� ltn�=�xкȫ��%&r�㡘f�.8	1�|�[���p��a�����.�e Eh�o��ˁؿ�UuE<���L$E���j٪;
ެφF��㑠Z�?����f��r�_N�@ً�FY�5L�!"���#��_ ���0��Ƣ�U|����v̶.�K�[����v����Q����F\F��NE�*873�P 뛑��4����MH)��X��.��J���Ǐ���7�W�LQ���gC��i�[����KVԛ�!j<ϴ[������
a.��KbS��д���� |H*��*�r��g��2��
=A� �!���,��l�"��?pj8��)3b��D*�H�^E�An��W��}�r�J��h�(_�^��ª��޾ҙ�zo�F�߽amt�DV'.џ#�=�$8��LE- �N�S��J�,��E��5���9-��Y�J�σx �<5h{:��l3Do·q����6�P4��e�xm���"���XRvM[Ȝ]`�E�C��s=T����z��x�r�ib���UL�����2��>��+,�G�޻�ܶ2;����&��!N��A��T�_%h,E��`_���sm���MÔ��"�4�,\S�	��ز�X�d<�&�v]���Q���H^	�ut�0`Z�+mAv�D�qwI�Ӏ�C@~��Ʌ-MT.���J� ����u郠�m��絑d�xae��nl5��Bv:h�m�:�੆���F�_h�,ӊpPGbS��I�����Qp�R�F��@Ȼ�������Lɥ��(�fg�n��f�T2n3N�W�$����Մ���:q>r�(Ĕ���O��?�oaɕ<�Qat#������ٲ����������>���� �NΙuN��Ҙ��4�9,��7���n��0�Pi��@�y uC�O���9�gG���=a�OI5�"�r���YS�����GsIy��ʍo �?�F�F��$��n�v�1`)1�^Cy'�{��dWñ���.K�鸪zI��^��:��,߸�*Y�D��H�yǂh����M��'1LO+l�Y�_�W����D��pK%�/�yH��*|��i�R^;�*���~��Nоܻ��uNS���
�s>q����!�|����Hݫ���s�ʼ����0�_��M�xX&@�n���~�0S����ǯ���d�;�t���7��M�M�wo��*�u鷗�;��-�����S�@N�����j_�6n����������#�{���S�#%u��R����:�٘dQtV�Q
G�jA�w�'e�-៝0��<��&B�����@����:ќ�:��j�4�:+qD�#__-��nd�ê�9_z�Kg� ���O:SX�L�J��M.ט�/�8X�%_�r%׺g��,k����f��<�4�����I�����;��� z�Ey��9�qb�#�5܁~EQZ���|O���GhI�(��@�
���<4y1�ۛ�LW��T�~�{)t�c�[J�;)x[j������`]��`օ$�jw�������<Fj�58:��� ��W4o�\;����D��:�MVZY���M�c�j����� Q��Ђ�JA$>r.Hs�����'��0�Լ)�-�v� 3*��Ҳ��Т���������4�j�{	�Qs��ӗ�L��p.n�klX�A-935k�e�H�K3+��F���H`kܪ�CvˍŒ�ϰf�W�Ӟ���4!�G��PtV�JB^���*{M�w)��#�~��WH)M=+AެІ�˲���?vϛ� �!��wo�^�
��������]���V�d	�;��U9R�����T���Yʞ�]uZ�<��>�n���s��j��˦����jDP8�P�z`�kJ��C��~3����`�EZtC,�<L��%��a�����-\��}�#_����������,.+p�m&�都ۚ�'�l*B��_�N�UZ���d�4�����I����]��ҥ	S:J�s�a �� Ņ�<f|fuE����d�iE�y��Kl"�
�ֱ�ؤ[��LY8r0 ��������7�i���A�� b�  �@�b|='ץ,N7��W�Gf�[�-g�z���- ���)��'3>u�&���n�%~�kZ�>A䗘�d�Q$.
��Ŵ�tK���l�!͘=��H\�:#�L��~.{�mf˧�#\�.|�d�
ўM�B�Ϳ_'B�}A�gm�괟?�Ķ�x(rD./�<M�P�1��55OVA"�����Ft�"�הƛ�%�&��AUM�'GQ*�m��&���c��;M��L�M@��{h�!ma�z��JX�z;���:�*�R{��P���n�ߝb4ד*vt�i�w��*���],|��̬�)MB��_\����#��:���ƣW�D�NdS|-�'%ȣ8S�ſ�����݋fiU�*���9"p�0=�T��>3A-B�>��\���Ǫ�}���3N2�L������,	V�xU��\�B�]R��è��ۧtr�C�����<���څ���$����k��P�ǭʯ�ЎO����:k�ȱ&�=Zz�Ew��j��]h`������>�9�L'�k0��b�H�5Q;�E�$n���k��]��nG����{�]z:+5]"H(sa�� rb�R�h��s){�-�گ�=���a��u���S�=������z���Yv�a�ؽJC�ٰ���(G1��
ܟ��������� �Ha�j�<>��#�������B�%p?��{��,����wS�J9�:��&�l�����~N��YSB�m=5KK�,y`���7���"�L��,��4���!�4V&CV˫�ވ���+���D�)��w����%RM�뭐2Pb�p����{�2�vs���qW~/cY���tt�X*3���p�W��L��=V�B���R�=�H�coO�'N3�"㭀^6�:;J�Mj�4��G��	�^\�ؾSq֗;����c��Y����a�G�8�@,����U��W��*=���Dn�~x���*]������I��������^&�d��V��:�l��1	7;��N���9��s(:;��(صFw��`w-�����NwU�a
s�}.bq��� �6�b��)Ԍ���H�e[�af	^��j*\� s��ya��vE�ORX�D�V�y���M�.�['���݃5�u*E8Ԥ��@L7뮦u��>���ہ�&�C����6P:o�n}��r; ���F�s�`G@c����f�l��r:9�,iI�pya�q����V��I]���(?Lb�*��N8\m�M�]p�n{kނ�U:�F_�@Z?<���\w�9#�a�J�:�4ҵO�zEU��?5MTc���Z_۔��&_݈��k���j��~o������'~,Q�6��u&G�=�D�[���e�� ְ�T`���|/�r0/�"Z�Ǎc�[�.��k��ر����6��'4A��
^?^t��I��o��4t�l��
�k���1[�<��p�DgX���uГ�*��
~��x8�aÁ7��m�p���%�=�$Lv�ãɮS`��/x�j� S[��|V�g'QR��l����\�,c�U�3N��}������/S���N-)V�ۇ�@�p	�m����s:ftS���ʢ<���;>$a��Ybv3�Y���W�
Ec��1<��Ж<}$�
6\-h�?=p�`ByM�ɱ*�f�qR�b86v�,�0�/�j�m1^�2�!�&���>�� .F%�Xz�����H#�+��[\����b����*�c���u^��eޯ��I��S��a���Me��F��$O� t��rz�O&������[�m�O���>o�����-J�����k���'���O��͹�1e�-� ����$md���G����^�,+(�"����dZ������M���z\4���xF�F�/�i��۔�������L\+>��K�ě^� �xB@�Q��s1�1�2X�>~Y!�>�����lٚn����hN��Nq��3��J����>+ް�����uOO�Hh#��ATm�D��Y�Ջ2��`Pn�p�hkKD,�f�ScE���D�9�Ibل����D��Y���M��>fI�j0��c�%^�S����c���ܽbD�;�	����=b�~taO��j[�P������50���/�\��J�OK���R3"����5㒙�5�O��aPt@�1߀<���HO��ju��5��P�@�l��%k09y����7�;V�L�������J=���2XtY��^�p`/O��/��M�8����$��fJ��������?��P���A��]kUĉ��n��ZH.)���<���~DNFШ{��ݺ��ݷR��q���3�[:8?�لm��R{l���J�J�"�g�h)~�x���>C�����%��C��MK�<`Z�B�J�"W�=�����%�~ ��s��aAQc2EEt�.��R#"?E!�fA��~�?�}CE���I��!"P3,��:��8�6;2Huw���b�5Ѝ�1�"=5�~E�^����	��8e�,k�$�[r���=X	X}�Y`z¨�wVyF���׋ 9]�NL���7��E���ā_mU\ cr�10�*9|n���(&��[�(�De��{�)���?ʰ_��s4�C;Zm'�����������@�s	__�!�LA�:�z®�x�_ [�"jeБ`%��,�(��U�X�HJ,�P��?Z)nG�LS_}#]xx��#2"���.=G�#+/n�NK�̇�3jh�C�Dhj�@�