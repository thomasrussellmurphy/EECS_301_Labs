��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>b��z�P��`S*���mX
�Y/��j�a�tE�+rސdc�x	���JmB@w�`�Ȁ���`���)�l��� �d!V����g�[��2&�3B��D��Ղ&zG�Cy�䰿�sˇ��.���ą�u8��2t �7�^/���|z6�8C��'���a�V������,?'�s�Z�i�ju���(7Q�81C����i6
��T7�}P~���T�ݫa9�4�V�\���( ��._#�z�7�0�/���CT�wĖ<�J��� ��9�z4��
:4׷c(�~���!]�嚕�E�@D�S�w�f�}�X%���w�mx�YY�7����Ei�ݝ�I��C��0l���{���'�h�(�������*Em�ާ����#{?�d!*ts�ϯ��C�Ǘ�'$��}�i�t��W�R_lG����:h9��y�_����T�q�řqju��bAۀx�;���b��t��S!�ǎ`�I��l8�W��P]fs�����I�!OݝS?��P/hB��BLh�c)�;H�|-�n^�����]u	C/`I�x'�n�m�y	b� J��J��{�����p7�%����0���܏e���6�Z�Ö_�������q<-���Q�Y�����
#_Ҋ��:���N��S�I���a�������ow��v:b	 Mn���"<k��І��'f��G�9C��6�at~�3�O�����y^nX�پ�i��\��3K�Qǲ��j�ş\���5�F�U)%ѣ0����^&=��N�8cϵ���鈁�-��rl�%&3�t����~T�`�䋓ԗd��lq��VI�"�Zy�_ee��~$����Vk`��lM���)�&�F^[��cɳ��yx�c��B��-ϥo9�9F;s?@k��S������Z��s	P���gQj?�� ����W܈���'��W��7�{���CN�:#JV�J�lh��j���*f5�j�q��'��� �B[��]{K��{9�*S}&���������q�R�a# �95��a$-�Q`e�Ͷ�'$��m!tXk7d���-�LK�ϫMX�1ҭ�q����uI6�So����`l����r�NO���
�>�/}e"�D��1��Z�$�>�6#	��bgqX�J̘m�2�j$�]s�~��R��������<l�Y�����}��H�K@�;T����si�����x6���'
K�9o\����3W��'��z��	n/7P͢F����]	��*U�'���N7��>�Q��'�O��C���Ҥ"�M<�>g��-���7i�)C��?�6�w�Y�)�8|}�t�$�@(����D[V)P�n���������8Wf���T1��(��Y"���08�Y��� i�c 7�Q{א*J���^��5�	����Qe��҇;�@���B9[�A/ҧ�GdXq�Lo�_��	?�����	<�wn�EY��𠌹'UC���|��RV�I�^ o��:��Gg�X9C���p+j�ARS>��هmʇU<h��7�,�-����]���B�m��-{f�tZ�X��| }q�����g�G
QO�oYUO�*�D�P��M+K��+,%A�lq7%ػ���I�QH�w}���n)�[��߮����H�;�1�0*��۶r�$9h}Ѩ�fѲ�?\x8f�A����.�������\%ެ#8멶�7�֠rgg��nw�M�H�
'vA�z l����H]b���N�ǿ��:Ŭb;�`9�T0��Hߟ�w^}E=�U�Ɔe�v�7�+Uo��L��b�^�a�_=�={�q�21I����?��^�/t;��Vt(�l*[4��L�u� >8����u�P[��y�v]���Z�E�bz�TJ�'�c�;�V��*J}�ۅ���'�D�:�����f��0�{Q8�V���vrvI ��R�;�H�]o�>q�^�S��rB�ۆ�*
�G��TK�m��W<�x����|�۾\� �!��`�Rb,E�&�i�-D1
��l��]��w�z���25^���դ<Ba�.;�k���Y����Ө�&X�%��d�Is�P�$:�3 ܉�c�cO���*6hVp-9H@�L� �uia�l��D�[ ��C�!�T|\�L��ET��%���<O,ٞR�r
�]��9�ϘJ���R�㑠-�!�����)T�N�P0�=>��fq$^���e��� xZj�����<f;@�F���G��&,�b>��)�z�@.���:Neduܵ;�XDv	��֘r����m����}ǭ2Y��|�Eay��|��>.6Zn�����3M�V"�����qd\�4sJ�j�����}D��f�t��9�k�Di��bv�gB<.ŉ���Y46Ў΁�u�j�/�����.�G1���6A��}ba��(:��6V�+V���*�����q�s����$a�!�s��"z�Vh#st���ԓ�	��~�F��u����R n��̑s�cTV2?�[�8�����0���#�k�(�k]�AZ��E�0۞��5�\>g����̌�*������}v.������7�3��VZ��}��&k�fP{Y�=%��$��n���%�%\lG|�'�u�3��>sbY2����&��B�0�}ecű��x�ƺ�w5�T�� �#�&�1 ��}�]��;$U�S���z;mJTVj�yy�~�&�I�܈��-9X4lD�c+M��Ii���[ھ@�z�&�픷H��Z�P-a�ex_�o�x�A�gLX�cքRFOu��^NG��z����c]r�N5yz��/t7�j�g�ɵ	Ɣ!�}Y཮��d���xP�����/��Z���P��%?,�{@|�1�%S�+\v���t�G�d$撥đ������J��VR�*1��O&sm��4��1(�M���<����n�Bf'7Z��õ�5�ZR�e|� Ԉ��}ˈ�:�:���Amz��-Ѷ�9�aI��{I �!�駻S�N�_�1���<��B*����Pt�H<bw�P�H�Ocjz`P�iRy?��cu,Ò�7�X��E�����]{]�\����>`�Vu����g�\�7/- �@7��7�'�>܅���2�YΨ���*ߋ5M�ǹܚ�7+�+!i����&wI�e{M'K�Tw�,F 3��"�ww�i�����i3�0d���^��5�������=BP�+���yfU�U�B�j(e;�g���%��C8	TN��$��[3��W�nd��7\P�ޯ��1,�#;:��- #r�Z��w ��RAm����c���^<!9���yn���~��۩�)���)W�*Q`����V,� ���4�d]�i�/C:ʰ��N� ��f,I�������c\�.����B���콟���q~�#�;���r�~��8�`��g>#1|�l�*N��pvY�Z1J�-���L�$�z�E�{
�v�{�7�)'�&I�A�V��j�%0�!A����d��N=�r��j�evB�e�L)�t�[ᦈ��������ᕱ�WM��a�8]���G��Rz28.xF^S���5_�@i	���d������Ǣ��p��<�:���\���4&��5�y��#<�E6��	qz����;���x�P9��Q͇֓Ci���"&��p�/��tD��'F��	�*U� o��fB$�
�@d�e�O� ��M����ԁZ\�m`B����+Ė�NڔB*��jD@�Y�)�fUme۞�_��Rh5[`�x�r�>�]hH��IoO��*y�K�a�-H%��:�dM�����!f�G���]v�>-��z���7(�a	@��6~E����B@Q�ā���Y�S-�O��="��B/S���:��w��\?щ����N��y����f7���ԩ�Pj�n�gڤ�4Ž����=ۜ{� ��y�xt:/�o�h�Cw���3�x9�N���>C��C��b1�й`�}v��˛'凶K���jK6N9֣��!��-���:��m�����V�k!��M�Q"�޴_g� EH�>pe�pyU;urW��!�>���H�m~a��ܻ�R��|f][�10pH�)0���G�6҆������0?�T��D�dh�;����yn!�p��z�-w��# `�>q6�+F�*!"8uܔ��� gf������*;�&����a����،d6t�;-�ku���Y+Iu�ѶΈ�x��2�'�X���/j5��vg��rb
�!�~au�Ѹ�TV7>�l��'��'�%p�?Dq� �h>ڢ��\\�R����9�?�b�1��H���x���9A&�i��x�]ٹh~G��J��C��&qM��̞i޻�"�]��5M8�_��D�!�����\�J`�%�<��(�FMw����Ce�u�-���(��A�YX��%:;.�%�k����]++�=����#È�tx�c�:U=+����o�M�b�ʒ���'�<k���h��}�vy�Ln�¦�����*�~��M��^|^��7�Ι͚Ph�i��Z橍Y�]I�Q��أ�{��T�C>����u#v��$�yzΆ�L����v+�5�<�t���{��Q�w��b%�[����)4}�|��QN� �Z!�sq\$9���/.��$�=�vgs�-'j�]�-��`��K�m�q�� r�tWA��^k�;�c���Ua��@$v(�Jgsۡ���H�=JeἬ޻bNһ��"�����꿨�f�XM���td��?���U��b��9f��R����@��a5���t�:��]q)&t��ܩ�"���7�V�W�0F��q*l��Vϯ�k���/��j�fREG�k#�Nc_�*౹��lz"�ezA���1ڠ��q����P�R�5��5:�)�p��?�����\9����i��,	��M��K��&n96H}ϡ�! �`�ja��IZ���SF�6�=O���85^Y�Y\�Vý�|e���Y���O�3X���%|>�yO@�`�#o���#��M���_�'�|F��1�ӛ�%2��`yea�ÏObR:���
����|�����9{�G���ŷg�_#*�
(C�0D�v����褭��� q�L���������7y��Gyh�v��x�%G�!oF��+�O�UM��bI?�a;7��E����%��l�0������dq���ɛ�tN�����M�������S�Q?�+>���sT�f�a����3��Z$WNw�J����"{N�j�ߍS��_���k���f�M�t3�x9/��_|�d g׊�7H�ǳJ���� z�n�|]#�r!�� 1pH?z�U�sO;�1�䏚w��c�AՎ�V���y�|u�]���1O]�y/Ei��d���sG����a�@�X?rp�?'�27�qE��B�И93��\��F'Εxo��6'�3f׮`w�V*l<�
T���2_�_�����x�N�l'��p�����胖�JK�:����-w�>bh�k����|jp�|��X��i������k��-*�徻�N��˸AY5��1��0�I�/70�[t"��͍}Vf2�*[�D��qϿ��d??=l�o��k#q�����]�@N�j�Z���!���䋎�����Q���O~�ҝ�n:�l"ì�hg����3�������l������	�N(���7�����* X�:�8�a�Xt0���充����T�4ft��5]�N�(Ĺ�DŸ4�U{P[�fy�m�)_�Y"kib�Ð���,��@\��qHB�7�3n{v�=��4yJ���1:	�S"��V@!-ϥ�5�NZuX��� yė}���˯LB���7fV���߄3�س^9�o�A�v�����ɹL���$ܫ�rͮ���y�vv�(�
1�����6�%T�y4EҐ�{��Vt��C���n�iB�t���_��w8�����z��dd����.&T�3� ?:,�'>�`P@�Q��v~a0W� m��6#�!�:/3�X	��������/�|�Q�������h���o}IV��"�¨��d��f����m��צz�cu�rV�8��`H�~���U���Y�[��?�ݾ�&�~`�u^����|Z�we�Wp����`�T�&��C�Z�G�V���Ȭ�8&�\��񱒚�)�0�>醂���x� C"����7�u5Z��&6�~�u�$j���Q����@Α��R^��"_[�v�7,�����)w0�$�0)�$�6P����tP��7��Ѭ���zr�[��\�:kr%���.V��c��2w��[|p0ƞo1GQ׻������+A<ӣ+���K�WuV�nc��)�Ӆs�F�̠od�I�'�Y��;x(��eV����η�