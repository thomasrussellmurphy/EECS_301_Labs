��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\���V�fnvx��ÍG_;�ȅe�~�>���9�>��Y;�0GT��}��E0F�_�o�Hւ�_K��PW���yȮ���gR�U${]N薡�6J��*C.�>��y�%�>�w�7L*�m�	@#�j�(3��-�~�Z��.�n<(�ȗh������G�� C���e,��ǐ���$�p��^>��%@��X0���lO)�Y�[�{�8��C,���xgR��t��G)W3b"�������$��F�ۥ��llDV�j$J�nR�����C����}f���J�w�(е�3b6��@�Jk�t����H��!���f5����>`����8'�d�ʎݮ��Yh����v��̬���y��3^�E[�K-�2IHY8�|�)�Tgk��7൰N���m͋1n/�:�:�h�ч������}���ŮH�~=A��R]l��}��B 
SWD��J����8vC ���G9�a���?��6�<��u�Ы����/v��k�n��$/R;�ǪP� 1C]&^�<��V�l*�,��ir��,�jP7+����y����=lxlY�QGZ.����c�}�N��0S��}�Mg��Ő���5XƉ=�oA
<cIX�ҷ�Qo��9NU& 1�K���<H����F��e��	��\����9g�[�pn	W��;��	_�;�f_�7�xvLn��{�N&�&zS����/Zm(�{�@d�/�m�&��!FHu�Bغ��Yx <ll^��k�YI�s�)�&eۤ�ިm��UKF��{�/jL5���* %��Dno+��݇/Ӕˉ������,֯%9;h-�H��y�R�v�;jGƀ!�Kb�yCU��O1X��8�

�mK,�;9���BI�
��8�9M��a)X�����YX����$ϒ::�1%fD1�e��Z�i���a�\�[�D����Z��#[,!f@Ӿ�b����8��}�ꋚ�qq!&|uW�o�0fY�����F�-��W����&.���(h
5�ei���>��Ϋ�cܥ1Ŷ9��V��g�!A�?��������c��'�CL�X6'��ۃƽ����=yzM���w�8�.��\q��B^��f;�j����{e6����v:��٤M&*�Dx�����fY鬚<h3�@��H�YS��v[˴�Ջ�L���=u7�4% g�0�%B�7�w���@
ೝR/*tU`��(�K��?�.���?���0�T�%�|�Nʽ�aDk�P��`�6w� ׹������*�dz���#��^����U�,�S��);�L��@	�b��9�"Zya֡�����¹��cى	f���Ĳ��rՁ�R�����n��1=���������&�s��Yz�!�w�}�.�J
X !;Jc���)E��҄�R�·�g�U2��'�[ؓ��9#�I�06�,o��[Cp$����Q��\��:�x	����]J2�<-�y|�����m;A\�"f�,�ņ���3qEF��3����uup�y�#�
8��J_�]��P=��1�m  �]����B��P�6a��ZuC��AU�S�8��<���w���#0���jRL�"�YT+6a~|M���&���Jթ���D=r頉`A	����@ӭ�|�~��Ub��&���|��]
>���Q{��|D���m�<���!���5Cn��Ei����P��4�9W�ϝ5�)V⏼4���@��Ï9�)cTCU@b�T�͍��p��t�\r ����q�,��RT�q;z\�	���+�����(RǶ��8�dbLN��v���T����o�ىZ����]�&�F��p*K�}�8ʘq�e@{"��>�Quw��M�K��m�Ht?Ҵ�z���nd���7$�-)S����Lp�}
3Ks��\�\�r���>���<ɝ�1�����I�ij5_��y��ݓ�/���Sr��0�{V+�-ƶ҇#�Hq�f�za��K���9���^����!��pN&Y�h�vތK-�j���B&��7��H�֭(��x?wX�$��m� ���Zw�QlO�E\��ʍ*�|
Ho�U��ΧnQh��H7W ���R�mQ�+t�R�O���.T�`�6d��6��M�t��Ԏ9���s��J�wo�˅��ֆU<���s=�AM�3�,`�!r�{j�vC(�%;E��*�;8�5�=���|��rY��o��/��������<@:-��0ޣ.��خ6M �-�#�8~&�
S��I�~�]<��a�d�G@��"����7��]s@N��Y�:�?�.(S���2-�	b�3��$�o)N�W"8a]O|Hw`ñ9��\��;��a�M�b{FK^����t8�`�я��a,*ͯe5����h�u0y�ɸ$<�qƬ��f*����lmh0�ו�Af �ut�V����8R`��-M�;kJI�F�e�Jv�z�=�PbR�s@rח�;���!)���ܴs��I<�0K�H}ͷ�Q+�yte�v�
��zM�N%�����w���o �h���K@t�8�P�e��N��'�HS�T�-=}��ٴ�j5�H�w_��:� ��/��z~�f����z��P���J'�Y�F���w $�IE���`q��w�h�8�ek��]���O�ė���r�վ'��7�m.��%u�{�y�LX��c���h�o 2>�Y��q���a�q�����f�Rwہ
���H�T��l��;��[o���)��-�N�M	Q�E�W��w�Ya�I��?�L��z��R8�&��G ���@�k>lf�>�����3�=R��A�
��[~]O�1n�R��������*���ޔ� y��bLrp�T
[�(��}o3�P�.��I��L��~�j��xg������'1�:~d����!�z+K�<��iˋ��M�

�y��vg-�
TO���Cb���U����5�l$W(t������<�f:��ZH`���W�n&�4� Ɍ(��&>�-_���*g�<�&�����8q���'�.���(��!?}U�/r]s10�p�\ha=�����ѷkɸ!v�Po�[�f$R�~����� y�qQ��l �0�e����Q�W@2%��z���/)�5T�Ց�� ����k��4�X+Y�������XL~��#{H�ɰ%ǞƱ��Wք��./��� � �	xB�1���վ���/_�}�kB�`k�ύ�Ό�Ш��hebW��)��ik�ŘZ���HD���s�T"�k_�I�U'�-i�YJ�w?��Q|�d]�=#�p�D�+��wJ�粱C�s�wD&F��̼I2�p�T�� 14Ƚ�Y<�r�z��o���i�r�\�o���Ə���%�������]���0V���7��q�������%�E�t�A����ҚFp�)<��ßn�C/�Y�?B������$. _����kì�Ko)VB�BB�-~)�E�q�5Z߁��V��(�uo��u+����]���J�v5ԫ��8?P�П�mm2�kZٔf�m�Vꤱ��Vv���Q�ݕ�<Ukkz��_^���:�ǹ�z��sA����Q0T�2���z����a�&��TU�Z��=-r��,�����Ѭ�"��R�U�)�F�'�d�-8��R#ƌB���çI���KPs��E��L9�nX��w������U�-�ր�}T�����:U1�'m�fi�]�~�V�	���22�V��8�q!�P�C�B,j��ھ������C~ly<�o�~p�Y�uZ�-��9� ~/���D����(A�ğ�<�:!�z*�Fs���ָ�'����
T�r��C��%���
'��	g3o���L�
���U������{X���+�B��`3�"�òY����m^Z���v�Ao��o��7S0*��&�H��1��/m����<T?s��1�7��o!ݤ2&����t�HsԶݐ��|��2�9����'�3�� ��T�:(��)�-���*¸�u�������+�s\"���<��
�'�(�
�u��O�IeFk5HoG7�֒l�$��`Эph����׸j\e��f�	kt����X��s��,)�
M^��ST>4|��6ٺ�UCG�C�>���UH|ߟ���F̑(߃ό,����;~�Zˑn9�XN��{�L���NyyF����JdB�^KD+��x�W���;iD����;���IZ�^��E���w��Zv�譾�=<5�*&3�o�q����7Z��<)#O�%�@5��!�tѨ����l!H�[A�9޻�J��Mw����!���f&c4<�n������_0�(^�2�FJ�
�ȷ
S����	����|�@Q(��� %�L��J���~j�2k|�K� ���*���bbf�ǁ�ǽ�j�Z�i��5B�k~1��$ܖ>A
�\��*��7]��uݏ�3�]�*��=�~Js��$<cl�h89F2W����+�r��X��� 6��5����P����ꖊ��Q���E��e&Y��!��x���6�FU{�R�O�Jh�g�����b����h�3���0U@��qN1�E�bv�Uk��dw����Y���#�<q;��}0flT4	!{u�nA$7�,�C�"X=>�Ý*;��NXm,�(=��J�	��b�� c��pT��bp���C$6�'R/r��^�Hk�D��S�J�5e3g�I�а,��t��#q��t��Y���ŗE3��a���i��$̧C��?Y��L�`QD^Q�O�9W_��jliT�:�l��B��y�~�Iߙ_]����ݪ�e��G<�ٔ�x}Yº��a��JF��[�h��6��7��d��_�A2��B����+�y\�0;� L c�1N�65���A Ǿ�������1J�h�+��n��?w���t1����^6C"x��-/�|n��d�yjv���	%��)��_"�01 M����������0���!"}������'��є��LQ���ɏ*m�c��l)�b}e��@������*��`�d�ٳM\K|}������`\�.c�W���%��/rz7��FG�B�?��@`y�퐦�u��p����DB?͞q���!\���J=X�ݽ�!mI8�7����)�b����������m��m�E�5��9e�M��p�����ɻ`�J!1*,����K�y�ѦCz{�t��0���d���0B���>����?�D6��5��~�&~�cF����
Mռ\C�j�������ӕ2.����#/0���t�^�����{ҧf����S��!OqN�ANX\oY���f����7�2\o�������.��\�F]��AԱ��w_�_���ڊ�����D?ZC�<3��+#�>].���X�Mq�/�-:CǦ�G��3�Ɖ�$��9sO�w��0*�۬��=��;Y�_���(��G�>��Z��>�ce��I�@�aܸ|����b�Y�ZZG�b�l�/|Ae0����_��Zf�uX��	se�)"����0��o� &F�"b~q=�`i˰�x�[l�SP�6r[ty�,�ϤCc��ޖ��N�I�R,����`�al2n��x7���(U�~�	�b�S�NX��pK�mf��ٕ^�q���g����]�z��oڈ���=ڃ1*>�S�Bd������a�6����n���P��-ά��(����)��դ<8����P�!4Sfm��1c3 -��uH=�ŝz(ly��ot3o������h�9��=�tAc	�\$!��ɉ�z<��e3w��>VfV�����o�+�iz�[�����7s\�i��;�" dҭ'maL�����:{�4O(�͢�:V�qO-S��.HUaV��>l\�>����ṇ�4���%?V�@�@�B�
x%n^"����;�D��4�RZ�����Ъ���W��y�x)g�ɆiǬ'����z��U��W�q^�G@�΅�Qv��.5��z�7J��c��$*%=s�F�-䶓�͗��(�,#�'aE�����|:f����]�� ��\{��B
�{�*)�h�"���W����j�X�f#x�,�a�p���#�Z�n�PB�-^	��l�:y�������SX�W��7]���S���\>�2�a��*
�V���_�.z��Ⱦ��a	���NX���V�;	���~��f���0�x���j�E�d�q'D��:���*P��0�qx�	9ż�D	��dr]�4p���l�tY^�m��$�sZ<:ӏq��,��t�=�A�/�^T�ZLz;4SEm�*�A0?G���Y��x��]�Cm��mR+��fmA㰎�E,�W�La~�����Bc�Ԯ�(Q$�B��@��}?���EK7�����2-0�����9ێ܆e���m1y�ߩԗQݰ�k���NJ"�����2�Q���B��&II�0>�ٕ�24�+�����Ck��i�'�5���%�2ߕ�D]�Ӄx�gN�����l�Lm[z>���G�>�q�6u!Ǐ��!��bq�!A%��hc7�о�LI�>�o��*[[&ܓLOГ���?(���`�'����d`n|�2
�C��B�{�2BZ�������Dͨ������YS��d�YN
�Xh��Lxկ�IN���<Z��,��[8R	77�[�k�IT�Ԗ((���Q<
����B-��)N���6�aJ}��ݞ��>3��t���C�=Sv�K*8�2�f��Kq�5W2j2��ږs.�`���ʄ�j0�i�=Qye��cJ���Q
�}ȭ���r��lXi�*l��Z���+~)�N�(���mRdU��i��t��4)8���a��zx�-�� ����19������;�_����J�([DjB���)Tz���
�ҡe�{p�;^�&*K�Dj^����0�PBq�z���T�r��o:���,���8%*'�j��"�l�ߑc�w�'��	�m�g+�+����k�iӍ�!���u\c��G�8�C~=r���E�┭e��7����U�������l|;�͎��f"�S, ���X����Ԟ'���G\0RQ?ks��4/
�9TnB�cP�����L�_!�������k��&��iyZM�VE
�-�	N4vM�_���	�*{jƸ;�	��K�/:����ն���5����8��RP���K#5!���Ta��� <�b���}������;Ά��r=��|�O4��>�>V+�9_y��Ҫ�����킸�$n��ݢ����;EV���Zӡ{��=���	�w�굚�2 ��Ba|�j��*6����OLa��q���J�ǀ�x�=�%� �� K{c+���)�qc�v:BU���U�¯��_*=�>v�&��s�_*g���2��8�̹��{A�S�_ʑ;-�*����L�N1�T4�o?F����x/�*dE;'�ѩ�̌���������$���j4?�����a���x3���o��:#��CvAn�eL���V�b�v2��@`�X�Q�r��W�SG��`�KVZ7�[8��B�q5A��5�a'А��4��P	IJpq���x��wɓ�� �gO1��_Ș��4�[�0V:�I��j��@X�+�U�O�͏��݉)˰��I�m�t�jY[�X3��Άi��0����h�6t��U�����?_5}��߱�[F���,S�	�=���w����E���,�r�wEu��֎�u�j[�W KX�3���	�u��c��W6��zq�(4ؽ8mN/3��$���˞���m�Ӑ끰
��C�dK ]Ӏja~;�Ʊ�`�X�$��-����n��W�7J݆�͚�|G�����2]D��i��>�p��_6/���(�[�F��D�A�3Y�z����^�g�ԝ(���� P��&wu�2��S�]S�z�PtHL�f��1!�3H���0�W��X�w����!�KY$t��2�՚q_4�����������
^ͼ�$�ؔF6g�#�F		ON�:$�'�Y���a��P6gqÿ́�Y��ڢ�t����tK#D,��`eXVq9)�P�~'^E[`f^� �k����;��~wh���8Wp���V�p����"�:u���Vp���8�a����9��$
��Č�R�$m���v^P����Xs�&U$-d�����-_�=W�c�u���o+�i}��	B��(x괵q[-,f��US�T�����\�����T'�_����9^'�yC�Ƈ,�Ōl��Ǐ7���7�Q�}rq{-҈F�!$�j�� LK�P�t��┼�A����P��"C` (�˞=�7L�z�n)V��S�D�i2]^| �
yU��F�MǬ�_ۖ��{|,^�.�g]ܟ=Fٔ�pe6��r8�T�j��s7�!��mdf%���I���Զ���1�C�=�f<g�ДXx;w��#���iVE��-��0ҷ/ىГr�""|�0�BZJ0$��]����T�]㾅��?�b���'�w�~�0T�1��<r���'����W	�w^:�kϴ��<�]G��L�V�}2���t�{�����?#ۼ[S���DT3j���<8fh7H�vty����#����>(ug|�Z���*��J�iYox�`쳹�p}.�������.�t��;6���U3_U�"���8�:�0_�]F��~�-Azk��䀘�j`ҭ�i%���Fnԁ����q��u��긲��
��
��N�6����<:ݥ���zu�^eB�1��"��J��x/�,ڈ�����;�t7J<�"��D�o�2�
�������mfI&�V����aG&�'�|o�L��p*h�7�]ʬֹ���Ol9���їc��&q0�e�L��K���Շ���Z�ve�tM���[���%1�<���6e⺔ʄk�8d�Z �{y���>�WjS�
�eF\�t����5L�O��ZP�X�G��� r���6W#40�Zk�]�GbE7�{0���G������4퍣���~�v ڗ��W�Z��!|�<^s����;O�r�d�I S�n|�/��$/4`�JQ��V����@�K8�|)_	���)���4c|�`ь����L�8��?~9���p���˭u/�h�нƨ�eH ຯ��Jx��Ux%��a8���6��я��M�VA(�ceşl����Ջ�1��J����u�]Kșp�W��\^%A�񟅸��vz�\R#邧c
v���)��tݤ�h����#=�pe_Tal���!���u�^�X�T�8;e�>��,.��a�V ��AK$��H)z�*rU�ߐ�.�v(��V�{�ݷl/9�(�����FW=�5����A��u�R��J�]�QD��Q��j��p��H;H�R`~�^3����ȧ��I�'^��p1J�DtN�HU������Ӕ/�J�m`�Q7�X�m<zyk��yH	y�J1���X<�3S��C�H.�Zu��\ 4[��H�"7�+b�&o�JHU6�t���������?�!��\ɉ>�;�k"Z�3}��h|���#�e/�a!0���?���'p��|��J�C%�a}o�`M�J-e��~v��)�������������u;�;f��Bd�MK����R��f����h�������Hܱ�h �I�~��pJPw�&e��,��a'
�'V����kt�',��Rn�2������J9u �w�������36�ד�YLf\����������[��i`m��rH�g����4�akp������4��s�bU#}��U�NEi�TsdO^ "Wz����dC&|�Z7���'�$O���"aͮy��(����z��}L�,��ݪ]��q�[��G�=e�W2�k'���� �|�[�$�� �{:/*?Ԗf��נ���A���*�L7�)�d0,Jɷ�O�^��\�6\����o��)9��W~3/�ea���J�c�9�K�=nGk������^�\0�����*�ĥ�;��!����)���Ɠ7�!:K@�G�ȀƘ�q��*�O��d���]D0�W/���(bxo�e}�� �/�g��HM�`,�X� "n�.���k*��clW�F�