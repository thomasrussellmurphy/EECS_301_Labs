��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\���V�fnvx��ÍG_;�ȅe�~�>���9�>��Y;�0G+��X�LP�(#�_�t��� X`�!ΰ��;� �����a�[���~�v]�r�H�R3ﳌ��r�I����f�kZ�ZYHv���`	��]���]ymf�rG{�wZ�j~5ڷKT���}����Uor��*?��c�V�d3���F�����ed�Lb�W��Jf�H�{I�m�?�g�bm�8M�R�B����7�1:�!>.:~B'ŧl.��d`n �N��[Gj�@��J��y>*�k�R~ VM���4y�Bv��К3�O�ʠdB\���p S��hd �j#�(��%��S��3�P�	~p�g��I*�^TB����*H2}�����#Z{��[�@�[��o<O��E��/�v�Yɣ��bɦn(V?����[ ��'��U,�����a��Q�_�P����v��<S,���t �����Ή_�;��y������ �	���ߕ-�i����� �u��^ݞ�����w��s�b�˼Z���9v\r/ j��(��mx�~U���a2�����rsȣ�EЌ������qc����>�:O����z6��xXN����yaD&M�`l�Q��4�&���핏�Jq�LQ���\�O �*&����a�8ғ�������
�ų��;��k��~!�3�!�t���
�g��;�0�IȸnE�R�����5�j�A��(���_z�x5�2
�W�Q*6~~G�ĶL?3����O5_���3y��I_�(�'����5���C����e��~w,�>�e/=g�O	�2c��_Em�s�o�X���Y�,��d'j�1�T������ !��I	8�/�_�;�hV����tj�s�\�������_���s�C�]'|q���du�$�K>����)��@)���	��y^Up�]k�ͺ���+9e|�V��]0V�!���T�a���kJ	�u�MQYt������ܵ��(��w>��PV%Gg��+]�H
��R�- o���9���Ǐ>�����k��f���[
�rw@��`���ǠLz+b�cؔ�KRS��wq�� �%@J\]'h%О�݂�.�����+�I�[�x��!�ʖ�f�� ����Nh:���}Q��	7�$���خ�_��~ �x	-�E'�C�j��Z���AD(��#����d���tR#+5z��u�-�AJ[7�W���
�����H5o1��AJ�ё�G�?Z�X��'��1T�d3MP���.$��
���J#�z����8B_~"���p�_�n �<�4�đ4̟�Y��r�H6���{�?;���ѓ0����������k��9�7㎓jS����o-���[�bT�XM� ���Ljm���u��?y��kf_T=�"�Nˠ��N���T<BwbE��v�YBɤ���B�{�_��E�l��=��/b������۽���K7ϡ0����!T�.K�s`�?'$��m�N�߻D�Ɉs{��x�d�i�T~$Q������/WX���./�A�O���B����j~;\�٬ahx�]&��7qZ�&=� ���!���i�n?�0�c��0zV�P�>��%4�iYL9�
�-4�|��5 6�6&ڇ���R�����ZӹH�L���X���J����鐄�Um�γ���X�
��ɯ��ч(�J+w�XkgsH`^�R��9��V�)e���h�����ha*��Oé[����q��ǵ�"�j�=���1/Z��hE�M�p��t�,�sߥ-���̐���C�����C<�:k����&�Ip��n�f�mv��18�"�cV>����F���;4��?���w�,�ω#ɔu�ˍ�͋��.��O�XTI���<��y�����_�n��E����9�"�A�����'�/���Ƿ�MJ�/8��䣘��۪����z1>����&r��C��$�=��ԙN��Ҿq�]]��˜�P�Ȅ�Cu-ˎM#*���-~JF ����,��v*�)�E�֏��\�<wÜ�1�as%0%2�O��h8�0)�(2���(��Oљ?񮓢��>���Gе<�fU���x��(%�	/�Ʌ���﹟f�܉�DFA�ݸ��Y�5���J&,�\T�q}uB�6Z����OB1^gňggdR���@�ʂ�M�V��5��My!h.�̍M
%���/��?6ZU����YC	����v��j.vC��F�4��`��AT�Ltʊ�K�%e����wܖT���T�1\��l�� ���6�C�d6@����7/�XQ��j���bG��7�ƀ��̤Μ��>t��D��K��K�(����Xφ����Q�� �Ů�T<=\��ׄ�`�I���k�Ȫ���^��,�����ʦC�X9&b/�	F�d:/v��;�;��\�0kg�=c�Ң��H�� ����_�7d�n�3�>��P=ۏ� �)AD���ϟ:�r����rlcv����f����Hq��)i>ߤJ�P���pO�,R���b���&i�X�j�3����Q�qW�jr��z���@*�ޕ�A}�#%yX@�CIK�ݨ#�Y�����*���\�r���n��|^3|6'Z�"߷��u������� �9�}��-ga�
��/^�+�X<��OJ2I䫗�/��;m�ALH-z�*����߆��q1Q2�|�G���N�YۡBOV��x�XHS��U��"��sjQ��t��*�v9ٽ7�ξ&D��#�����:�>�Ʃ���+t-.Q��;��/�G�� �эR��QK�S��g̘�չ8�|�+߿"��ڙ�\�1��gII���r5�� YL]�`7ĵ{���;@�5����Q|�H�>��o�K b���	��f��zU+%�v���:��u�}�<�B�G�˼�_�U�����YBs���u�Na��.KM.��*jv���gܚ>�~��h�Nea�<���\����D���9萤��>�x�˝RH��y��Hp]��%�qc益�2��~�l�7�ߴf�)��DG鶑K7�bh͙�k.�?��CM������Q�Ngq���E�+�cn�Y�4 �����%@�S��>(���v����a�po�7�������!��3�f�_�AF�^;b.LE��?F�>8����2��*I�o9�6�4�W���`,v=�	�^<�I�.s�.�m؟���`q��:vJ�8�nm͢���A��LN��?�����E���e84�bO�3$���#^���Z�\��*m�N��e
���]^%������"��<@P�#������Aeҋ�J�Z��6�pSsR�u�܇d?�Y�7aX]��.�B�t�Q
.�97h�,�I���!'n#S��9;K	蛛�&���ڪv\�K��L���x�iv��3�G���5^�-����U�Ԋ腖>U_�L�K��A��S}��8����g�,�R{�q%�Zk5"���i�KQ^�x���#��������wM}Eȁt�u�רM:N ���@M^X�����04_}i�9��I�5sxT��Fi-�G���u���8��'@d\����$�Pۮ�x]�t�cE�xl��شnjD�d�%������~��	�N,��#OY�12ޫ�s�.����$.���/&+X�m]�>�]G�Ô��LP;v��b.����>���O�~y"��X�ӴwE�#��q"/ά�Sb`�Yp@`{���(�/��]M��^�=�$T�Zʧ�T���}����Ƀ���?�p(�����.N>�n��ͳ$�B�� xԦi�\��n��v��� ��f�.����2(A�,#s9�v�N�w��]uZ� �p�i���C��B_��������$�T�06�G���*$��>�S���Rm�R�	��qH�Ȟ�x�F;A�;NR\��ҭA�)��ث��P�s�d���^j�����%[M�ڛ�C�#0
���K#~ܫw�$���4�yo���p�IL۱r��n2?M�0�~�U7i��}* ��7T s|�W�����MqWIu�&��>�����"t�U��.�RB�i����.jC���`ޱV"փPI�΍��?S�����[�xk�X:2�Ȓ�R��9���x�5�-gm�l�����&6�5s��Obw��H5��ߎ6���j�ƫܴ�O:�D\��Uk)�ivԉ������7����Q��4R:sx¬�V,��|�1@oЪ��N��X������k��H�4�*֒H��|ܖ;~�wE8���� GuP�]����9���S���N5�-��U1�z�A�����e�(���p��E������J���;s6�uaО������^F�V��<g\��Ky_ïZ<dNݞM�K ��ȏ�3��wӟ
�;��I�w} :�v�z���Aٹ��x�N���:G=ʉ85i7
^�`��s��8z6ׇ��s-�512�oϧFaA���α�å���[�]�+;.���*�FCV��x��h<0=\�H�{��m"#KM�L�$�p��HQh�HWඡ?F�q���� ��TA�v�52k��E�\�[��`�|1kw�ͮ�%d
'>��q�>�ωn�:9�]<F.�v8��վ�99ׂQ�?��=nYg�H{`=ñ'���+��5~�m��Y�܇E���}f=>��Y�"�G|_�dͽ�t6[��=ѦZ��d��8��t^
0�\���R[<��KQ��]l{��T�k��'?���,��v�vq�g��{Y|��2�����)E�/�!�F���s��V����;BB{A��+L$�2�Fp��e�yp�ٙj����2���������=���=m1���)q2ʋ��a���&$����������<�/�3���0^�UT���ד­�@'����ʕ*
�|����;����s4�˚Q\�u�^�S(���ܕ�G��vC~r�_�J���a�x]5��N
h������=�{��7�￾'��@cuU8f�=V����yneM�ؠ�H`㣂eM<m�|�� @iȬ
ɭ;X;ò�� �~��@�$��j��/IS�޼� �=���ŭg�1�w�#���l�U��/�&~�"�	C�p�K��V�fQW�����J䦟,ik"}Z�{�\�����[������o�]�a�5Ǖ�ݹC�r��ÆzA�4�Y�z�ⵦK� F�^�{�$?gm>�'�jx[���d��G��S�U]؈�*YzGx�uD�&
j��o�SK�$��?����3�{�<�P��:�����^B�n�2�˟g�7�s�v1��%����q���Z�i��7���ƍ(~3�e��2�iZftlj�i$�x�鵏�b\y-�K:~h��%�zoTI)~��>O@���2Z����(���v���`�*���^.����x�^����Lzt�`.4�4k`�޳���ޏ`H��O�wn���?��(r���\�3;CBV3>E�>�~6�E��k��Y�_ ,���5�Eӟ*VY�o8h��}�>]҉��n6�J��� ���%���O�:��FJWp�#��7l�;�㊍��cFP�2^��XM,k�h���YaB����qC����~������dh9�ޙo���=�NKW茑>[��Um52ܐ,��� �ƼΪ�x�����q�3�}^�Y:t��L_��U�'��8�1?�����4����Sȑ@�[�^cJv��dU�|���x�[�7��`�Pt	h�9�TN��wm\�$�!ň�V�N�V8J�7�x�\@T��<�m�9GG�"�K����!i�P��Ci,W�&i�Jӹ�x�6�� B�d����Ey�l��4�U���}|E�~�&�Ed�Tj���6���@�d����Q1��g�%�ҵ��_M��E�g �䠚�'��Q1y\�R��@����b��}�\3�Üh'��ƕ[��aj����hVN_��³�����}Wӄ���e^a0=��=M�]�?��遯W��Ż,
xIf������sݞ��˷ƛ$%fV���H������+-����Z����"�0�����5��	�Tv�0������D5�Ԡ6-���F�9[���\��&��%�ti,k����~�۟?;Fuuֲ�e��;�~�i`
r_���a϶aeg5��ĮnV�3
���}r~x��Vr�^��T[}+i�>���D�y�)X+����7��?>\�wgӋ��W�H�;��g-�V�QJ�|E:�wS\���yd�C�C�'3i�`�-�%o,�v2�������d^^�k���eN��-G��IE/��uͨ0#�t�3�X���zL	 쓺�x����}~����^�'&��8q�<ZP[�,
�h?�q�*�S�:������A�ֺ��u��:)�_P�����<:QN��;f�9��F=/�U�j��rJ�y9!�@Z4"_&�iK%�A��O��^���A��w����ꂉ{�{�b��F�©�98_����)�"َ�;z�&P�t4T3�/�!�p_q ����Ya�@�A��B����br�>_9���Mj��X����Á�aE+?��3xll�����^\<�%%^H) NI{t-���.0S��U�>����$!�]= %��FR�~O" 6�d�^�]�� J�,�γ^f�N���c��s��Ϸj}��z)$�W̄рo���5U���/�g Ǯ~+&�!r'�:|tyk\�����<��h	(	C�L2���`v8�6� ƃ��d�=2�/�'�׭��BN���-��+��S���@�o/װe�6����� �GYo��j�=�(�m#��g�
�����ja49"w�����T�A�퇦��/�Iin�Z��d���ʻ9�B#$�o)_��T�8Å�PPWy	�;��5��!�@A�|�c�7��3�7c��ݳH[�Tg��^T��?��^o�ϥaN�#���A%��.�*�4Ua"a�+%}�Xg��~����7V�ޥa/mhH��zK1�5�u~���F! &oVYJ���D�<��<v�/P�{�/G�x�����R4�I��t�����W�3��B������-:(cfׯ�ơvyl��4$�1[+��	x(������e!���a�}8NZ쾴�lc�%����Y�B��t=}���.;U��~ݙ�W��rx�g�/�vgS�$M_���X�?��a%�����.}C�8 o�T{��Lo�*���u�_(�!�B�,�Vܝ{�Sy'����h!ۀ��C>u���_g4��g��k�c2L�0���r*�T������_heוH��em����=V?�T��:�"�W
1���ܻ���$4��r�nXI�b�K�����I���*�����A�'�b95���Go�?ղWђ%y�o��	Y��'��O�d7i^�h�*BX���4��r�lM�+㕄e���?���'$.�93/[9�@G�ߌ�j\4	�w�_}O��Kd9
y�;x��̀�4�K6DOpd_�����6����(~�( <�N��#b��{?G&�'���ia�]B�L��Ϫ٫���Y�=M���k�8�`q5��b��n����]�����|@t��ɞ7�N_�S��=�*�H���I�V��O�jZc�q9S|�(��F��}'N�t��e�>c��&{�Ef��"�ګ�
�/�͸j(�M��+�P�W,��bA�v3�?��8���$�s�a�@������=�g.�jV�.�;ç ��4*3ؔG�~6���=)����[=b��ΌQ���̛Η! ��I��K+�
��H	�*�w;���`�d^q�<�y��}o�6+� ���i���.r��'^�1�{��Ùj�	�ikK"�g�0a-w
<�uk{1;���P^��cX�F'ˢ�]3�|��s�SB�23��8Ͳݏc'o!�C��^X[nw�m_��\ְŦ�c^-C�<���d�G�4)h'� ��%��:F3\t�ڭϠ[3��,�#d��JH���ԕ;��H�C��(T��[}�ʤA(�߆x�VDP���b�?@~�+�y�i���ȱ���ɠX"��wdP�Atu�����bX��]߿� �����6 �d��°��>�l�4R�~�<Y�R��SU�5�=!�gsŋ�����T�8�зŪ%��Z�aE9[:�.�}��~&c	�*��K$Ьl�T���O�7Y�*���Ue/�(G�R�6�q�ب��z~�_��8�W���6�)�ҍ}e���Z�=`^���d����8����^��Nf��M��P��[:�=�߷�k�����Ŕۓ�h�li������Ns���V�a����Y��������M0�/��8Ś�v��cmA��+���~�W{DƇKr�_>.�A(:��c�x?��~eAt����f�v�^'�Zts�bc��X+$�������C��yrtg٥{/W��d@��Ѣ@2�!ql޵T 5�������G�t���~::�J��K|t�]��0�}O���7�����GH=���gN���I)�����O��ϵ�z"u��j���r��?PA.�8	7;߈���ݭ��T!I%JY�Y���
���@�oӃ���Nh�}��6޺Kx�]y~u��M����f�L����L�_�r�	
�8��j��Ϝ��D��#�l�7�O]��H<g6��ân�L�F�1���b��,�^��^��gp+����#tqWa�>{���żS9�/�w��nΖ��鼈뛌v�+5f� 1�2�z��l/�1�'nA^axhƠ�ȗ&2��#��]Ѝ?r:G%J�Z�6w�T�q�o�Z�_Z��(0�i��6%�O�L5p�?�>�^+��w���վ?Ż��nQv�Z�MV*-'�u.C�"��?o�xe�Ȫ��������}��ʟ<��1��h*j���*=��aͳ��[Tۯ�t�"20�b�;B�1V��5fi�D����C6Ѹ