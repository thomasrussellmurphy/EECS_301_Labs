��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\���V�fnvx��ÍG_;�ȅe�~�>���9�>��Y;�0G�J	m�_;���?�[�f.(ܬi��3[.��$�]1�	��IhX��sNs���,�7��ۏ<��i�e�-��Q���A�2�y5f�,x��I�0�c`�l�|JXs����{
E��q?�b|1/�QŁ-
��>X���k��	��{�-It���j�b�.����9;w�^I�����jJ����2�< 0ynu�\`+���Yѫ�v`�=���/W�̭�u�ǟy+�er��1�����M�2e[R1��ۡ��_�n�43W_Wʭ�ugs���,��blʉ��;w��,"�'��ʛ�)<�F�d�"G���ʐ?���Њ^���gw_N��]������@�3�̩�IԴ1*�+�
fT�~��+Bݾz.gZF��'�Ag@� C������VX&jף���$����٣GV�Ŵ�Z�Z�	D[�񔯋T�y���̮�iϴ����?&����k���v��C��f�;j�2O�T�i����)f\�%�֒=��=[�X�^Ǥyt�g4�߉"mrJ"<Մ /^i�!H��*n4��X��Iz-:�K�D�Q��i�2�b@Wѫ��� $!Iꮼ�Z�B�=������2~���!J�UrDTӞP���T0�l�8͢����R�vL�^7,��؂�={�J^�TSXS��ZY�>�?�t�%�$��!qf�j�J�~�@�R-�Z�q���=��C}�=��d�/�]�=ɒ�V��X��!:с#�`��Pȼ�fg�M���gu�x�Z�e�Г��I�eR��\�����M�".��z��򞷣a2X����FF7��-	�~���aŇ���	!H#��$�+C�?���v����������q�XL{�Gń��2�"�H
}��Ns��y�_"l�9�k���-W�y	��~H�M#�Q�yu�x�Ǒr5��9]�+�;��x���!u5S�H,uf�.O�V3��<Wb��2X��>Jv�/L)�%Y8Y�-�	��2�	�ҍO���.XsI�y{\H�\����q�l�?SY���
qFb�*����Sv��6f�g�1z��=��5�Ȕ^r-�譧�Ktx
�'�2�XO�/�H�a}
��}�MK����Vڮ$*��N�gl��+(=� ���}EZ%�u~{D?��~��H�5-va�����."���<�s�q�r�D
��c�(�O�����1WP/���D Z+D�J��lwO)n���9��VP�]�[O9���ɒ���NI����\��D���ϚM�j�H�<����l�ј�Z?cYd��_��`�[���r%�t��ܮ����Ò�Qq�-@��+r��ɀX�>���8�ߊ)x��Ǫ�qS����K�c��<��eRX�S��
g��CǙ[�V� ?
�;M�dek~�(ӏ'�{�s��4��VOM�4{�ē-K�d� vÿz�{1�R>����p��vJ71`a�Ko4�s�l��
�{����φ�k~�U�r����?��[s.Nq���,����J�*�̗5$6�>�]�>:jx����܎�	K���Hp�&,�gG��Nj�4�[�����K>�����|K	�أIڑ��*gy:{�i�����D�%�U��U���r�)�=-Sn�i�=q7,Ѩ%�,Gj5�-�̓�}O�Rb���<�a����CȰ��Δ� �-s2��0���`2#s�>VR�$���i����\�*�/j�؟��Դ�P�����e�¥v�7ǿm^l��9��-�ЩQ���4
P
)��#����_T����O<��S"��x�M'�_|��\��q�Ƴ���\�pao�gHs/Mni��Q�K�+�$�=�.w�_�}�142���Ͽ�����I�F/�w�iW���c�rX#��}b��:R{�T�����]ت+�@$>KYk��ͨ��'���9���J�/`c^����*�!�`K��g<��z��9X����<����B��xG����U�#��^Z�G���
L] ��;ߑY��4���Hd	�w�E��V&I�������3W�f+���͵$W������f^���.���<�ԇ乸i���L	�V~hw�l6�٬����n��5t�q��O;&M�C1���s-�`�܂&��fͺj���ֳ;a:��Cb)p���C��`Q6ו�`d� 3��mŗmM�c�mo4ڧ!K����o�o��h/�F:���X�؎T+Ed��Dh|��Q�p�m��$�ɟ��E�ӴU�qAYWz��U~?࢙4T'w���շ�p�8�b3H�l�a�O[gN�z�#m�|��	��߰QN���~�{��@�qų�0�9�B3�k6;�(���m�wZ�M�8q63J@8�ڧ�ZR����L��՛���I ���y��*^p���{&�([�cǱ��)Az
*�0�"��,�N.B˥�g�RJnM��vGO$�D���j.%�G�!�թ��|J�~e�Of޹8j&�Q��Z��9�Q&��_)�����
:0G?4�.��QC�%0�z��@�zO�wB�~���(K���«��t���P�=H�vU+�-����7L�� K�`�F�b���@�-7Ԫu<�Jނ�~��#�r˲5�jxRb��DH���֚9����!�%W�,Ts�A�w�{��*�귦��i���M���65d��}㌯k-�
��x��v���<�W����EP��L_�$Y�Gx::Z{e���I�8�B�����w�!�1���}�ΐ����<�in��(k)g^�5н��\�p�3cKXN�/�g ��240��"�����)0�L��ߜ���}/+Km��cm�=����$��צ�.�Bמ�1<=.8>��Q�p�.�w[����e���o��?�ܻ�y�ߏ4:O�*6r��@�6��8n����]<���d-��Uл��)�q����I3�u�o*)�pp�kf��s=����z����n� �
�\�b�c
J�	�_Zk��߅�����|����+���_���s� �}+�x�����*ɼk<���m�����2�&$��b�ܗ��ƀ?T�ȸ�"9��I^��4=#�5O��ml��QU�B����^�;"�oX�t��ðؔ����OC��|f�y^5�AޣL����
�)QKþ��0��tW㍟`�� U�ފ��}� L�f4�Q
^�~�L ��N
ӂ2UCɘ��*�J2?퉦}ұ;K�gE=�_A���C��V�iB�j�n�v�^�%s)����I����t����j�E�4���D}k	.3��4�t[�eG�y��`�K}6�p���Թv��+*���:@@�Q�eqC��u�Wl��J�+e����v{<�;��9W1���VJܼͳ�i�� �-�2E�Q|���)%�.y�&�x.~r!(��=�EB��eE���|1��4��yː�˽��7�z� ����$J�(���_�z��@�L�]����.���������xà�N��+92�@��Co.���bxe�`���5_��rD6M�D��zw՚ڞl�3 {����m�C%�� [k��EH�M[���z"�T41J�x�XF���yV���6��R7ο����}	�7A����W(v������G�%���8�6�����".�I���+͔�/X���i� �e�n�9�#Ha�O0ȿ��}�b����"�,�n�m���=�9�T�*����qY���5I�h��}�j��>�;�8�
_z����虬.�қ��m��i6򗓸
zl�UĪ����4��:ƑqpI�Q�/'���,��N
���CLN�����\��	��\� ؚ�1_uQ�G���fF��nű���x>u��s�Ò�N��5�/a��U��\�sܻ��T�������*b�3#fqI����Eu�>�kz&�f���}�B����D��-�����ݝ��*/�/o�����K�V�B���H|����'��r=P�\i��p�#�#�W�:sCC'��}���gҨ�1�4n�b#<Б1���-�&���\8>�[ZJ�ү�ST���$ŔuŶ�g�"o��rd����^�N/�IF>�Őv��^Z�Ě�5YV;6�a���Y�I��oȁ�9[����_����X̆'�A"ps�L!�&�6w��[��{�Q��x��?ph���H��<���v
��hX���87�����u��oP>N
S耵�5��C�w���S�w+AB^kƀz�R��؜�B���;�(��/�f��C�����_�0���*���7M��9��(���y~�۟I�M"�(����J&��R
Ir��RyPR�w��3�y�p>��)G��G���?��n߸��b;#=�Ì�H!>��!�Q&C��d��nꕶ�������n����Vf��C~Y�@kT�������V��/%=�|\�I���զ>�����b�@��?S8�<�q��?�x��a��~���:���]��9I��g�g��5���=�k]Q�^�
�"���@��i���C0�uQ�d����3��=�������O�D�
T.�툚�Wi:��{����Mr���:�A3D�۲���_�=
$�wȪ$�{�j��\��u<�S0���j|�}q�`ԭ�0J���;6�]���CO��	�Ճ�]=���a�n�
���ȃ��p�Ѳ��U)�(|ځ_�����-3P��1^��[���Ul�C�?�a�)숦��,��\�[�6 �_=�o������2m�&a���"�W(s1uz�� �N[����� B�.�i��]HC�j�W9m"BO��Lu*���QDl1=�+;��e�ZTS���>�_:N�c��&F�u�E����}�����J�/�ļlf��ھ���Y��V���Bͫ��/wzb�#z�kE� �1����F�/Α�%l����W���(����m�D�ܲ�W�%���tJ?�n�EX�w���o��#��B���c*/��AZɏU)���ↈk"��X閡��s�>B�Ce��D� /��2:����
��u�h����r�"��cQ*8�d)�U`t�H�=ZW58;�s��M�P��Ù���Pvw�|3�	������X��UӤ�Z]�&:���8�,ʑ�ܫ��J�!V͆D��H�0�U̻T��)by1H�*A�Ae!�lUi�Y���~3��ϱ����*�휵�A�!�I��S�ڴ���� tI�����;w,O�1LϠ5�V��6�J����j2.h�A�Q�^Et�����mo�%��i@Q;EM;$X
��Ի�%KT�Ko?�h�\�Y��!�V��I3��K1b>�^���z�=뫙ш���ž�UM����b�p��2��Y�t�>H��l�H�4�2��.�~�7��0��&��ԿK�֭���Q�S��d���3K��JF�� Kd[/6{�S�y���9��S%��6����y^�f�tϻ�ԨoOp}q�Z}�0u�^I�a���>.e+�J�W�Ϣ��L{�y;���,.�}[���ü�7�"0\��!���d?h�;���S�qC���T��5�6r�3��ް'�c������Nl�� EJ��rOG�u�H�T��Wq[Ds-��3g�@(�!~qN��3�j����u-I5W�R���{Ŵ����/7�d�å���`�����3j�Vzh�V�(�/{�eA�-�^#���y��8���N)r23�@Ϣ��u�đB�2 ͛�'u�.^�>p�f�I�r*%󮛁��$(�L qOmP!�e�;lN�`�(�B[������Tw��R�����0���ˇ#5�zƏٺ�uY�+����R��}����BV.q��ibN=2�#���S��2�
�q��b/�<ibVc�� �9U��/f��e{�O��ز|�cvD��	�[��y��*eMo�`>����o��C��\�>RX�^!SͿ�m��
���@⥎�3!��>*^ݣ!n�R��v*!H+l�(���b�/���^������-��EC$� 닮%�?#�_W����V�+�7���XE���5��O�_�-�� hdJ�ie�^Y���1��<��<�Ϸ��>���JR�D� � ���/�r��8IQ���@e�q�a*�i�8�k�]�v�>6�0���;M>{�
B�]���ڌ��Q%�k��[���a�ؘ��.���w).���u�<��	ˏ�D'�fN��51m|k��`-��?��ܹ�4���=�z�Z�=:�oK�1�ٺƭ��G] :�S\=c���$�Z{���"�+~�6��8m���#��[�]p[�2��K�l�M80�x��Ve9����3���P�O.D:�>V`�U����I�q�P6~�Yk8�����P"�j�m����~7��`��F�MZ���ᵹ�QnJҐ �D�`��m�a`�Q(}��"�i��w��
MO5/���j���6�?�����eڧ���"F R��GU{m�����*Į�)9�_f��L��4jk���~�M��b{����W�$帣� 5�L�<�l�X��ƑV߰�r�[�h�U3����`�F�6��#)Ϩ���e1�Zh8���k0}`���������ثj��@L=b����L	�5�	��a㠺�!�g�]R�ǚ<E���4
�"O��'|2t���ԙ����2�{L�:*N�>�2h8&r�h����Ȓ�������^M�Y��'ɔ�z�u� ���r�KBq�(A4XX.ug�eN�tA�+���&@�g
�w�����Q_����W�2�,��ܑ �D~���Ί�.aQw�J��i�h��e���6�
ߘͭCU�J�������əɗ�[����\��K�p�|�T�#���1H��֐� �T��`�G��:2}�m> ��N��$qL$Z`�5+@�(���DLȰ�c���]Q�jqBh��f[$�qY�.n���H�r�{�k��4����Z��ۊ��pƵH�r�?O~S���D���t�S_�K=�V��t5�?�;@�qb� ��,�̶Dd��;K �Ȉ0!�$]�H�z!`+� e8c*���BL��{P1ʕm�+�aR\�K A��D&�}�SQ9A��J��G���R�����/�0��۾0+�J���t�K� �:�S�C/f�ؼ<��k���/��M����((�@~3�ܽB.e�%�' ��/'JJ��ң=~�6��R�����X���>8s�ZiT�^Z�/W��#I�������CiFFO�?���v��_��9o�Z��B����8Q#U�#|?���|��g�Tح�4�<��2���2�����ԡ�n����"k�Q�s|N�9Yn�.혩����p{���_�TC}�f��WmS�+��l]�_���"*QΆH�7�jF���*	aȠ^#�'q聯'�M/'Ud4�0�L�$��?�WH�.Q#�V�������xF��hW����m���j6� �W���B9[L82QY�t"R�:�����;����u�������t��g�ܖ�Z�[-�����!?CJ��PP���
�.���N���W|E� ��!4*M�`[�A�#}YrE���61�������S�?4��W��������'{���O`��jjJ�?�d������i��Y�2UǢ̜�aY'
�m�d�B(��p�X;�XB�VP wRs|��[�S�Cb.�4��̙�6�BzCM�%c���MC�J����F#��?��h�tv�����<�?�My�,�>�զ�����N*�a���G�xG��	Ϋ�q$q{H�e�漣T���[�p���sd�u��N��
E��S�!�"�\6��E� -أ:Χ��)��i7���d�LC�H[uz-�S��j�N�-��b-8 ��n�rcI������yϩ�(+6�c�b�[B",�])��7��)Y���t�"�Q��Y[�ݩ���������f�Mb<��}��G���.Ƹ�ۤ��;����-�O���t�n�F�iq|$��J�1s���GU͒(8��k�\(l�t.o´��QG"T�M?�"f�1��۫T��?�����z�%/�Eb������[���rr���}#7�D`�ȨȈzV�ı<��.�h�j�G��f��cp����,�i,z�0��.�S��P:r�����R(.�w�RH�F�,��,�E�:��|`�{�s�w4U�ÍZ����̧�%��BzHk������
�x9b��v����&x:Y�i-߿e��s�j���)��*"C�Y��bpOR�^Ѽ�~�݃��A�*BHzdc�]��܈ck��i\}/�0r-U)��?��l��T�>(Qn�����Λ���k��q�*R�Zv6�KZA���R�W?/rO���Q������8Q�q����ᵙ�
����-ן)���>� l�"5���O̈N^�{1h��:��ެ=Ͻx�[�V�5�5(9��AB�I?�������F������4