��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�i��a
Α1S%� �uj?�L�3��TLei-3^5]E�$�Լ�N��a��jքy�E����L;��,��Ų�Ǩ�)��!a��\�?��"k��.P�d�f W�N�{��T��Qv~���HY��L�i�H��n�7����l�<y9��@�Q5����/Z���?�|�s57�I�1���S�@�Br|7�� ��i��ʿ��<�Mud�(G-�2	�Rm;�%����;;�4+� 4�W�z}k���iB?�j�vV�e��;�P��/aԙqh }E�Ȼ{	���V�aosR9l��'���k��)ƹ�G�P��2�ܐK=ᴐz|~�:kn�~Sb�pת�^���%ۮNV��N�~�D!�»gLʊ�d_�6~	�P�G��+=��n ��B
��C+)BF����	�^'��cPm�k]�U�j�&ߌ���4���=]"p�Sp�ѷ
u�ۭ���y뫔�KI��n�/��2�+�z��U���g�|��e���i'pB�4�����u<֓�ۻ�4��$���)�^;�f��2Q�:(�W�*�fr�h��֒3�^~5_�S����l����	,�K�聧.��_��	$<���/;!Ce��\c�r�Bj/^bjT<x��с?ϰ���C�fe�ncm�l���7�X._x���և�#+�;�W�w�
�B�{����.p!���:���ݬ��+��-G�u���k!c���|�.�s� �6��>Au3;Y�4�������@i�q�+��a@]P�uB��l���;��B��ɻ�yt�9;y)[P�am���Re�>y}t˫L��i?*ݩ��L����w���ٞ�BA*��ަ*E�ti�s��{���{��l���eYC�7���Gj��9p�2(�:��k�l.t�g/�t��~ÐN�&�0��h�<�e2'��@���0q)۩���9�(c�y��w+8Ux~�{�]5���������}���$��4������� WW\�e/ a���1�妯荤�Oў���?@]��uo�e򝆺�}�/@�̛,4���Q�W����]�wT O*ۺ�(n�;�x����X��@r�]b֛E�JG�F�0���8�����L�J����\�L[�ea�7�a��ܢ�/��⠛W+~��9�Cn�I���[�u���C��B�i��Y~@C�S���+t26�b�C,׆03\�D�I��U�@�����F��8	ɘ�/J�~��n�\��/{{7�2��\������L&W��0"=�C3Ke�l$1�8d���,fZz���f`&ar���av{�ѤCp2�X6\�Q��T��]��\!Q������R�� "+~�˨������tAMhb�r6h�MDv�RU9ƫGҘ� 45���ӬY �$7��6z�7F��g���;������{]_;��Ϥ��#��r�HT<=Ԯ)˿p
� �(= ��N2
L8e��	��\�N��� L�ւu���a̶��ݳ2a��G���@5O���k��?�$�W��/�t��,��m��,5m3E��-'vԜ��d��!~���)�����k����a]�pX�P��O�B�E���LF�Y&�!��J������^��Ι!�)��T��im�c�)x)vɐ9c�KI���.���EH��A�z.�f>��i%�K�T�T%/�Ԙ-�7�no2����ɼW�b�~պ$r�>R�Y%�2-��i��m�b�4c����H`�<��Y�¬t�!�{ ��;����vɝ�im���7��{nP�n�@?(c<1V!/+��x��Te[�y�<I%AW�L���zj��W�Fuɠ�!c�d�XF?���Q}-��J�N���/vX���A-F���1�_�h�\����
�B,���L�2���̢�v{:t ��i���Z�]���)1���n�ƱOx!�������9p]�W'�7���`��wL�؂�=�Ҩ[��	�����Ù~yD^P�g9�w�]ґ�w�G�t쁶s��t��/*�Z �������	u�ݺPG���F����;��mZ<���%\�c�}��&�G�OoK�!��}��,G��H�1�5����̃�RO�У���y�P��K�b��TJ� �$%t�hǕ0�|<;G_Cw�����y�i��8ʚ�)lc�(�~��A�T�-s�5�	"�˝i���q��SUC�Fy�L(�,��f�#X��2�Njӣ�/�6�I�-t�V��ʆ�|�OM�T�	8�n�ш��`��ji�A����Y�Tv'�����*ò1ջ�;w�@(9O#�J�(�7[T�WV�d�,�SZ�=׼,R��(��Mӓ�iC�	ͮ�,̪�`���ֿ�r��pǫNg�m����K��9S�C۔��E���iD�[コT�p��JU�9��r˓c+&�I����e���p�� �)�խC����(>�c�j-M�����Q-�u%n��� �Пl�"�q᷆a	>�~����w�k���=� �(�:p~����"����<};Җh4�P)�:>N�-���򛨣���w��)`W������P�w���V^���>gHO$-9 ˰���0ȯ��V�E��kKl,��'��3���z���,!��p���GxxaX����ǽ��(����߉��U�6��k�],z��#�Ȭ�D�Q }f"ϋ������O�������xmvrha�?_ww-�S�]X3����Gz���*ɉP0�;3�h�#eJ7M���C>	�F�c�b��cJ�\Ѭ7�V��l�'����E���Ȉ� ��hV�z_���j9�hi�qd���XŬ��'H/rcFg�C��K���q���\/�3ϜK��0�Y�%21���Ba�:��c�/��\�@	�d���]�� 	�͢�/��T��>.+
�L3��d�H���������لd�����6���\ %�0!c� ~�e32��Ug�l�%��zH�;����h� �
HM�Nd���[�+x���^.�A#h���G�#L�ӔB1���g�`�����+4������@�p�����O��'��$e�c��\ґ�8Z�#� �wj�m&��:�bn�����bem 1(*����� �R�|T(����OՐ�ҹ<�A�F�5�_��8�t�>n�Ai-��Ƨ�3%i@��錜�Z]�/i��?��ë͒o�(.頼�3��	�paf�mY-/jE��)1�]���%a���	W�Q��b���=Q�Z�J��g�i��6?���X�5�C�h�L��57�@�WvZ���+�I�g���3F���dv8�U�N��Q[.�D�S
&��(L9��;	lm�sK�̢j�ܵ����fB唭�J=�w.ʡ�����c�v
�ޙ"���^�� ��<,�?�����!b@N4�������`�/�q-i5�b	�Z������3��ZQ��)�6��n��+K��G�+�4Q�6T��W�ُ�W� ۾p%�UIw�h�P�]���&����	���~���A
�������py0��~F~�FxWD�������q)e¼`�?�::Pe%8�Ա�rn��E����� �Co����n�k)��]W*~
�		�:)=/\�%Oq�Ґ��?䲃��)�AZ0�������?EM�S�6����D~'|0���q�d-�{���)�W��]����w	N� �l�U;���qO�'JH��4��RUD����
�nP�2���3�L3�)8G�e��Nl�2�͸�T�/�'E�3���r�
���e�Z�%)1���¡\�
�k���N�X���]�*8ž�lʙ<Я#��C�s�LGT I鮄]e�<w���8eq����pQ���5�f-:�.��������V��M�$-��M���iz�d��/�<��Fe�:n�������T{%�IJ_}\*���7x��y�0�]|d�fэ�q���%0H��r�NJ?���/h�7$Hk2lxp��"&���_uӊ;2_�XR7�bzGd�(x��~L�aO����#����M�եC�z��0h��'3��E�xv�U�am���Ͳ2�WKT��c�ܿ����n�j�"��cH9���|�XZue9�2���U����A����W86���ǅ�632<�a�yiB6�8�_b������(�8Wg5��>c�_6ϲ"R1��/o����0��*��=���.�r8}ɏ�U����3Ęrl�v؆l���D��F��1)� "�|b�%��r�*޳~G��C���
2�gv��PK��7+�0Ν������n����h	D��϶7kEZ�Wr�W!�z#�6d�7��Ϝ��i���hzxkL�;��Ebx�!V'@�,�8�GY��GVO�����w?��YT��,7eQ��M�$
}��ޘ=���j>��$G�a�}w��B�p���J�nå��$RX�g;b���d���G=:e��A��^Q!G����T�1@P��E����q��jհ�#�����t�`��d&F�����a�ʱ�����`ađX[[KkÃ�$��=�iy+��+�D����ci�|�� ���m&����>J�X}�f���S�N<U�ة�:S����&&��^�'[AYYį� 睅�+��1p��k�dr����gL{m3H��b�dI{^���x^��
Ȋf�;���+�OVh���Y0 ��{�_�׋�c��5ꜱ���<'��
������9Ş���Q+�#������ȶ�ʥ�_���.@w�<������'�'�܊����O$�P��puO����U ٱG;Y	��Y�I�S剗h2o�CE�hO,Z:���Hf�v���� ^�Q�<���۬f =��>�&1�Ċ���%�Gc�������x��X4�e�g�g4w�f��@���3�.����[vX}l8����̓z�O��Dq}�.�
�~]p�m�9q�p�[�k�Ԑn��o��,T)���@q�P��wt���Gj�㇤��a���,yt�Տ�[;�����R^>@'Z	�`�U༭s'Y1sŇ���ӧ�?�yG�@z���q�]|��Q�at��X��E�vG\��l�";���t�U�ұ+a��7�
x�m�����J0h9Ew�	�1�
+�q�Y=-�glQpg+��J���J2�O�]I�ڤ�w��,��㒈y��v]vѐcj\]I�;��a�q�\�.39��q����o&G��(n2S���/�xq�dk
�]�m?\>>��-���o�<m���n��dɽ�&�daJ����s��`dS�٨D�$�<���0�6�\A�P�F剁��O@����,�i�n�Pt�:���ф�T)(�Hc�(��bQ,��쬲H[T��iBx!#�V���Z�n�Y}�� �-�� l�ip�$>R3��Bܤ���х�=|�,*����2��{�h7F�4l��� ,1�{�D��'u�$�V>Gj�VP�w���D3�m�fu��1�I Q���y)0i-O��W�(�-'l;���iXɈY���9�	��f���n+Ծ.���"�	�Zo���V�ğ�Y����h?���OL\�J��D��~�^L��%?7�ҵ>0u{�~�}˾�e��HE�b7����`!�#ޒ��m�V��B��8ԫ���bkk��*��q1���,Z�k�'����+��}?���G�=�q�����V����p�z=�a8�V�Ӽ"}08_�G��%��#����K���%��\�2��#�l��ɺ�T{�"�_!�i�Bt����e�D���R����f�U B�����T)<�Mp�I�(�����B�'�7�q",{zޓ�mN�5����A���x�XH��+0�ZGMc��R�����6|ӷG��/<;�Hb��Mj�<���E�$����b��d����m����C<��mj�X�����g�e���ϋ�~@��#f4N�@�qS�G~Q6:���b%Z��*�fhW]6z��=&0��-��ݜU�>�/�#��W\��(q���G�y�EBͼXw�	��a��ETh0�;�����d�f�s$y@/��Ӵ#�_�M�DQ*�C'l�08��[x��YͻޱuL��߳��(��q��{!�Q���d��������ߗ��G���v�vUR���?�W.G�C��'���|������x�\�MfC���n�hӵ64۪n�E�D$�U)�F�����X������tpA�^��e��;-���B�S��F�i�|�?���u��K�K�	�_2��׹4����x%���9z
G�y��i-F	��eb~�O�j;5A�og���˾l	`4�Qe���dܚ���M;ꢋ�.��y���nn[���A��̡�`/S�����$�r��׬n���0��+P��\�����%���W��U�P{�(���{
G�/�B�G�Ey�0�(\���N�	 RS�}-����ʐ��g���bQ��ݩ'�ƚ<�ͯeġ��w2�'�o" �/�+���fCVUD_%]�4[�S*�w'{��~p<-%.��y�XvK�%r�$Q�b�X>^�!l)_��X��fƭ���e|�!>a��ű�(n�0�w�?�$3K�}j�榑bR~�ԕAԭuR����]���H�
3���A-�c�ǵ�Eo\�"�N����������nzTZ0��/'�3�<�}B�#�N/��ߠ[1e7V��L�ݏ�=b�?���*��������|�u5�1���T��$��Q�_��%X��&7kR�o���B� *(�~i:�V�2)ٸ:�4�7�����! �9����N�*aí����|?� ~q͎����>u�@���D�ynЯ�v�U�֬�q��ϱ�O7G�2�lnM�CpJ(�v�X��L�k'�� �v�ӹ�0-�����{/�\?�j�]MhS.�̄O�7�2�k-�T�87�+�D���f�n|���{��jCG�*��)G�,}H$>���Z5Ս��IuY�R ��L�@��5�.�Ձ6�k4*�5����x����'PD[���w����Qv��)��B1�?����t��;�����{	��'�vh�s*�i�*:0'[<��������m��>{���P�Vf�`�����7` #t�Z'K]��@��a�F�ZY���ơk�>ؐ��j~���yM�ޠ�NGޕ�����+�w�b�u�4�pL�zf_m�Ǌޅ��D�Շ%-JF�I����P��g��*8�!����áQ��UB�f~�n��:-��b$⫛��o��V�}W�ѲH�B���ձ�<@)M�s��)��tqp�@�dY���S&�MC�kw����HF�1��~��Ȝ#.��U,��P�����Q�_p�����~E�>Od���6 {��R}<�y1��(�W�7�l�{�jz�5Sj�w�Zx��2��Je+p������vU�Ou��])_[�U��:6��v�H��G/+��m�������� ��g���wი?̾���\��J��G$�?`�������S�ir�χm��G�9#,�c3Hz������%& 'k4�D$S��
V����(1p^D5�p�'���N��_�������]�:J��'�D��iI�05�l��4|ũđł�U�Mܐ�`�ܽ�]b�eCS-��i�&r�s^&|�]�?5�#k|����e6(��Q���%���'��ͣ�U�l8��-��z�Y)�f�`�	�kV=���.&�I��B�0~�!�@8q���	1	�@b߯9G��*��G��l˸�ک��/'¥�{��:�"��tM����"�)Xz�[jV2�{t�rh�)z(��]9��y�%�k�˙kXN�$��/��NhD�K�Y8]R#����!������͙�/�@?�T˄�z���taJ��(�xa5w�_����Q̖x\i�5ۢu�?<����"zw<�2�k)]��/?LGz�Tk�s���J���Á/[��
����y�g���
!�Gl5Ħ�y���gS-�q�$_�R�u��Go(����?8s|���5�
.�Z{�m�cd�ԇX'=.�+`9*�fM�R\7�k�g��� �}ܠq�o��ކ��/�<+K}��j
�k�N�2w�j�s����h�bR�j��[j!D�}��U�eBS-X��:����=a����*�ˊ�J��jJ�(�KY��Ԉ%���E��g�94���ZEԨ�Z�o�}+fd�8v��䥖;��o�H}_2�-��q[�vY��9�A��)8�!�g����~�-Ւ�Q�T@�r#���R���)�o��'G)��aaB>�p�m\�J�&���H)A1��M��Hs��Q�� �P%���/�fN�"9��J��g[��2{�������+>���ݶi1��uŪ��of�u���e��� �c0�
F���$��Y3��6ʝ'm�j�I�#�J��,aC��/v-��,�b�g7�qnᨇ�:�C,����}0��(�#�t�tx��>�qa���Imff�)0z����� 2<�QlY���d!�!]�Lm���~�-t�d�͏&�7�V�kz���W���2HL5X���|�9�Ȇ�툷g�.�>{�y���wߕ
Wۦh1��2�<n���'"
�j3b��kދ�V��d{��/���|<�#�ٮph���T`�<gL!���տ�+���n���h@��J��8���U��%+���K���Xޗ*JV�
�3b�b���������i��ߍ�'��]a@���mT�<k�O��`v�����.�y��y9��q�?�՛���#2��C���n�N����w�)�+~����[����ɘl�`�S�5�ۿ� �M��P�S���Dd�����hL��p��=vZ�0,�T4�\I#���\�]�i�3���#yLLk�C��B`��?�$� �E�S�="$4	0��4M��N-��1��wm���S��꧍����Ј���H�����}�����:$�`d�"A�B
>���U�#�S�Eb��`�2:��ӶP�ϤcJ���R��n>W�LY�z؏|h�{���t��yτS��3��	�i��2��t��,߅B�Vgf^Ce �+}�4�+���������N��ا�-���.�����DՑ�5E�C� �1$�9�'8�LH�������g��+ ����_�p��6
���V:q3�xrb�Vh�W�<����`?{��.��v)\���yd}�$�Rz��$�=/�&�#o�Е��C�~�(]�My��v�����W3�+ )���$8iD��	Ϩ�'��,��qh��;����U���
,H��"�������)4���y�}��+�`�r-LJs�ۋŮ��Y�VɚD�σ$3���Cz�l�z~�+9��9'3�Z�?�c�d�Ҙz�4�v��S�r��&��ZGCt=����Jm2:�F�.D�����2�b��&ge��d��N~���um�Q��b��@�#q[UG�[Q3��-ü�`nd�U<Qxn!!�]����4��Ie9���3>�4u���
vE�v�E9k
��h���8Y��ɝ5�=�pY�mԊ��>����y�I���7����=k�6(�Qo����p�^f_�a�p��5/��̫��{
v@���s��	�sP�Y��Z��Z/�#"os�B|B�I���.ߊx�g�j�-�B�&Hz�*E�6�c�%�6�T�p+�R�ݪmRdi����DR	>q+��O�%j�!�M�n%
�v[���+K�DKE���C5��
�R�ϵ.�_XՐ!��*X�O�B��d�ew���v�#�J��U�Y2f>�ČwKE�`��ʄ��R���3�����^e� �E�~�����}��}%)�iu�����C>ف`2
b,K	�A�U]�(0�����WJ��F�;K��`���+ZZ�nk��\��#2��ۣӡb��1�S���x��ë�O�Fܷ�:�bM�p��xK�ʹ�<Y�q`0�)�éw��̛5��PQ\)p��?��B.�E!=���Ys�d�T�m�/Уᚍ���O��ՔnU���U�@t+�F�곬�yJP�|�/�J�]Vt��џ���ZQ>�*4$2c�`�R aО��ԋ�Y��7(#�r;y��;���NJ�SDe��=�"�nQ��;`�~T�,QR�w���������;#��� ��c�Q=�&vK���F:G�!�^"��<�x��c80���˴�F���?��2��$��G�DE��ވٷG���1�� ->��b�W/=b����3�,`��_�L+�m%�Q�J�9W��3߶���	�xT��L �M�g���c��vK��!H�s��}O�:�#v��\�^�l�%��8(�mZ�35��-0�r�>�"����Q��7�v��椪��s� _�%Lm�a`���ggYج�sV�dD7�VQ�澩�y�C꓂���Z2��I
�X��9+l�����0�LQ�{r~*4৑����K1��[Eޔ���#�
	!��B
�Dx1�+L��6o�R{���i�`��C�:�Uǳ��s�㥇�C'��)�V�>�ݨ��@�:�����!� q�����sЁR�!6X1����6��.0��)"�����_�P� ������A�]�ux =xw����ͮ�d~OS��ҝ舄���{��&�1����4=�f;t��5�A�a�o���f%�q�bSz%/�q�/�`�	�E��W2�\!�B|��W�а>�G�n,�ifP��5���'�p�b+t� ��NZ����������a�-�ls���[5n|b;"N�⁆���ՙԊ8��q���/�)n1`b���+�-W=8s-e��IFy��EV�Y5�L;�_�ǈ�NpSj� ��Z�2g�e�}���Ͽ�u��*]�xHhT0�L,Y����.ى9~�%�+Q���7��D|��T��tD
j���̆pC�D�_?C�C�2�]��=���8=7���v�z��[��
G2S�!��$ڻ5%h�/D���!����#�a��C#�
�)xI�n2 ��Әv�4hlw&�|����i�N�	I���g"x<t19�˔Q���!D� ��I�xU�I1-R�`4]��`(�j@fڏ�ۮ�0Z*X����K����,�j큄�T8њ��a!���П�{n%p���hM���Lڨp��k"�萐�e�Q�^=�rZ����(���z3)� �h��b?aDm�]˛ �7O3 �Z��wL[)p�HGDi�'�Vل�q�-fU�]me��r]��`�Ğ�v�eWD(���E�5���ۡ^b��:��6.�W���I��R��d?���_.���O��u�$�7�s}�z�X+�E~��l��N<p�3�C�%SM@��<Xo�ӛ��~<N����^�kyi�g�ȌŸY���s:t^#���$���N�H������f�,~Z'���]Hb� ��+J���)�́5
�N4@:9.-�v%`�[C�<�g8�&�(��=M��
�Hy��\��V���_R}B|q#���� M[�q�n��_=�=L��Y�-�5A��g�uf6∧�'G""m�U|6��$ˑ(z��[���n��4�	��v�����e�^�e�#�`H�#C��c�B���eBE���t�֗�ey�=�C���
��+�e���er0
}4��#�� �����3�rŒs]0O*\�C�;�j����D�z�
��aFﴪ؂��"���3���7)���H-��3�����	)����񭼿@#(&I�p	}�'`�
=�ХOu��Eu1UH8-ˬ�7� $1�S�����"}�"����"��������;��L�&=t�t3W^J�ո4
��	����ԡ�J1��M��/\
 P�0����_նb8B�.cF�:8��S�UA!}iM��3N9�<;<,lM�H�Y���L:�z����ɂ	���&�_�5�"ա5��7�L.m�l_�F�Y��N?�t+��%���A�3cD��+"�LOe6=8�j����&r0��
7�˙�+a~�d��aQ����@ź��oFf0萎���|O����KGJ�:��=��{��
];n.�� �0[��rd�d��e��CX������C�z`�G���4�?�Ԍ�œ4bf��zh�(����(D��_*R?$��^��C$P�9)8b��W�yX̧��i�mQ"��f���5o�L�4jp�;jحD��X��J�Q���^=�lj���R�Wg�2[_U;WM���٨ط�q�#W~%�ﯘ]u����Te-��袪�5��߅�㭰B���~iٛ��l�	ѷu%�s� �t����+�������qI��k[Ů��ٝRkOK��P�0�`���`I3��-��}d{FO*�C���cE���3fCkw��W���
O��N�bO
�������o�y!�([Y���z�Bq��1�0��V��
kY��/���U�]]���f)�c�����H`y�yq��1��i`-��%��\����]��]S��v�dW�D՟t�D�ڢ�Z�%i��;�>����Xy*-�1o�k���'����,���c�;E���g��\��b'�.)���\/X��4xjY��-��]�����6��uD��b)K݇
����.�Iگt4&��>��k�Lu=�Cm6Mm���S��;����J�FjnW�-�t�06�R��ҍ
�-/CVV%'�
y��s���%��%�G�d���~���<�Hf�]�s]xE�y��v�E�Q8�V�����̘Sl�II�H�`^>�*ip�A�BM=2��U&���?�j҇����9�_Yq)���&�r�E�x�4爇^�o�ٻ�!V��!u�H�w�L��7����z5ϓ��{�?g�9��_���c��AH4-Xd|q?�4�yP��*��x�-���Ye#�~����%���R���x��s׷ }��3���0�3��!���'w�����Xxh������p�#�A�fɧmU�u������?�1�p@ȟ�	�C[+]ÐD�2=�;[��v]��6���Ҵ=�L �j��H�P���Ҿ�VLwԯ�=�ܰ�������
�M�#�44dCy���w�|Q�*CO��U+��H?�IIL˻T`��s8�^��l&�.�b��Y��mpi<�Ԛ�:?�F�2-���1�V�
+c�`H�1D=ف��T�!�a��'y{O�_G>7h�-�9<3�S�M1M������_Y`�������N0G[!�7�B7����/j��j+��ب�|��W�n	���b�6q��������s�UU�������V��10#A����\���=>�ۼ�k��b6�6�E8�>���R��7�k8���?YK��������� �N�|�=�9sX��,V�^-�ƭ����4���
��!��P�?~��xT�|82�r���ϲ\��F��;���n0�ve>)_�T3��������%�CL�8M��Y,���^%iJ'����h���+g��uQ�N�5[uyB�9��N38���^���t�m5���+)V2Q��כ�4!��h>6�\ү!��(��UG@����5����E�~�LVf���ݬ�7pw���F�AH�,������.b8(K-�����Oq�i�3�*���ע{'5 �Q��B�
n�԰�6�ix�׷�Ѓ���x�ԁ��B�0ZXۀ�x�����Z�0���^K:$�<����Ѯ��kL�7�z¡���b�����<�O1s��Ǘ�o�t�b�Ա�RE'�'7��9x��[�����������������:��Y�����j}`\9��#�0����A����;&��z3�ƀ3h�#6��U�Ρ>�:�`BK���~6�vf*�^
U�t�۷{D��}���K� 6K�_�]Z�l��m�s���|����#����]�H�o��m6��b"�u��LB��y�8�+�-r#m�A��AwDv��9g-�*����i����*[8yg̞x��*�N��V� �rM��"c "i��~2�B�T�V0}'߮��?�Y���h<��|}�C�|�Lf�wq>8����� �z�n�����B�_��~U+������>o�\��LX��&� 0��e�Eg�r2%N��VG3� N3Y�R,��q[�29O�2�p���d���Ą ˲��dà�=�=�}f�&��8	��������=��n.خ���tn���hU_���Q�#E�Ǚ�A��O�4�!�6κ��Y%�!3i�����\�f+͊����	j�gh�����^a�ndE��^L�F�����F-$��5���ǅ�6K���J�U��(�-��d�g]���aeg/�4���1	r3���Kbyn������FYZ=�,�2|��	#��gN�"C9J���_�M �4c/�8 #*�+�^�qw|l���âv-��ز ����پWs b��+�_�t��'8|�B��4�dE�[�f�P#�F�� �&���V��ߟ� &c��H'�((�E��]���Cj�B|u���0p�8v@\�W�O10̬�f~ί� ��c�9V��h�tt�w��#��:R�?��g��i"I�U��si4�/u���XK� �LI�"�=``�x�������\�|��B��cAS-�:Ѓ����&�����)A∌5A��,ǎL�ئr'쮡�ȇ���5�;����0z�J��?�~��xPZ�����!b��h��}����K���p����
�ϗ1��C3����\��T��&��S�M�p�?����j׳�qR��@��h8�v��K�1_z�����Ƅ) ���I#�=�W����v�O�i��� +x3�f9;�.76�5b��.7��Kw_kղ��h�;@K���b3n*��^+��%�i)�TNN��Ҏp�ۣ�SX���,����W&B��x@|�Rw����Af�R���=�f\���r����6�ʷ�	���\'�.�L�>�F��`W����XGM�&C��qՏ��M��P�mRf�%��M~:�.����Kp�#M=^�+a��ׇϥƓ��,�8���e���[�Uۚv�����=Pxm�KX��+����v/!<M��a�X��l�PJ��+%-w�&�.�@ܯ��eyB� V����Z<�`F+���	 ӧ<OݰZ�c���+LV��ތ�P�֌�4I�gH9����f�Uي�ZZ1� ��f�1���R �d�iG�?�@O��S2�$�CRwM���cz�' �	��u~��S[�� D�Ph����Y�63��Hg}��^̰ �P�z��D�Ӡ뾰�F�䍻%4!�w� 	�����5�c�۳�`=�܌*T�V�t/���ӋK������TW���pA5��k��u�̞�Z����:�M7��i2L�a!(�`:���'���z���qt�F�w�	�� �	�@�T���5���1I���aDX��,RԱ<tF�כ�4s���j��_o�0n�~�&'�}1<���mF:otGe�6���w)��#��(�ʟ��?џٺJ�-�N�)�N-�a��Y���n�͘�H}_KoTJ���a��9Y��L�K���
����/2]O��6[ 5v�B5jR�^C�{BE�c�:���a"t*s fȰ7=At���0I�=�Ӗ!:�h͵X���7--��9eO�^�bCKn��	�/���������|���o>�6�7p��n�)���hL�BŃ�,:�beӘ,o)���%}�0а��^#_\�bAƷ!k��btv�"����ҽ��ֿN�Y����⚲���^�8b�n�G_Y�P;�$XS{��C��(L��uZ�g,_~��Us&@UB�(</�/���/2��+�]8�@�եhz�Vo�d+�eo+��}��8(�;l�n��[���D��'���z��0>G�'v��!�Fa��/��3L�kG"�Y�0�4L��~5�2�k����[�ø�/1+{�����܍��ݠ�ΙZKB^`�҆*k���(/&���كJ��U0W��w���C�z_��%�'��E��hV�ϣ�/�a���p��ۼT��zD�<��d4ܚ���房��&�\JJ�� �{�i/��E�T�Y���^�v�Խ�̉at���Cn͜�BjLc�4�7{�z�a��3
s^���<�@���ٯ�*�D��f�(���(ȫ�b.� ~��/��(k=�aJ U�c_�jY> :6jO�	���QkA���}�z��9�j31��9/�i*<yr��6P�g���4�ڳv�:��a�E0��g�����= �]��:�C�h��\�&'���OL��>��e���p�M�̐2`�GK�Lb��gu,���u�P�x��Iκ��rh�$#1�4r�UxRs�ٌ��^���]��|p�ة�ύǬs��l[~�a��b}4�s��� }��Lm�5�K4�E'5�e/+�&�ۅ�|u���oX���.,:]|����N�o��^(�u�Z�v�M|5�8g������k �Y�v(����;܉7�)�ki��^5������k`��Cd���� ���� ��:��CgΦ�tZۇ~]�f����P�S��/	N!�q@��\NH馊��h���@�D�E"3�	����e�b�p7:�'��}۳\�w�yV����?�6����x����6	��&@�B�@�D��}�N�P�������:m��n�d�%JEKkD5{r������[�����F|��Ӈ�3&�&�ys�Yh��7�3.���kb��y?ᓝ,tm~�H4�s �IG����(�//v����e�a�D�6FJ<��5�'Ы�׿���+�j�)}EƵvz(�ݨ�b5!�H�:��z;�^������R��췬/����ۢ�R���%�e��+��у�����ɮeŵ/п�1����ꇬr�:����F�'�sQ��Dz:g����5�{�2�-+
�>����ޮ�:����hy!z��۬���-����>I�f2���6�{�,}�\�x����=e�I2i����秎��3fԉ	P<�qe:�m���g�>���o�%_���Y���f!��cAɇ��5pp�3�t᜝�B󛿡9M5�aª'!�|���+N��3R�������#�NI����Օ���)�>r�����$��;K����*N��ȳC{4_p�H֭2gsb;$�fn��\�B�� cB,�x�'��K�� �Cj��1�g >E��ϷM@u	<I�d���݄���#{(�U1��q�m�㸰]=�� j���M%�u��X�RB6����=|N�ǝ�����6��@��ݔd�M�ق����)q�o�Z"B�mS4���(��I� �4���kjuҔ�yf� S/���FY�'���Ԝ?_gWv��RH6Wo�7��/T�X��Ҵ�4����ܰ��)h*�Y�|��A�$�n ?�]�^�KH�N��-�o{�?�}�� R!� ��[ 
��=�D�#g#�L�#�f�ު ���ռ"n�v�4`���:���[[J�����)l-2��Û(�DȾ�*�zh1�1���S����g�����(��t[a�a��?!;�d��+� �\���l|y	�2�./�]�[p�Vw�>�~��l͌|�m�z�-[#��τ+9�¶i^#���;P���8�w���h�ya�P�Ĺ2i(yٴ=n�_8�L�_�6d�#�q�[fw�LՊk��0�d�4���#�~З|3�¯�)�0�X�h�cG���d����&�EF���k�����$"3MV��c���/�A���ܮ�祷�$HP<2*G�S�U�Q�MW�3MN���k���rn�
�������~I҇* Ȝk�pB��)�A���3�
��3V�ͪĐ�j=T���>�����ü.ñ'�f�'���f�-�=�����0�L��()Fm�d��2�~�t�����&I��L�("�z�~���|�[������*���s�Ʈ+�י��6踼��J��h)<~1�^��`��s���.LaЇ�9�g��m��p<��@O���g̺)����a�?h����g�V~��=|���[`y��#x%�|V],@���E�J&'�.�k>��"��s��?�Ż����+G��-��=<|]k��]��d�ĻW��Bh�Q^��&�4�_�Y�!��T� ��IXq�:��wNz�1�T��s�9���9\�������W�K�&BP=��Ş�@���I�, �{���'�p�Sp�c�8y)W@-�/6�a�ʅ�v�=삐VՃ� (�Ǩ�hKR�6t�v��P�$�Ȣ���U?�P�F��o?�k�Np��"m����}��(tJ����FQ�f8�c;��@9 �l_s�1���Y�қ�Jk���B�#?5�}!�+���fQ����E~�]�Mb-�s���
��Q�%����6��.����j��! ���dJa�����2��?�Rqy��H�\��	#b�z��E٭ Q�#��=Y���8���k�a(�OUH����O�B�Q�T�#)�Hz93���|u��2M������i�����+�`'����sk'����rm��9E�ݤ�z������)�� }ő6���۰�9����FN�;x�J����� �r�/1���G��FI��~�ҁ�ө�o~_��C���?	�֖�ݺ��q`��5�"�t`U~��a���̂،)��3<����nq�)`��Tg3��Ky�cn�i�
���?�	�[��>]v�'v�kj�����zT)z(Ό�6�ƭ�Sy�"�K�Q-4V�R�J��ه�i%%��'YʰS%g�Q��4����ء����-Yδ����)���:�7@̴\Y�{���
Y��r&�˪a��7t�¢9	��"���a�}����:�����{��{��E�o���IUdP��0sj��R�E���\4}���8�ʏ;��9q�cn�о�Cw���+L55�*����0��%Lr���]�}Q�}U!��}T]��2ᔆ�-0. E<dzָ��$������X!H���ءB�%�8��� ~Ɏh����5��Li�d$c��;}��,{��a���:3��v�S��3�<[I�d�EV������O��U�d�H�-���^�z$c�ab����f6w-0V�i�Z�Jt���&L�*P9��yE8��`()����u�ɜ*HՄ��Nч�trg�T���_Պ�(�7^һ���⅌	�JO���PB؍�y��}aǃ�i$��fQ�D�&�Fվ7*�	�}�n��\�l��˲.��GҨ�a\��_7}0���r+�#�̙N>nmv&֘������%�@D�X0(%�ާ#��[[(uO�v��g� �Χ~WH��B�7�I4f}��Ev�Mv=j�Q)��~ŷOz'kz��UKx���by�-�y�����To�/�hg���T���A?���Υ�5l��*L��_��7�G���"���Q��bG�h�5+���~l 	�M)����)rz�?�?�ی�r�/`|�T������_~��?�x�+�_� =�?@���@�c�elmI�}a����2�����j*s�Oi3���-������[6�4��{Rp.����4�B�F�06���K�k�l�3}?��Z$N�B�l��C��C�N�8?���6N�ˍ�����z����죺$_"!J?�ߣ���:9�u댈@���7��X����J(�����M'�LI���������բ�!��)M�v�0��h#��������wUݝ!.����[��)������4N.�,��̶ڳ��B�.	\Y�Z��
/�B!�R2Е���2Ru�Gl��$�'����y�|����D8��������sPق�]br�
�Z@�8����;��6�pqM�� z)�̜f���a%"�<����e{�W,���y`�%�l��,^��J��oG,o�l&���t������n4n������]�~�����Sc��_/�g)@����e?5��3�
�B���csl�~��f�O}��2�������\����f~?V�vP.8��vv�� ����)�HsS��;�g�.���E����o뒝h",7�G8�0~�[�'��y
�#��^zM�},�3Ͼ�溎s!��u��J�5O�9B�-��-�����=��,��\�K�;����ٗø�r渭N�%A	@۰��n'%C��� ��C��ȧAN�_�)œ��%Cс�[2)�����'��RLL�mY�����_<G�O.M��b/b���kr�,`G���^�v	m&����{}��T���*��X��n�M��}��F3���6�cy�Dc����&8�1_#؍�j����e�-/�Xҳ/�rJ�����2t!�����/њ��W(�����'�FM�m@!��A�?�<RYC�;��B�) %�0,�@땫Bh�5f�K,�@[��x�����[���_aL��'���b�<��]b���=[��Z�%E�������{�]�A���Su̽I@��wY���K;��=�0
��=)�NR�[�(ooky��z3��X&? ���J=X����~a���QU�@ �A�͛��⁧ju҃"�]���;0�o_�s`9�<.aД<����xȍo	�4e���m����q�QK/z>�C��m��#cr8����w��0X��뜫��-�ty�X���C��<�6@R8���8h�z0���Ey����I^�Zw��+ ���>æ� Y� J!Ps5a�t�����G\��&�����c=H��;#�ز:!r���"���d�+
x���H��F������xA�pdV�
���y	�Z����k��������:���J����� R�m�B"�w�i�9�P�
��6]˿`��6�*�w. ��-��@)NM�aL�D�I�
c]�{)�b.�3�&h]7����Y�c��q�_MV��V�����~�VH(���ױ�R�E0��k�1[ixg)�$����W�	�?��0��&� ��ᨵGq�M�zd�)�]'?69<~���	}�0M��{���*Nߌ�
ZX֊����f�{�vy�i�ǗEd�A5��Ѿv��G����,x��(F׸z���b��4��PE����QXO^ih�����V����.�4��>�Έ�vD\����Y@�o��҃�B���A��x�mS�Χ�U�7M)ԏ�*�ɔ��xsM(<ce�5�J�"^ Ex��u�i"�y����z���*	?�lv���I-WL5��}$0Gcm��b��|�z�m# {败�}���]& (o?���u��H�ǎ��[��ج"��;��X?C�͚�;ֳ�zFk���Q8���Rχ�F�MR��|��+B�q�C�{��_�d֏Δd���PS��i��ȟ��[�YW	� ―D�f�A[/�ǚ��Hy�/��Nd���д��ujk�����	�4�̃8��� w����d�N���j��iX�3�h2��r�5���V�@&��w�{@��*�l^C(r/���b]�1L�S��FS����k�t�eB��>�:�ͮ��X	oRBH4��m�-k/y��I�%P�Ÿ��#���&K����#?��p��F�!(6�e�l�o�``YQ���2�r�Mو�,,�1���+�������g:�)kn~D Q������b���I�Ev�Tk���̹��۾@~o
jͬL C�����f�G���
�W�t�~�4$u��Q�fF����v�]+�!�M���Ĺ������͔R�3���P�ʝl����
5#ԛ�?(���VB��>�C��y��p�P T6���W&`e⽂�0�͇�o٣xGI�����RKK���4�^�����is) pW�
 ~�j��ൂ�{<�6դHO��K<�4��K��jF�,�%���m/7��]8���UЭٟ�vҖ���Ǉ�ٰ�}$���fL��V��\���2�9i��#M��d�^�hX�"x-4�<���=�w��<�O�J�1��f��AE�V���?H�l���*RI�Ȅ)ÝJ��E,k���0�V�5����:1���7A 9�`NWWm���u�-U��l�27u��%��ų
Tt�Vy�1�5��S2���!j�υ�h�\���`�&1�t�&�Ij�cr���B�n�%5���"��K'�����WQ��5��0�932'��%��?����ᦽF������v���'�aO5�/�$v2�ƕ��II}(���fh�ݿ�.�%�M������[բ���u��!��h�.�;��lZW�ˍ`������ϴ���}�$Y�2�Q�����܍s� �A����r��ՙ��֕�x��n8��MVY{��y��CI� y��?��)s.�+���5f���#G��y����?�� X�1r�04ͨ�Ǹ1��N��Y<b1O�|��B ���V�f<�$FUY�Q����E*7���e��W`�]J[W���N��;
�Gc�e����ڎ<�pJ��{^�@�]�=������:�Q���i���5���ñ�S>�gH�8���|���6�����f6jt��<��V����l&��Y��a�s5��
����!�����C02��3����	"��݁1�#�)��!�â19�?:*������{�ġ�J�e$1�������n�����׸/U�<���~j�(�|؁�w֮�:֞��?vH|��h�|}�F5�ܾɃ����$hfR�oLրS�~��*D���-Q#�vׄUܱ\�kh8�B
݊��E�Z� ͱ�TQ[�ap���M��\i["�A&�ߖϦ"1�t��Z̙����ηܖ��%�x���x����^hVś��;e��+}�M���}�i��^�֤O��(͖-	i��h�k�a��$jl�#�9u����v� dp�֐�dZ$������Zy{�j\��+��M�Q]U����\z��A24w�
i�^�^�?.��-0���5�vļ�����uEI�:%C���$�}p�W(�s�`����BD��9a��o��$m�l1ˑ�mS���p5>��s��W�_¶�"��`/����_h<�6����Cp�&��r�р������Ѫ�'
E.;u�~W�B,�Ï1&֭l/f8�X2&SUwи��aXa�G:�X��S ��(r�3���iX�aM8���=�	��[�Yf�w�|���"���}���&+�7#b�@���C^`��O�i9WO��M�ک�O��������;a��E�ݛ%I43���� �C��Vm����/I��6��(݁Nu�"�Π��}���<{�Y��ʆ��mdEKd�.8&ӛ�	ES�]��f����f=�������\�v1�Ef�o�$�hNe�RB��9v;.l��۟���"�b�������ݶ_�WHǡ"=�L�H�_��-(��f�+�2���hՇ$ظ"#|=�-���I�3�Un��_2ȼuE�I���2Z�� rgD�+4�|qҨMq��Q5�R& V��R�����$若u"���U�$2У�>�Q=8M�!�Ұ�t�I��Kxh˱.�!��X$�y�Y��=�)�T�|�x�H���R;� ���e[���zD�9���i.�xv��1���j����BbwcnZ8��qiC����s� FR�D��aJ[]"*�f�f�JqdL?�����X�������\��[�����Q��0UҜ�j�:7�K����I����w��%Z��Nm���v{��#u8��&Ǩ����t �yyV��K/������cG9ٔ��"p
�nG��Q�3�@�l-#��'�0��]%��y����)0Y����K�ĕ�_��*�n�?��VU\�뱏�:g��R�Y��� ����2�gf���ٛ<�h�
ݓ�f.U'�5:+���F�!���\("��\ԧxz��#4F��~J8{���ps��s}w
�є�E<�,�R\tU�N Z�9~�R["��=���T$.�`��Ի��n�Y�1�C�����3 d#U��f���C��M�%[�f|���vi�gx��Q���B�t�4k�ѿ��7j;�;֝ϼ�Kr9]��?��Kh�~D�'pa�pQǷ1���'|�]���Ӡ����-@D5�����{Y=5���L�G��b��0i��!6��X�{L�y�I��o��2���1hx�/{�Y���hi�fE�HF��*y���"�Na��=�5U��]S:�C1Y���:7j�	�	A5�F�4�����WB�eݩ���b ǜ��w|��UU�v�ݽ�tѲ��Ž}$�6]pJ�ϸR�a���,�1T˯,}g���&��C��h ���K���׌/�b�������\ �Cl��!șY����B�8P؅��&c��Ǝ�������&�ќT)Χ=��8��I��O,�k��9��~sm���8��Z-�@���Bs���Z�T���t@13Hr,R?J��'�dt�o�7�Vt؍S���u�S6��=�B6>@\	�y75-���j�6�u2�_)!(�����_6�0��y�>�1��Em�������6���$G>�80��·#a,�K��<*�ī�Ճ /�z�����F��P	����z��Sh�yB�1<����{���3㰽8��^�>	a��B���Z�����u	ߒr�9ߚ�z%�IF��UuۆU5A��e��P�m�,h��)&\'���`�h����4�qH�N�`�ª;�}��*����A/�P2´j�K�>q 1>b���F%ؿv�T���-�1�b��3�I�Y�[8���-��g߭�N�X٢���'���2�u~љEȘ3V�	�3�V���߽n2�,�(țG\��ɉ7�]0�E�����R����
*�i�3����P�?�0$)LzV��2//Q�ә�)m@���m:��8`���
 �KqW�8,����(��h�݆��/�2 �2:�{��:�6���T�f����J$���a�'�I����·9�J��_ke��M���"�@��1���~6�$0��)�kH�m"��oy�	Dh����uwm�1�:@�x(�.;y|A
��ϓ�l(��M�b�Z��kBZX��Y��+�^��-#��C�9��ϝ 
LK��3�F���͕���.�W�gJ��+�j�S� �bR=sy�g�2���V��Nx���"Mz<�wi�����L��
�U�ݽ�jD�4Ky"�+p�sl��E>Oo��s-��v���3��R��G�v����-��	}2���#���Ҩ�����_'H�X<i��W3x�~��}v�o�\�;������rՓߥN��53 ò�is��֤u�=�w�:�M���P�c��r9�f�=��E�;�F��*�O�'�+1��7?97��-�Cf�fQ�zȀ���d�u�f.��Q�6�y�7H�gɝL4�/�ls�b�su\)_\'��@�j�h��nĲk��DΚ����_U7�Gʭw3&�~�m���򐗿a�4�����9<���m�5O\��Kh	``:���_��-W!NY�D����E~ӱ����Ί�2�=O��OYj�p+I�}q?*���y&>��T�����r"b�ʏ��0�����jUHu��j��xEK����
��v�Ɔ��N���}a�������l�i�M:���D������K��#����*�����o��;�p?hb����i$'�TL�<�[�/��MVBb.�{(ny/�'���N9p�  v�H���y9e��<}.�ғ��9��AoX�a5~&v|l���FH5�u�=<��� n�'eC�'j�;$/T*&v�\�OQ�ɺ"�I}D��N;Z`)"���I٦<Cҙ�@�~��{D�� ���{{Ԧ"���eQ�6�e�X��<��F�wQn"-�ų�)T�k��� �>p�G�ل�w��q\N*��>��`�rVp�t�=��Tj�z�<�)nbӾ�oɍ1�^ �|�+tB��������7Ύ�'�P8�v��-�}?|
z� LT���*��!UQ�3��윒<���$9����\P���zg�EvZ����� `�6�7.�5�(v�Q���������j�-��&��{"p$�x��v�J��:�V+����Mq�d�_���;V��#�"�'�-t�(�� ��+���}����N�EZ.,�˞-�z�������A��Z��d�r���川�ۋ������=C��{-9G�H�ag�X�9���x��#Com����"��M�Ei�S�Ѱw�LᐴQTcpA%��^���z=9C^��A��bDH�����EaI)�n`ퟜ^��;���w���Ġ#���6��i<sv���"}`��`�u��I�:v��ƨ�1��8���֌������d��s�F�����pP%��`�
I��|�3̻3�%c��(���f��+g�(���:�O:a�}w���]][����-�_H�_Co}��P�$z}%��v��^~? %���D���~8S���]�M��Gg� C�~ȽYI�`!��LVE+����qUH�D(a}@f��+(��R�4Ʀ��Ѱ `����@'�FJV\�/��@�Oq����*�����䮯�Wi���LeG6 x��}�u��U�zb!�װ���8��1>28�C�����w���r�4�]]�f\�ޅ�����k�����'͂U��>M���&�8u�&�Ė�����o�:rA-�y_�`�g��I����:0@�;���[#aDE>ٟ�r�ች0ҙG��2kU���`dO���s�C���s�%��3��|Ѣ��s�'�J?���ᖷ�3����O>��F�9�طsw����i!��Ծjۉ��'�����;��tI~O�H��-�r%'��e�r��@]���r�XwTC
.�ee�"|3��6z���#�dgN �/���%����paA񢏼J9B;��<q���їS`�s��hv۴͖�5�᧵y����@"C"�ZQ r����Oz�5Q�����6����h9�̯3��P�*E�8��G�O����������%E����@����*��d�����5����g��e�3�| E��߉�W�M���%պ���H�T�8��:���8�*,��d�f��<C=��z�G��k��oq
	�H�=̒[Q�����~CԖb�o���	�`b7e?�����	��W�Xn��'1V��VX�1w��!��ԶL9H����9��G�Zx~���s�=ŕ��jvF�� �E��	 ¼$CH��QZ�8.�5��Bt(�58��|�������ۉ�����@/���K9���0���� ^�K�Q��iJ�8��k�}-��<���l�7N2���̐�@}��������.�?5��
TA���
�Pe��8#�3��s��[19��&;��=m�8I��z�b#�fִ��C<gOC�즟L�ϛ��`�ʴ�4-OUtKӭ�Kl*�Z�:C}H*��tI ��/0f�@K�Q;9�J�J3���w�Y��c!Y�SM�n&b\C�雰�NNiz��q���}y	����A��ru���O� ���C�n���镏�򤘳p@��%�d�O�����T&ƾ���-���!wE��}�����F2�k-�6<R�Mwsf��Cx(�=�p�G�K6v���4l�v�����U�=�A=A�O�(J�;��di��(����rQ���<*`a}�_lD�Z����� �и�A�2a�uJ��9�j� �3
]�8
���`��c�R�+I�a�GG�<3Z��Ɂ���
�X��Đ��:��X���V
�r��OOF��f��uȵ��F��^BjvG�#2y�&3�� T����0�̗[V��i-z~����p��3��|���� )-�{!V��
��3�H�/{��7�ۦ�c{o���u��������ֹ���d߃�Cw܂��oP�K��d8�S�0��&���)c��KBe��z\�o�m�}/��'wq��ү��ՆOvhyA��Ea1<�Wk���A�3��l�H焪�_J��V`�'��l�FSLC$ё�.��y9�Z���)M�����nS2J&.�VL}41������f��%,'H�B!�*L�0˒��3�i7����b[PR��	���B?�P�=�_x��⓫~q�׏iLԹ'Se*�^�%�OC�����hc�����B�&8��g!dɾX�N�Kc����'
�>�U/Pj=� ���&
���ӟ��q�D��驶z���K�BK�e�J�S�.c�Q��G䥰!�W��3��@���	 a�8�ӣ����7�)PƻíK�b����m�l����Iŋx�:��U�-��@ʩ�H�	I,op�~�R�	 (�G2� ����h����Al��Wr����G9�l�N�� �_��bz�)$72n��DG'
��k��@�:�^V�8�]�'�C�U�?��͢���ƯNa�ĩj#��L�K6���t?�z�D�ڕ��'K-IJC�!˦���G�l��b:�N�7�x� �^ґ}��!��)�<-�/F��|:剧�$u��:>��M���]�4�l�ἁ���~�n��V)�&K�dz?��xlNu�ʦ�8��9\u�ь��~D�y�ju^�`$��j�?�i.tu(��p�+,@�5��+ Vݛ<0��SV�;�K�eV���q0�u��,!*�Vď
�2�p�������4�)�I� n3�'B}�B�d�=`����hzi�&9��V���<M�w�>E1Tc�#���)�^�M5G���P�GpAܑ
�GZ������z\�&�qB״���"C�����2Q�� "����<����&х�y�)9$� QGǓ�	�
���P�*��������|�|�c3��w���י��cu-m�ݓ�իSX�7�aL��͓��)��Z6��(��ˮ5�v���P�ܴQ��#o��
2N���UZ���>.�(����Aڋ��VG���*����_Ru��M�*�7������i��9$�oѶ�^����Y.i�������c	���p� �Ƴ�~AH&ȵ񑸿T.Wt�5� �4��9O�+�qÐl_�vhn�����'ʦLJ�e�#U{߽���\���W���N����v�QU��U�"����J�{�G�=���3�& �A���x�y|O�r�;#Y?|6P:h�h����F�vz�e�~o"��M��PS-D����3f���0 ��gՕ f]d{֚�3 �Yt����Ԑ���&06%I*�3��\uE���I���?V�q-��G^,�UD��a�LK#����k�D0����p�J�_8����a��D�`�԰g�nU��e��5�u���?m�־�2����D�����z���qf��7��3)�m�������BHw_N⃮'�4��Y��ߣE.	��iI_WM�w,
BH��S\�~�m1˒>^#�4~�4�>y�}���Q��]������M�c����`"qE�AA�q�6.��̉���=�)����s�WoeA�����I�b�`\�T��~K#��a���ʼ��`����n(�%�������0GZ��s�1-N��L<���Pc�>��:��/��o�z�UOz$k��8#R`����g�O9��W�sOc�����#T�8��$K�>���ϰ�尢=����Co������e#9M|�*�E���-\�<#�m�:L6��L_����Fr���{Z3j��o�@I$��sl��/��F����2��R��ADk�^W�|��H��e�IvB�@R��@�K ���<���*�8Ʈ<��(�
Ed����������{����ۛJ�p� g9��� d`��B�M��{���Z!hl�;�5�m���(�����t���um���A$[��Q����^C �2� �3���)����mup�5(dn�X,��� m�)��./�0J���.<����"juD��U�H���In�P=(NDO�͉��3A~��J�c�%��t;�z�A(���-�ٺ1���n�o̝�;?g}\��F?8}�容�aUj�lC#N�M�7'q\?��B��u[1VM4gy���u3ܭ�T�ybM�0��/�>юlX�;�E;930���T�������ӰG�>�Gǜ�&�vY�&-�]�ڶ:���7��]yU���=�By��7_ps����eTC�$L�VZ�03Q�(9Vq x���:����/Y�+T�8���C���Y�dJK�rO/�������zTҬRz�d����2�{+�W�u��$%!Ҙ�9��1y�9,�V�ÚmQ/���r�r����6r�d�l88a�ace�%�g��ֈt:aX�;�\V�����)׶Dn�f L|����H�yP�!��%�,Ȣ�i�p�BqOM�a#�
�G��������hW�k����v�`���vo��+��H�B�#��I�cj#�ۖ�i���ɥ��jg�~�3� !��)�˻eۋW�9���:A���Va�~�+���闵*���UV��	O���m�;�3�6�c��K?��К�gafL:��-뿴@�D�@�ʐ��~/��&ΏL2�R�fZ��(P����N�#d��p���k���|J$��N���-<l��ʂ���y#-"� �d���37��ފ�w�[���YV��ik���S�eT��L�=���EC�k�&������#z�+ư��dP�6ō�h>z��kp>�ce�+C�q���(Ldx�L���^�����#�]6�����)�TI(���>�$���1ٵ�p��tQ �(O��kU�E��l8���	����$'	�����"�V,r�T^�M5��J*���T]�;5SJÁ�m.}j���{0te&'�0(\�mBz���@�� ��p��h�i.Ay-y�$�jo@Q԰pkӄ������g��+���|���?��ܸ�fOd�N���
�M}���Mw-Z񴌳K�1o�0�ˌ�ȵ`j��<��1���� C5��sG����/���F�2�b�׬�/�*�5�h0��0��KIo��̓�����*g��̪1��t������g��1~�G���h{�':wd\#����Ă�(���Л�_�����j�X�ۣ>h@A=f�� B�Y�	�C����T�fؙ�=����`�a赒��;I�0ZpzZG�+����ڽ��h�"�eV'vRQx���W�./�r�ˀo �	��>�	^U�ٶ�ZZPR5�&����C�H��6�����	����Ň�a�-�:�S5U���0���	��v&=\���*���z��K�e�Y�,�c��yC3�ٴ�V���60Yt���f�H������Ƽ?�.B��V˾a�[����q���ɀ�֓�4�`Zzi���^�U����ip����)TW�' ���z��'*�<�_�̶�N��g�O��3��-����G9Bt_�`��Xl�Kʪ�<ֆ�S:���}��z�SG�������x��Ϗz�#@����E��,Qz&/_1�RNy�l�`�0���@�e8V��)���B^��D������.�x��&�x-,���S�V"@���#����"�OgS��L��+�ko�{��_��X.@����u��]ylЯR�Іa4랝ֱ_�|B�ĝ�õ�N�/E�0��U�j�����o\k���2	��`S�ˤ��'Z���Hq������?8(�G�3��ȶ��P`Wڊ�=�V_�q�(N
$:F�����Ǡp[Y��>C��i��h��g��~�ݬ�"D�0,_�!��\ï��tI��x�����"�
�v��>Ɠ�F�H%�3�x�%�R�u�q���4J�Gǳ){��/��:�A�f���܏G.W-�r��O߶]�����W�J7�kz�ѳ����±J����v�-��7��0�9��P�k܉-���iE����`��< �������d�6� �U��������_�".�C]I��wb�ݶ&P�כֿ����C����"�j�
�],��z #~��RLa�\t���[S̀l�����P��`���`}�X)ߌB�����f�c�Gf
��[?�ЋI
wN#[�/��!������6�I�] ��mk��E!j;��� ��=��hٱ�h����a'Vr�k���}�!��Jk˅z��V��q>�۔�G���c���ێ�H@%[�NY�F8;�!z��/.j���9t�y�D�%�`���I�?��֥j��~	����\����,�~���� t0P+*@	��c^��� P�/'�Vc����ѷ���EtW��0�ɬ��>�����X�1�B�pjw�����~����@�Zg<���ф�t�*��D�B��)��4pq�O����6�^p��]8�J8I�,�g1/��O��/t��'�>��2�V�{��/�k�윙iդe�ؖvA�@��_~bm���tG�ydG���c�_!vu@��?1���k��Z�D����W�/�(�t5=�); x�Ro0?o�٤ƶZj��K�@�.wa8�A�a�@j�6^��3"J����LR?:9�k�p�`���ns�Y�|S�}��˗��ڲ[t��x4J��R������6�pۙ}e�7�v�Ƿ=]-���(����$pK-���k%�S�Q���B�e�h�b�I�_g�>Zf��6Y�l	��TS�"?�dg�;��U5|^/���D�f�FY/K�U�I;��!x,�R`�Ѥw�/K��_��������C� ���{����dy^a��� �I(��H8��GD�ۏL#��6�-�?E���$��}{��L�Ɩ�d�I���p�e�g��f��|�Z���'�]3�����T�Cա��d3��J�c^��S����?���J����/= �)��-��S����{eXXn����B%�M���5qv��R���ȥ;��Ga�X�1B��� |v�B�h�M��"V�,J��]�m+���b{��u���$����M07/*��P4�o��H/��U�o3�����ҵ{x��ֳ�g�f|fmX��4�9k[��i���_�j�_��q�{�:8�Z#�^���;H�1�����ڦ�,,>� ���\�Ȏ�㦚��Od�k�*˜�i�x}�ц&�����.�4�������8:H�Є�Hņ�} �-o�
�����`�.C��a�Ź�!���4��PF�Q��$�|��H���L�Ը��a�pݥ0�#fH ��3�'S� Z����\<���1�{�h�JhŖ�����=���q=���Bh���@���` ޤ]a�V<X�&�����W�թ�p>8�(
�V����ԃG�R ���TS��^�Ӟ:�:�,�����1KI^��*�Z����3N3� ��l�A��,�ё����c�����m���wA�݊�N9h�}(ؾ�B�xK�o�b9����!���%K�231�)1�D�ч���~!X�#�]�lD�-��W�s-	���L��q�K<�)�~��X��WU�"��ˁPAz=�}{a G�U�"�P}�0d˺��c�/L��|�[�7w��5����(ˍ��-�J�	A(��$qŨ��_Ni� A?
�O��?��Y7$THt]c(�*�K.y�p6�-�H��l��F�=�SSP��D��>ʰ��b��dPg����ru���{k��O�v9��ͭ&ڢ�A��o�廤R��.�}q{跱�{��b{;6�Տ�E�S�x�٣?q�M/��p��>����P��!�%BIm���e�#/1yV�z��!��Z_b8�~[q`٭�t�!C�Gf!6�(�2'J
���{��	�\�"KM!١�I�έ�`��MhР�T3�7 \<X�4m�ޢ�ٲ;nL0ѧ��E�S��-7Uġ����U(Ap����<_]uV�	��������Cef��@	�,a�m�Q����\��{Ʌ �{K�N�2 �RS@;SK��A,�p(�rpts	��7�S���+�uR1GE-|��A��ܚhF��௝Ly���0���k����B21��:�)�U!P�:�"�_Ì���y�C7G7��ު��P�<�n[ޑ�e����HT 9(5^�aԻ7"���$(SPbӖ�j��#�<�ې0kpw�K*���I��3*�E*e5â���տ(�p��X��������l&*t�ݕ�ڟ�����T#��9B^-�W�)t��|JD�;og$�#����)��=j�v�� ����r�6�|q��쀽WaIy`�1�~���]L=�pH�ʼZ�f:��
0����.�V`hE_��^��I @�9KΓ�.�X��g|o f0�U���?0��\�v�1��amg��0��ܬm5}�m���Q�F�2�?F�ⳣ9���VA5�{3��g��\��+f	Ԋ_��
�W��0F�2���1J��`���g��%з�o��h�
Py�5g(S�R?�]�%��j`bJ�|�C\�l� l�s�ۘSL��J� �*�%P����tSKy+��Ь\C~/q?���-���,���H���⃳�J>�cL����C��7^�թ
dm
5��^n������O�\]���.��`��|�o�ҭU9��m���*��1,��yr�=j��,���1�����lGˎ�	���Ͼl�;F���ʔ�I�G��)�P|g�{x(Z�4`V�v^]s�+ҏ�����"������!��w���M�\�;�K/+i�G_��$|j�]"B`������9:�J(T�+�w+���P\������}O�Z}0�X�3\^�I��;|�CCPZ?�`����ؼFr,�h�S���!
A��?�7%	a��.'h�Qm���:���n�(���W�'�[�Sc=����$xP�^�F�:?�p���[��u�������Z��<�������[K��)�hW;��i^n�W�MGE���7�W^�H\ns)�t�~!���K&a{啴��ခ8��p����/�&�wX ��ۺ��%Q#���t��e]���I����k$�H1�zO��*��+����Ū�QEBߺ��Y�5�c�D(��p;ǘxMl�{z����'�sժ��nļ����ǘ�ӭ�8���[a���i3(ouSRO��r�UEZ6E�j�8Z=4dQ��}"<�g¥~9��l�:��O~TlE�b��83��������Y`�-�����	�{�A�o���2�D��14:�j�nI��ț<Չ܍j~�N��X���[jv�f[��m��^'.S=V�=*JC�a&�q�%�˂9�@�8	QoQ����!�U&jSu��2`�q�+��Ϳ?M�qt�Hu����5'���n����&Ζ/?�
ц�7�8w�O�Mr�C3݌y�cB��	3��=�1����9.\�?�:���.-п/��+�T�7��Zx��w�|�=9�������mួZN�<.��~��%ew1��f�D�c�8N��l��f��O@M�ݞ��~�K�d��$D"��u[;1����L5�͜����x5˖)����D]_�]���A.�L���Z*>;Y��|�b�@���|���T�PݸE�&�K��ݴ�������F;[���T�udO�?5i�ʷ���G>����e�(�e�<iQv>�������nh���st0���g P���F��g�����O�$VlC!�4�.7�?ɳ��G�S���~���=s
)H��\���Pfs��}�3�#��/HQv�qB,�P칙�h��G8�7��KZ֊(w���d���BZ������[��}H�NjP4����ý;g����6��<\�����7�0���ϩc,x�^�A��K	��n��}����'�_��sX�m���/'RTt��$�L��Fp����f���ymj!��OV�+��7�}
�Z>���jf�K���q�8�����*�	+�oЉK�B�c��i(ܴ�r� ���$d�ܚF��x����}�WD��K�q�甾an�d��k!oz�lv�:'����B���b����q�p<ئ.����l����Db~c!DN8�߾��|+"��9*!k��������s#K=��IO��˳��R�>���P:�v�L-�o���(��	XF��[�K{��'����q�m�BM�.�5sVk�ʥ]��^&��b�$kZ�v����=:1�s Jp�g��=��t�@cw\��wZ�LNv���&�P!���6�K��	�-"�zQ|ΰ�W��A�N����׮a��*ZX�Uw@���^7{�h���R`��Q~���1�ȳ #�%^�\�O;�ׁ��i��x^���*�4�d�U��Q�_��C7��D��l<��PH���]PƓ� !��l�k�ĸ��Y��O�A)�V��L~�ΘI��<s��raԢV~&i�$W�hzi�霷t.����;��h/F&qj��PS1�/km�Y۫*��p�N���BU2w.���p�=��R�%4p8ґI� ^�b]A�W!L���	_�}��$�;�� �*yH��j_�.����.bf`�������,Cy�Y�j0��:�YKFv�U�A��j*�n6���U���\j�D �vi;�<e�V�D�*O�[%�2�NZl٪M�8Ͱ�	�:k�w��X.¬7T��ڦ!�d�#�%0����[AM���m�at���_�:��6�o��g��LT/�Ft�a ٰ������ƈ�_P��W^,��:M���+��{HO�w8��)�%R0�Z;") O�Ġ#�׸0��b�~ܖW�5�nC�KP���iy) �qwr[�d�P_�8�.%�S^ZK�*;h�z�r��-f�d2P��d�b��VcG��ر��y�Idw�[Y���up06����R?� 	���Jl@f/�����5�0R�*���&k�y�)\ ߏ6�G�(�����d���U�=</P|ɕ��`������o-;%�Ș<m��V�0?�Ozʴ�!��F����Wu�9� UV��[@���,.��&F����A*� Y������T	?�^��f���F�UOEq����g�����vV-�\�۩�x���'�>��INE���Ŀ��\ө��n=�o�����n�E�l�Oj�G�]�i��pSEm�VY#�9赳wY<|fk����c����K�Cf�S���;�k Dj�*[�r8P��}n�����J�-پ�}r/���y@0m'���5�"|��1�S�z�kfY�a��X!a��6uh^1�k�ؖ!O�|	� t�M4��V�ihf���-ђ�p��`�} 	*�>,sCLn-)0f__q[�צko��a7�nr��./�)Њ���iY6�)w�J0�%��W@<b!임6�7��ͯ�����I�ŮK5�"�pN	�.Ę �|~��Y%��܎~��l���R���נ���}�j#���닀��;�ًF��mM�>�kgW�3�1�Y����3����߽�嬧���6Azp��%"������3iƆ��H@�&`4m���l4�w��|�s��C'ۯ��gVd�f�]AL��� �#����R�tz80�u&Pa����	��O,*e����m)�|��)�1c7�LaN����ʅz�I�&�����ƽs=д�nNߥ���/�wb�}Y F�g�02���f�{�Eg5#��=��|�g�*�X�oρ5.��37s�d���/1eB�g� �/�JGSVp������I6B%>6S�6��`؊o1�1w�nx�<���_g��p1#��{�P��s�<����3�j;��L��[��4�b�C��I�j0�!+��9E:�E�|H'�:S~������]4X�M!�㔼�N����N�$�;�T��U���o���
�D�?��Kf���Vm�i�t]u*���jx�7,ɐ�����\���Z��m�?��V���ıy:���5���pr�jʑg��ۭ��=g����ǨJ.0��r�K�����w�'�P�.�	H7_䗥%�7!%�J�t*�2P��wT����1Ǟkpx�OGd08l͙7tܰN7Z2�ɀ��Aj�-�yN�����3�Yg���?�"�Cs����h]i�2B4�hx��M�oƇh�:�2����� :���:(��D��f�ڊ���7�T�$&�b��L8��v1���YF���R��x���m�,V��W��#�7*�iv�HB)Z3Bо���T\���Q�l�������5 P�=�}�.�YW,��'��M/�Ty\֍�#��� s�;�YΡ20!�@#�{�H��O0b��l�ԵA��k�� x��/C�����< L�H9E`Tٟ�'���1�`}g]�:�"3m�I-Z����UJ���;	t��]�d�/֐�U�^[k4�2ȑ(�嗞��8/���_��,�3�p�s� �6�b�K;cؓә^�����+�3%�zeW��hr�/L�q�o�d��ἳ�ꛋ��k*��YoR�|u���mb���Ld-� �\
�n]������`l��Y�o���d����f�fQ���乳�؍7���i��1�h�-'+�7�߯����N':4��Əu[�[BSף*y��h���mQ�L���c#A!z�h�-��G
�#���{�϶���Y�"g��F݉A�r�_�/ƴ�� |~�mCD�p�QHT����j[��
Go����
�Nwr(%�����yHJ�4�)G�Q�4^���W�7�c���zc�}����{�K�w����0&?XHC'���p�41���'K>�ʌ�Ʈ�Ԉ"N[4W�2���)^�����I�;ay,^��gY(��1"��m�ܬ��#���@�v�C�t�Ԃ���(&��8��	n��a��4'�y���ݽ���+;6����[�q��a��������9iG�T?^�XG��!E��5���o��⪕Y��.Qژ�/7'�M�,��Ե�UU!ps�P���J�8V�9�Y�-�p%W�^+w{�O����x���"CAGQS?�L�e����g��E�� �bd���'p��,��Ja7��ӕ%lF��q&y�)[�z�z=���|ztu{��^�]$u�C�����@(�.�7g.Z�GE�%��b�x��u�EP#�<ܒ0C�VٔP�ԟ����ut�)yf]��7hn�8�wc4@#7�x���t<���m��Y"����b��u4��x��VU3��}D9�(�FP��н��ܥuB��f�.m�`nȞG����Ey3����Xh�#=-n^��5u�O��+�0a�ӯ�+5Eee�@�R"�惕<Q,X�8m�8���������-�1�(��6�K��m�KQ���U�I_ם����MU�K�#��w�j٩��JR㳭d���<�.oi&�BVq��.��k���i�x276کC��V3��zV�<V�2i	! �s�>Ǚ�9M*S`L���2KC&"�<#��*�K/�ܾrA��fM���UvD��j�ٵBQ���OR�,��BO���
گ}�t�UL< � �͇ұwYUU�d�F[Ɏ%� ��	L"��iRN�4������]HNY�p�@~#k���.5Z��=:�*�oh��v����$�F`���qQ�э������{?!�B�l_��C�:}VX	�����ڲ�������-�v�4r�q�}�@�q�;A�P�+��et�E|N��X����bX��K��/X�|5w�F���Lˤ6_�:8�jw*�q��85_	Hʡ)C���H�C�P�+�����%b�%�Q��,:�5mnj�����2��� ��UFG4A
,���o�zJ�@B�B���[&��T����b����x�<��Xn0s�p��	f�����*3�/��D?�Z"-a��c~j�T�ڛ*_x�A�.E�j�Gޓ|����~S�ݔ��>\�j�3��}s;s	.���.I�Ko�/*]�c�c,�}6�V�9#�BN�Z�Z�	ͳ��JeGmݸj�t�JW�k�/W�H03�~y�gfB�UV�X��kG����[�I\���\�6��# �$lM>'LyJZ��[/��Կ/a��U����s�W��ץl����{8�R��
��_X:p�m�I�2!KI�yX�'3B�����I�|4��6<w��B#�a9[L�-~kLW��Wf���N(87���>���3UCl�Ϋ�\���vmf_]��>nf��W4��Æ�ITY���P	�ݶO�)o+&����甎� ��ǡ��N�������fD�Z�ĸ��׳2�f��^~$�v MAL���ʱ�oTT;���읅q�B�3��Z.���z��Q��rq���K0מ��x'JJn�o�o��p����#B�Xk -�6����z��68�B*?�h)k��y��8�f�<THs��$+\�`�Lx�f���L/���vˮ����	���=��Ob�u(��V43�����^,"fW��Pd���vdu��K���;O��}d�@~\0�*��^�a�K�'n9�� .w���x�|�+�OB�NR���k��E���<C3����W'Г�
 UY`%���X<��I(4�~i�{9=(���I�\�;i���Z� �0e��>���D�u��A��~9��1�=�V�!+%Ӭ��4��W�z��^���@����(_'T����]tk[]��jM�/<�˴8Z<�B��� WDݸpw!��ضVw�]&��[�JcO��I�jV�C��{�֌��`u{���3��&Lm;;�m�f�K'+�A���s��r���V� |�_/O�9�)��/�w;O���'�(���y)�9�ѐ�UE�W�a��0�dv6�{��ewI���Vދ a�m��UQ�}Ca�J�(�b�Ǚ����/�V��:%f�UgI4��>���1X��!��j$~�H�4jg�$�����#(w�9q$A�[V�7�KisJ��ع�=.pl���,���H��M��Ƥ�Oa*{r\��{��ԟ�V���%�q�w�42�qi9�+Jkfۻ+f��i냩z� ѣ��CX�c����a�9��I�Z�0���������^��?-��bd��K�T@a�SRWZ)[�81_�X��6=�����z���7�s����M�|�:J��x?||�`�Q���s�ƛ\sgVY��s�>�le���4�J#�=v����_U�\KX �O^O�i�Z0��"��$���6g�ZzL���d��A�����^�q7f+�7�3�%2~&Ȫ�(!�O�6�цY���J�~'!��{l�|[�"!�\|���V�Q$�����Ԝ1���T	g�	y�Q���&�ȭ��ȊL�ꈫ�IyM�!�k:Jt��1���]���ĪjB`�������&X�KC�<��7Cq���sp�b�Ǩ/#Q�U��cO�.�7rW��V_M�X�l�0��)�K���j� �&98
z@����.����T/��\G���BGn�PCDl����"/�I���(��ߎN�#9�)�P��p$1>��׏Nx0b�(�]AR�G�y%�����"���7^Pk�����Lؖ���{D��t-�d��/6-݂s��~�Od��5�g@6�`������.�W���l��pنH��Y$}^��Gg]��3ղ�g3�b
�@���%�B�:���m�D#��g˳6s{W��Ց}�uS���t�x?^�a.F��]��e(��=򧑲r�- �5��X£;-c�}�V�#W*b僉�5ɬ�꿦�V4�v&���"�Q��Y=�X�U�}&�V�����+�������Dl�s�M�����:	�uy������@y��V6`k���R���z�<P�<|��nډQd��7�U����|��01�h��ɛ�L�[DU}Ml {�d�Yi��6g4�ٲ�~��1�,�����s�NR�.�-)��|p*
���N���ؖ����b�SI]�]\V"�k���z��v�(���n�?�=����WJY�� FGͤ�|��"�������6���c��Xްy0aP��ce-̉����8�`�^��O��>n>z2��
�ڹ�iVr��qx#�f*NSv��0��2�5�����f��<��@"� =��)"į$���bS�_63~`*������L� �Z��!�*s�>�p3?z����R4���v��-��9 N��Ȇ�!�P��� �@��*�E�����Ed�G��.�+�^Ni�w��C>�1�ۉ�W��+X��-�2
��Y��p9�Mk�y��4��bⱄ[��3��$��g��+�[���"��=Z" aD�b��������_�4Å��}�kɐD��;�V����9A���	�ѧqv����E8��]�8�{kB]�56eD3' �
�*8̙�	-'p�Zc<B�6굯Y3��!��+g���7$n��cB�xI9��[�d^�gP��a�_�x�{�����T_�a!'")�iL�6>`��H\C���L��>�'�ٌ2�8>�&��m��ʋϞ��������bD96�9_?~�I�.v���vb�s�,���ԪŸW8ǐ��:|u0��,�f��r���-��*4V�:�vz[~�-��6�2=H&�i��A��n��Rv�*��ϡ�b�=��S� �"��{�~lo:�{���/��R���.A»Ԇu�>��y��' ȕ-�͕n��Z{��XU�G~	'�d t��&�j?ߡK�vĔ�P���K(�ػ��ނ�9V�V<^Acu݉���$d
C_�k�o�;VR_8�I��9۶��BJ��4�'�R=���{A�D<�*�e��h
�����#�7��{fJ; xY����3�o�q�j�`x��c��`L�O;��:�0}5l��+z}7��RN,�q`!��J�Ξ���œ2�^�U�x���eSƚ��\6�@]�2��pI���&��
��MX�܅�%��ш!�K�kWR_�{���dԩ�r�#e�`f�Ua���Yx�~����Y��������Q��D^|��Y�S�`p�mhJ�$	��I�H(����n����lڝ�R��/E��KAsmS���e4CT�,�;�����M���-�%�<G��>���4O�EE�p�.��$��؈��K�~2u�H�0�	\ҷ
I �ʀ^y�`�J��󉊏i ľ��2�������Jܴt9�S&��|RL4`%\��Q�as��Y7B�(�X��+��j<j�$07���:J����I����F�>{&��BC)Xԧ��A�9V���gK����}��6/�WL�[���P_��8ʜ�ra�z�O�Ӂ��5���Z�{�K��e��з״B� 7�p&|'�d�SN�>Z�z�T��nۍ��a��>��d�$4��q�>Y<g{�}33N�D¯�ٰ�j(v�]�y)�ޟ�����KL�H�	����'�WNo`kȫeO��m��~.��jU��Ow�ѵTE�7�-��m#��{���_��̫P�]�n��)b���̏3~D�@.����<�9wӽ���=vS�i��B���lI��GR�b�����>��3 �ͭH+�8��=0'�i�b*�n+�ҕ眴 ����Y�o���%F��򣵧	A^ n�`tE$�o��R>�e3[l�0�~g�h<�(|�3�����x��5s��6]g���%l3;$铺��pE�G0Y��L@�D���5C
��k$ߤ��0�\�w��(W�F�M���q��ei��>�����Q	Y�l�N��-�#k�b�+��Í��w3A�>X��'.� W@�(g >��pw��@ѵ��8�r���g9��2y���v�}Z���������ĲJ�i�;p"�:�Jy9�h|jJ;���5I��u�a�M�J�v�k,�.G$Q#͘0��p �` 1�5���19
�Be�����Nt��(\�����%t$� ij����K���I���5L�[!����^�KI#���z�'���t��\eɢ\ԏ/*Ý�'���O��Q��7Y|'��r��qh=��0$��S���M2�A����r��17j�tЪ�E����\Մ<�d�c�:%�$�>����[*��F��A/�{��s����(@_���Ad<D�X�d�:V~�8��W��]_�����2k���������~^�����º�71M�$Q-Gx�W(��M�7��@r�ō���ig�E%Ԩ��ֱ0ۼ�B�}^��O�}!��m�����k` 4.��]�Ȁ��[J4N0ֶ����jBJu�V��ʊ��3��0%ĩd�v�W��gT�%��0 ��A��":tHi�[�Xl�2�\m�AnU�+9��T�U�+M'���>��������q�fu{�dv��������񺂆WI	� OsL7a�|�"��f*]�q�7���w��y�N��v�&f�u�vM����0hij��[p5Ł$$����� �_��ұ���s˸#Ί̀'	"��ϟ�6�P��2��ܝM_ �m���(6bU�+"�#[|�U���V:������.��#K���U26=�%Gك6ځ�5����=T�V�<f�������h���st�b�,4ϥ,�ˣ�ċ���Φ�{����ig��4��3	���@]�n��Z��4�j	�@e�^�0J۪[��K�[������;i���7!89c��A�孃�����ŋ������o�;3�q�� ��m���k�THn�2�9���3���xo)N��H��$Jw����29qU\,��"����䋯Kj�X]��N���~Ԇ˗�gm����׋,��@�B
%��k�?��2P�<�uR�y�*��yp|�L���� � ��������qa��}�#�[e'ڮ�c�T��w}&a�|�b%ÖO�nt�Kq���B:Ie���[�J�D�ڍg�����(��ݝ��yғ�kt �P���U�;vo�sܖ �(s�wV� ��/����a�<��Ow�E��$��t�Fq�O.()d���v�l$@�l1��w�r�;�C�*�Us�,�H�lh��=zQ*�~h)��m�:7�'�X�:�E�V�Q�������WP�<\�S��>=:k=`6�P�[![]��w@)�bd�YF+�E����/`WkZ���QD�N�%ּD��7B~2Jӣ㼰x�_ΐ����� ���k��-u���{%�ݯ�]!B�;vԢ/S	^�)�oF.����2E^�*������M_��9jd����5ˇ�1��V��ĕ��y~c�t?SF�=�ҋ��{��o�%֖]���#S�1��qk�&�Oa51�����i����z~µ����\;�/�p�T.�4Y�3_A�'&;�J�F��������bg�h�	Ŗ��ߤK��
����`��pt��N�!1�p'D�#�@u�7LW���*-&=BO��6���۷A	'�3j0R]��@,�G�� �r4!�t��kE�h�O��V��=�sz���`�����G"���re.��$d<2�+_�t]?�LQ'"��=gg�츶+�A�7�z_UQ1�U���3��}�C]�� H�������	BxJʣ����?��Q|~{-[�� �g�}��37ߥO<�F�,dZ�Xi���_���;�Xe1�6"y ��v�V�)���3�0V��^�E����t��*�}�-a1�U��j��Lٔ�e�wڦ�߱�� $��q�E)do���\r���ǐF��xB�����F�t��Se�¨Ä�@���!\0�4DľUp"f^6ǚI/j��|�b���0��WvcQ��2�'k�M;�z9}G���ƆK���<�w+�,�����]�:ed	�j�O��,� ���p.�@��ڈ*!n5M�
|Q�^��ޚ�'���w�eb�K���_(�k��p��uE؛�@V.�e��Q�xK�g�pO��K�p\�������5����`���*�_�~C�+1���"��63�b<3Id���B�ZP�1����U�~�����kgB�1JS=h>E���_*> �ژ����]��C)�@c���d�lY��yg�JA�KƆ�k0�ɾ ���7?bX���~�s��2���Y��E���丈G��c
� ���>C��IL|�؎~)`�NY��M{Cq��ޟ�lo�aǆ�ۑ��*"̀�v�ԇ&��:��za�V�\��1bO���/j�b�P?��|��"h�����-�H�����mwru�� ����y>�3lU���F�����8��B�]g�O��u��m�,}ډ��ԭ�r�����?���֏e3���D ��j��A(EK�L�VY0��NQ�Z�V�V�:��n'�Rtj1(�%��" i	����>V��X�`Hހ/��4M��!���;g�ٿ�ؙH�J�\�ci_�N>J�������^��I#";��X泟�`{�yz<���Ԫ��/�[X�1��g;b�1c���$a�AwMee��a!Ƥ��\��~����1-� :gDM�;�Ё�lе#�(�Ie!��t�ob��Bn��e�FjiH�z�;o��N�L?�(�w�U�a�����VzEB�9���,��x�~�5�6��NB	�w>���i��Z��
!u�����Y�fJ�ׯ��ڄ���LA\�0�����G	�����B-?����y�Q��E����-*�0:M�q��J�('�m��;<V%j�y�#��ͪ�G�A��iz�?���):�R��.Dwpt=5kR�:(�"�ٯ��;j.x��}�̚c�����p��V�)���%Ӱ�!�2������ͯ�.E��o���Sm�������B�z�����"��l�唥�@[(cy�y5�3薹e{O�_�9a���lv=�&�#���Q#ο� .��e�*������W�H���A����jl��vMq��N���1�l;���~*�|����О�ȋM������b+T����1�F�YcE�B�
��yN����1�M��[Ñ/�W�����k�@�d-�w���k�!^VČU%P���s �^.(�#��N���l�"Ȭ�������{�)���)��A���Y���Q�����r'(B=2���5pKIZ����[$H޷��"YB�T	��Y-h��R��Pq6�-��s N�3c���c�4$���L��z8b��ϐ,�y��#q�6��(�����+����Kj
lZ�í��|�x.�IB�d1.�T�F
�f�ؚ(Uƨ7����p�h���7�s	�/j���V����u���uׁ;�i��A��m�9��п�:Tn��T�IsW��=�/�,�������-f�g*\3�vVe�l`6Z'������(��P�$r*�{u�ǈ�C��D�O���X�J���S�}�B �n��|E���y�����b�3hUJ��)�ƿU�_G 5�GǱ���BW�ю��vw�a��8S[\B.p�e3MMOwûE���]v���-z�p�A9�r��~�\��bE����/�(z��M%P>��5�d����vG��#	ɢ1)[;s�]�vp�\`��x}F�E�J�@sX6�Ssun��q��m-����G�tT&m*�0n~��S>�$�x�,Qkn�i���`78��ʻUô[.b�	o�'B>��ol��yѹ�f��̿���G�_�e!���~�n��;\@�8��;l����j�i�� ��2�s���~�i�51b����]X��T Je_�<0��#���AC�2.t�"�>�-�����a>��<t4��a.4�7׾*���yS��B@apL?'w$�=�U�j�,ɨ��6s�_����C�Ozsqz������#��@v�T�p��e4;�'!6�ȗ��'o����\�s�jP�Hp0��������CDp�_!��������M�
�G��p�S�4�l?�Ŧ�X���f�\�AE�����FF~E�nn��,_7�\�����\M�PF>Ӂ�W3Fl�yD�V�x�VP+^.�g׏�q��J��ϘSG="�;Zrl���B�'�7sܺ�䇹
 ���C#�R��I�l��[~rƛ��]&zj	����$~�+$��~g�#P>���܇����EH��!	 �����'�=j�ݎfa,�a�9s��o_bqΞ� �`�rSu��!&"�b[�*��2Lk�_�y�*�B�z�jG;d9�Y�p����T+
�e˓z�Tu1k:
E8 >�{�A3?4��Ӓ�����N!b�6��� ���U�r����b���������Ě�����en�
C�dO!�G�p��Z�X���A�G�-(9�:r��BۑPaϰ�=�y�+`I���sG�6<fv�5�_�c�IR�է��"~�x��(U|��#MY�<�ZC5��~���U顈�w�G�y�F����H3�����ϩ����l��|	�1]��u�5i&��>�P�����2���� 0QR��}���q]�~����h{?+�7r<�l�w��Kz�5>i��4B�<�K���N7�#E*�~�f��oL�Ba*~Z@��9�Yң4d3&w��L�����f��ܘ-A�,��6rc��w�D�?��F���q�.��J��A"P�˟��k��{zR�̗��Y������p�$�{���=��ZY�����U�zҷR})^{��J@��ޤ��(59:��}��L����t5��wM�|�*�z۪�*?7����_��K�z(N�Q����������L[8��\Fw���Y�~cN���^��t{�(e�"%g�ޓ�u�'^':���R!�}R�}\����GZ%�
����Ͳ"�ܡc>����F�Ǘu�8���{������3H�wt�I�iӮ3��wB���y�3��TS�ù����U����H���b�1�JǽS�㞷���jғ��	����H|����a�w�M���`Z�Z�A�����K�o:�k����h0�t5}�w�I�"�kr
~ǁ��/V-슡�%�ЮL�]���S=W�b�q�2�K�eB(�>�:� t�bY��f)�~'�F���������dJuA�S5����fq5%�5b�~0iA6��I��_�3e"���T�D2g��:܉��j�o���:jKFUfQ�BP�S�4w�� �$����Y��~���I���g򜜈�*ް��������A�E���a��t5�B�A���"q���(�G��g+--�5���}��b��H�5O���y�śd��J�7n1����3 �;��?g��ek������Ym�E�e%�@���F�L~n�WH�`����noO�3b>0���9����������M��_�è�L�4�c|���̂>�f�_3�,tܖ$j��^b��^B�g^��ȼ� ����aʭq�4XU:j���q�pl�+��s� fk��zC�C]����qt���%HEx�3������wt�l����ڧ�w���?o���ίtY�B>� ��η��^�-z��M��ԶӺ���� Ű��H}�]}�!<<?O�,�e1g�&�.~�5�fA���`�O�n�����]��²��h��Q�ݨl�<��L�b,�5je4��^�"����c�ZN5	���w`Zx���o�����nn�S��X���	�G���\ �*ƙ\F����Y��Fx�Ԕ;k�(e\���Ֆ���:!*�_�p�qu1�t�);i֐8i��ź.�*u�u/�>qJ��Q�W��B�W�y�q���̫��jV$x%0�h�3W�`RR�Շg�.�X(���L~�iY��c
���
B���g��k���.���0ۚ���)�y�_/���#Mu�.�ޯ͐ң$�ʣ\_�Ѩ�Yxq"6��|+opv�|L�5�?��:� lbo)�H�gM��G�X�e�sd+)�� M{_���~zvl����y��Y�g���Q~���}uսv��|�F�+�p}V!<�����HE詼���w*K��#,b��;�?���u�v��W��zDc-[��J���M��c|&�#���ir�^�L�������"��7,�7套r��;��%��ȯ�y�R�7�Ե�۾f����/%@�H�I�;���u'I�1����a�Y��ޒ�Q-c�p�쌤�l�p��]��A6G 75�X�3 �p�1���?��)62�"�rذ�:��{�y�U{@@3f�a���ԛ=9-MMHR{Κ��5C�au� ��Y�,\�o�:�������R�'4��Y������ΗG�@ԁr��R�(�1�����ڷɂ�p�!��4�n��f�G-Љ(Ȓ��J�]��M�LŢjl�5��Z�#�C$|كq���E�p�GF��dZ��M�C�͠��^�;�m.v�\�Js#DuЁW����P7��������i���'6\��6[s�N�*h�(�O71��P�M��،!���$T�m�M���	!�u�%m}�ٟeX�����{c��ƚ0@+�VH9Q�%^�g��������f���l5$~nϢ�B�<q�i�������뒾l�� D��4�2n���mx�B-���"PW.:՟�$�RP��6��q��;�.8�?����!b�VCس�&�/$�*�����z����e���B|�)��\1�w4k��mκv{/��eO\^4O��y�@�� %y*6�P��f�3*93�jަU.�����l����
-��_��22�G�-@�*�ıp2���Kܪ���C���� F���z�����\��ε�.Pp�㹜�#���<��F �o����6�U{L�����<C�G:�6�P��/��_�hfz�&���>�ս� ��:{6��KV��d���nj;l[�J���v`Y�Xy�GY�&��6G}j7�/x)r�_����X�/��8�a��L�}��~���@g�a~
��}� d������®u%���9!Μ��3}F���JqG1lXXM~Dɛ�6��.c�S�1Iß'<)�O�'���ʶ�^X��4z��ЛR.�97Nc�T2���Z��52y;�!K�^r���l@S	���'����*½!��������m�3M�E�"�����^0����~}/a��=�e�/Zfl��ޡ���n;�s�����Y���Z�nm�Ы<���<}9���j%۵�ku�J�*a�$<Zus{<��4��Ԇf.�i��;��= mᔂbg6 ξT���ȵ"�c��I�{﬏���<Y��[t"�X�qN˫���9�Y�V*ep[ wtZ<�~$�yiT��6�_�}sU�O`ې ��b��Tb����z�r��.�|��[έ4Mm��$r�i�f_���@���G�6����%Ό�减���	�g��gxrf�*	˵q���zU�VՑu0��2��R�F{^�o��<R^���VF@�>�;׼1�<���\��6?���Qu����μ�f�������	�Ηf��2j��u1�~�8h���^6Є����w-q>P l�(	d�v��^�.���@M�j~�ǋ�ğԭ6�o���[�ĎV~u����des��q�*��W��.@�=K�fm�:l�i�}Ǧ��z�:�&j�Q6|r��ʅW������p�y���H?�b�]��ֺ��S^<'�eG���4�����Gq	P8z� K+6	���I$	�Z=w&
��P�߇�Z:,2 �_(��^�e��y��QRo9��#��6�l[�^��R'$r�&?�\,"-���4hCP�?�V:�G(4�p�0:��� �MF(O���$����b$#!�F��!1����,�=~]�GЋӳ�Wp�g ���'�E%oS�R�2�7�`w��M��٫�-�G�L��³]�x�[��[��;���kv.9��"��{���'o+q����ڄ7���������N2�)#�I����(��Vʟ�Uڗ���ϒ�����t#�T� cA\|0���-է���re��j�9�]��!c��22�v���U�݀}��&Ҧ����H�=4ϒ'�rr�~��aS0��MN��̳4$��i5\=jr'�N��T[8�4��2y@�k�O*c�1���\�[Z�_/��L-��'�4~�,%4S]f�-B��ktm�������4����v�Q���C?ԫZ��a�H2����}�H3:-�G���9�O���W�h;���s`M��W��8��>?(��*���d3IRB=<֘�T�ԉ9J��9-��Ң������s���wA2��8�5v�� [��L0=6-�
`4Z�b�N�`�ծ���@d�����>�rR\�<΃�U$�A#�YB�?�!�0�c��ޱd�f]w����)�:ZoB��j7��J�/�/?�HL
�$��)aR�OI��=��/z�#aH�(Ef�-K#�/ʡ���d�ơT鄇ɪ��`YΙO��<+���ݛ�ʂ��2�R�C����!�]��,��u��.�~q�Un����t2Ͳ0��gzcf�g�t�Eb��>�P|.�X�v�%^/���x$N_�R�}�F���`���N���0}׮׏���x|�v� � n$����C�Ɋ�7���x(�.^��x����5�����]y2�Xw��`�:������gN�U�n���� �j�{u�_��ߓ���)g6e��z2ws j][�\`XqCJ̿b,<�����Z$���^a��1m똈����1�8it�ˆ2�%��GB><́G2�I��S�>l��*��y�`}�yޭd7o�����V��m�Ч���{�d=d�8C�����(�B�j�j�������8�
��N����Պa�<��K�ZK���z��VKiɋ��b�2Ky�o8`	�^`�����F+:c���Z��������5�S�v�>�+�M4]�%k%���V ]�R$��h�:Q)w��d�h��p=߆��P���Gh��p��kx�����D`��F[y���S"��8�^��-�r6��6�VѮP1G7��V�i\+Z�?_�X9�;g��4�) �U�7�1�Qo���g�_'X�]Ĕ��@�B��&K-���O�VYH�����d?P�Z� P����̪��>wi�oʁ�7U��k�@�ƪ�dJ%��q�u�1�Ǝ-��H���������]:՝@F���=��/y���Qz�3���G1�ơMP1Īs9�t9��k�T8����.59x���5�~Yqf�D����?�վ���N��;�����n'O�y��J�� �B,5,w,�����IνZ�o��lxy��C��D/:V���N=�c��J�x-4��.�����NW�jtv̳* 泰�^�Kob��^�e��ff���N�K� �F��M�5��|��ɖL������o���3x�r��ݴ4�^I�~��g�wV��s�e�`P��K>�Z)���n���3���������O��h��j�f���tFu�0��^n�5}7Q�߀���qO�/P1�j��;��j��:֑���jydߦy�h�+h|�h^�	:3J��k�|d��&�p��β ���w�"vv�-��{g��MY���\-���l�,��v� �?�o�eb]=Q%�*���5�ۅ>��q=���C�2L���m��vt�t]���(���I��=�~����mC26��x0��E���h�l�ϐ���]���7�Wt�DM@$�� >��%�_��Ұ{�ek�Ϗ��&ky�7�7��^�m:�3�2��|��*=]=�w�d�w5����#�°zp_�-�Ҩ��z�]4����s�*9�J5Ge}��y��W��h�~�'����AE.�� �*P�u�i�|c��ƾ���r"�]]h�� z�[A��e��Lrg㳯�X���c�䕚牫�> ���f;�k�0>�M���܁ 4��ϩ��,�-�P�
)�q9�5��W�Ξ�d�l����.j`1���1���ӂ�X�B�qȗf4�e/��j��3^X��=M�H��뉯�|�n>�����vJ}�+�/��Wl��br�vD=�i��l��~����"����lc6~\}�f��q���Iȯ�]�{qČ� ��I.���-�Cz57�+Q�%'՚��賔�6�"%�I2��~]���ׂ{��#=(�`ݮ�"/�`�	�����=?��m��An��:�*TS��x{�JPf��<�5�d��o� mCk�|� <���5AFP5ZehXo�K��Eu,��Ӥ�2�F�M���� ̱�|��R � Dj�����?��n�6�v���}.9GF�M�L����y"s�0Dx:�c����cvX� '&�	�|8}Pb���k��t�\�Z=A E�5���׏N�c8�Ф7֞3��cKbȏ������2(��:"�$�R/^��%��r��&�� ���º�(M2�إ��]K?��8�O���<a�D�ܲ�����3���Q7��~�	��.�%ڧ�̀�GbTd�*�����J�����a;���JY��D�]�H_'��1e�Ը]��r�<�P���f�\���*s�b>��'���(���4��(��}+���W*:�8P�9<5NuA��e�l����y�{�;�1a�w*ɈnX������� �h2"	��ˀN�^P��)*ȹ�W��w���1��	�U�����c	_y��fA�`[�1�7 �e�'w!4S���!�`�cp�b�4$�Y�zLJ�ނ�۷�@}j��d#�?���)3�	���/���\�ip��P�D$o Z2L�����i���S���NsX�[uX9�6(����ޕ�d���~d-��j[�{��
Ͷ.�G@w����
zg�
�:����V�3
IFG��\�Jn�ǰq4�i	R'��^H�H��R�͗X���%�r~{3��ܓG72��z���b#���ǃ�>C��z�@���>|�� X�-j7��ޥB�����K
Xj/�G�������K�g\X�*tlp/���/�+D>�k��t����z̈�]�P��Zv$�D�2�#o�g���Ae�<e\Y�m<ĕ<�h�wF{�C/�a�ݶ��T���)t���1�+��E�|nm����^�MK�ԑ��7��Ӷ�=��	Y��1���m:�+�?q�����e���RJS�C�)�N&���ys;������CZ��Y<� :��ZJ,�Q�贠^�Ғ]J�j�o ��"���~��# }?Є�ީ�eIr�RVk:�`��xI�������X�Y��S�Ѥix��\�M��S=�����V���vȄ��+��z��J�Қ16�FG��r�T�h�տ���� ��q��*�x|~�ˆ�n��P�6D�GN��1 �Ï=�0�4M2�~|mo��U$^X/%=�iOru�=ܶU�P�$���tW�!���"Ұ���fB���Ʊ�>M�r�ț�ֻ��^��`���A)bS%N�J��3&W�L�m
������<N�����P��"u��:�7�G"�ר�1�usv@���q'W5���8؏/�[���h���H`
���1��٠��8�"~5US_"� �m�(n�O���F�O�~�;�DD���	mam+!������	ܥ���4�ke�BN�%��w����ڄnp��߰-*���^i缤�hW3�jQ�W�y�Ok��O��i��k�_`��10P"���yN�9ԖS(�N�Eb��0�����&@e�)�P�]�ַ҃�.���s��_X��f��U������й�+�יִl�g���2T�Q����1�d��{|30�z-�����vҟ����|����,�sǐ�� �mxG�ăkow��Z"28F��U�����m��W0�B����G���V
GE`�W��.�x��h���vDDg$��\)s��0L$�%@�*g��8ˈ��xr�l]�sM��8�vn�D$�Sʘ�/ �.����)2�%\�� %�5w��R]���n)us�xJoI{�����gX�Q�G-����^�2��}/�����X�/6�=m�2�_��=�
�2%���=�D��PM��L
��usP�6�۔4ަ��c	4Wu6*0^s��� �G8�e�K"��E��Yap��"y~�^�7���ʇ�V�%?�Y\��t^�F{�.ή.~FM�M�X�L%�0$\��e �<�D���#�8m;�j�=t�Ω6���˭���.�*�s/9PHO�������G��ʦ�������nYn~��9��)w����K1r�����ġ�o�� 	�C�i�_���nA���K����4�zt$@�d�	����͛bu��?]:�g1أ7n#h���LO%��+�fvu~6����8߃����à*��J�'���lL�M({d��2Cǉ�wh�
�n�$z��}��yZ��aB��i���,�m�����-W	O�N�Ey�^���l��_��3!��.� ����~E��
��c:�+�Ը�H���'��:MɅ��z"1�w]�A7ӄ�!&���A���<&��Z�}4�m� �� ��Rqx�X�	ۄ�5�|�"�s��/UX�����/=]��`c%���y�Ã���o�L�'�ĨH���_�Q|"O>���xyQ����LIt�ҡlŷ��z��i��n���r�0A�D��o�v>�~��P�����Y �w�g,7��L���	o���&��/���_��՜�+,P��N��Z�6r�v\��ً�;a�2�Y�x��T�<���!���x���嘎az�Fh��XoR���w��nU.��L(���M�]�����-3��~W;R9ݖ�$}"�5A�А��BQ"7���v6�^�UP4�E~�#S ���^��b��� ����kc�\|j3%��N��4���fzT*�>����@�4�����V@�Ҙ�B���M��
����]�_���I #B�'����3v�Z�� � �2_=G����F�L ]�}O�hL�iW�E�)t<ù
���$�9��'�P|�ԉ�;�OB(Q��Ƌ�N�{�a9��>`f�2��1����A�^\Gd����&��N�Ge��L�H:��*K#1u\~V&���T<�&��a�T�Ț�����|���ِ�ʒ8$t|{C��m���2�J������K��xJk$l�Aֳ�7����	x�>�Ĕ]��%n ���1��K'���#�dS�6�.ȏS��ɇ�
q��Ȯ���'T��F|����M��D3ej�Z-�q��[dG�8W�ZHfŤrz�1�ʃE�IQNY�U��_FPx9��1���?@���c�_s�a]i�fYqx��*�����Յ��6�Bt�XTO��`�6Eπ�T�Q`b0�KA�z�O(D����}Pq�hY�B�.�Rkى��I��)+�iR�eSђ���q�L�ڜS��u�b��6k�t,#;'$P�J�^s�:D���&��^�ń��5����s�^�����,'��X-���N}�%��+�;����j�C%\#���[A餎 #{�t�,wD-3��$T���	c%fng�~RMQ���x�����|Hs��=�Cd>�[��Ada<�2!ݣ[r��f�К��(�Y����_B3��-bMKG�����dn�ݣ�=W��g�y�#!�+�1AUe>}�k��V�-#|Q�ܠ��o�@�hh�&,q77�H2����DZ�\VZ*�t��SO���I[L��~��'t��I� �5n������L�f�	��>g�H���D}�6R�H:���fG:�W�����vtB���+6��E��cM���X��)[�k+N��M/+H��k�)�(^�㈪R,�,�K���UE'��6J��1~��C�&��6����1>z�s-��� s?�y��AO�%���m{�D�ʟ��*%7�Xg*^�O������cء���=F�?w��8/�.pG7�2˨�
t�$�2�̽����wF�۾�D �,�֚p�C!7�`��;?�ʧ9�9\��="΄�\q���{�_�����z��ͤo���Q��,o3��~��e��'L'��"��J)�;�qH��=�hr��d���
��u*" ����[o�� ��a�3~ѽ&b_BS罃.�ج塌��C��~���RL�m3�pEz̛���x���b�����Th��k�t,ox��8�~��[��|��?��*��bTS~�T<���'�Ə`i�l
QS��w�p��8S"�FS��}��V�h�G{���J�#�?�����1*�i�;��$�?��)�E�w�%���qXP*�ރ� �<���E�a>a=_"�aÐbd<���1�g@�0Y�c�]�LE���V�������E�]��e7��	�ϋ��W�����M�+���W�8�e���߄�V��I� �t5�F�-1�¸�D⮢/��8$�޳�o_
8B�>��-vW�f�,&���0�?��y�pB������b�z��{9�M6� �e+l��}q�lN'��5Z����ezzʅ�x�^Ɂߺ0�X:�A-D��{܂�^Ak�J��ȏNL�,r+"���k�CM���/������'|�\��&�G
����R,<̄|�͵VM���3��DʛU��Z|������6{o��e�-�����%!�[�an��;�拀��_9�2S�]]��j�H��Z%>���~�qj����-��v�r�w�#�´�jkTIl�WT2�|2�.�1��	"�mb���ܧ�Ξ�x�P��w�[\�ӛmdpʉD�u{Կ
�5K�h���ZʕϘA`�{Sݦ>�x����2D��;������;�nۑ�G�RC��@ډ�%���o�	`{/�%�m��V���Ѫ4Q_�ekg�j2c�I�8ƿo�Z���\��X��*,@�A1�o}[9,ۧ�&��+h9��NR�����T����^d}��)�V໔Ȭh���j���;v�͵bd'�y�WF��N�Dy���&j�ܗ��U�n�Q���v���ی��oE������j�[^ÃS|+[a���k�HMk1�y^�4��d�������.���71��������,�[���Ac��~�\�f���5��!p�j�a��v�GP��m�
�Lُ���j���N�b����g� �x0���b�Uڽ�A����p�e�'����<��ȋ>⑈4j���Ŝ�O@�Y p����!�2��zB��p���b���%�/ML�J��ɨ����9�x��H��}��K�$���ޖJ�!+�_�ق�.T�� �"O)f)Ŧ�9��|���6	v�I�ҕ��>��Z0���p�?��ƛh��D�X�"�t��29l�4_�|[?~�5ܦ�����&�-��ުqVn��0mF	��ƪ7�Ͳ�a�����)vl2ض�'��,��|�B���J�a�Lz���p��I冚y(�X(9��ޯ�Bʅ�CFD�88b^tf�x�>�N������g��L����2�;���""����pA�ꖆ��P=S� λ��`[1�˭O�5�\6��D��@�����SrCAO~p�s����
B��p��M�ū��e�p [P����%g�1����{vd�!b,�����	P�M&��c'��L�jO^pN��c�A��ʨ��|�Y�oC`�����3�]//�6�����arr9[+�����m�*ꮏG��[W�-�܍e���������ˋP���`�qBT56��Θ�O7l���D��vC����D2\�L�riU��)M#�	x�f�r�蚷P�~�7���#q4����:���̓+]щ@��� :�����¢�.���Q�/�/����H.�b/��.j��L�"3�5Ld� e��vv�)sAV�g��@�U]K邟K�'�~�r�/݋��^&��#Dܾ��8 ��9|e�3����n�-���Q�'�j#��k_������1�����߸ZN�����7�k�k~�sc�e�h��@=�X�
��jj�4�Uo��>���wf�E2��T1Ԇ�Z#܃P	�!&�T�H���B��)Y~��~������I"Cok>f�ӔꚀ�Ķ���jJq���y 
�?m$����� ��A:�����jvco�h�GR)}\[]:�Vc��Ԕ��۔�닆PF�8��-ڹ��x+U?	����T�pAw��j�n8>uƒ�S�;�6���+B"�Tփ�g�:a���W�+������Bgp��-|�wy��2QSLA���p�=�wS���Q��{�SAih����z�����X�Z����������e���-rS}v��6�/�Z	�8P+�~/��.Rz��ؕ1�b.2D�q�����U��ppw���-O�c�N�aw��&Q7�ŷ�fXH�aWrq�r�|u��c�:T����f�����͏�_!M/�Ί�O���s�����C�D�(2i��H��!}�$�*Wf���4��$T���A�ޭ(�\�;�g�A�)	p��5��S�x̜7'n���Q_��O��U��^f��*���P�\�7�x�S��lA��	�s9��pY�y�uj�:�_�'>¬m��M{�c=��y~g���z�Ӣ'
�^��8]W��J�������w;��/�" Mg���Ti穬ķ���F�ytUTg��R�[���n,7��Mj��I��^�ue��q��q�O6��y$�{�����k�v�Gg/6�R=��l�F1��O�.�q��+ �JVAQ1̓��̲��Uҽ��慯����U����ܿh�Q�R�Q���2S��Aj�O�s��������|�1��au�罥�i{��h�w,$�ֆ�Ć��"�z���RT%X�tA���~#�|�~�h�>iD'��Ng����/�M�Q��V�1�����Zd�?ԣP����
��%|9�`I��Q�F}{W%	���ׇ��g>{y.�}��d^E�va�m�8Q��� A`S�b����M;i���^�]���E3�F��4cKy��&Z��&����)�N]� ���U�O�	ħ TE1��RM͓��}v<5����v������lC�Ja�k!�?�-D���ƍ�c�Q?R�~�N������be� >u6n�0���붒r��)�����|���*[Y�u�&�ѰKAy�B��;�5�WW�Ӭd��y�|�<�+��$�	���;�b��J��jXg-���"ْk�N��5w�� ��FִC0������
t	�H@���O;�{�<'����#�����ԇ7 I1�}�4��*G6��Det����MC�𳝗���M'��J��tQ��XƻY8���A�%�1���}�
/(�+g*�6Z�%��J���(�q���z�v}���8O��)�m�}h��/�XcVS��e�<�$�*���ȗ�Ym��K)_�1Ԧsrτ5��<~d�Z�6�� B�C)�Ï@��,m�&Ms��5J��+�9���{�II�la��Ȇ�2�;_��)�쳐��SY��%X#(�ȵO�Rg��6-�����aA&���)!�>�e�'_��s'}���2�Hv���ժ~l�gtO�җ�`]{�
���ʙ6�s�^?�{��c�.D�Vl��*�o?��O�_��F��c��G��Io����|���+�R����@��pc9 �?�3Ե��"<�j{Lmx�+U�rHL�L��M�C��2�Yc��^F�+G��3?��}�*X@�`�6����DS�BNϴ'��w

q�8_�z$��c�y-��;?�B�%{ ��D�'�Ð��}�+��"�����9�B�?:�x@B/�C����sݗ��[=����o)��3��Lޝ���Yy��kC��P��]�v������
��IiM~I�����@\�,���Y�ʮ�Pg�T��t��(sS.�e��G`O�6D��"�Zg;�4"��Fs.�\���~N��������K�h�6 ,dh6�X �r�,�*�3��f��n��]��"��2
��M��������m�����9�-�.������?#Ĝ�GN5��u������qWe�Lݽ��o�>A�h"�з[��/��릵s��uD� �N�\+��*A1XR�d���7V�@Vf'��G����@ph`�q!BX�����'�Su\���dw�낌T%��=�i��/e�!�Z彫�!<z�Cn)��!�\4��G�`�=�Up�l�����pF�i32z�[�&��z���d��/1)���K�k�B��?e��aS��3S�T(�E�݀,!�!G'�材l��+]Gh��Pޮu���a�a�h�C�n�V^^��;yc��#�\9�V�Υ�d�c���Ec�;���e�Z�p΂'�F�����1;��PB�#u����*fq��up��=�mwL�%���f~���9�2X٦^B�?��4�����r醞���>�j�r�$�� ������}���������;e?%�A�dp��F�ד���Ie��0����\�G=v��I��6�kڊs3�2��p|�`(._������@�x_l�ә���qN�ΡYF>�dX��?Tg�2���
��2c��#?C1��F;�>
w#6U��#㍣M �B|]t�)��vg��#@1�.!@S��m�b���u�ub�\�T��?7���Duʖ�A�o0�wL���Vk���B�!��(�%������g/3Ӽ����3%|R���ǘ��(��a��L��;�C@�3�q�'<t��M���kڹYP�`��~}\����]��z�����W�a��A��ɱ�o���m�v!�ܤqB� )�i�Dr�7"����6s��:/jfYr�ھ[f�)g����[M2��pY/s��,J6Iz�Q5N�=��X�A�6A�򴂋��%���Jqa :C���Q��(ص�����`����o��S��|r��.����+�pN"E2��}W<dzuyS��_��?K��ώ��ɔ����1!ޙ��QXM#�U��B-8���o9�А@s�a�3O�3H��g�P��O�[S)e�%H��lN�pG!+u�.��c��ւ�,?���3v7���PO�c�?�'����Ƀ~
��G��B�4�8ˀ�5-�ր��@��Jk��*Ԗ�r�W��΅YQ��g2}�'Լ�����Lu
o�����T�$�;	2����='ʛe��^��+V�Q&�Fj"��䀐^���~܈@0�����8��Q�7�o��[�Rf�54�1�>��7)U��	�Q��wb�̬�E/g�f7�L�$gB��Χ�g(^a"��b>��D@[2�e#2&֓X
Q3�Xu�b����t�A��	��k�,�,2�Q'Ρ����_��һA�P�\�~"�?K�NI�1��.^�%�B���[�����E8�L,�Q���w�ʙ
cv�]���� m�wʑ�[��G�F3�z���A\�C��6�b4AT��Vz�8�9C��*�� ��+�a{ڔ�2ج����c���P�Z{`�݃�r$��'�v�<�?d%��;���o/��p]����HA$���ٕӠͻF���;�i�V)� ��_"�6_��O&
P����PzѤS΁�IL��/�gz���ǻ��������N&�iɁ}���˲-������ jcȽ�';�ܯ8�-�-��ܘ��A������Z69��/�n�޹��w��A��'r�c�%G������6�y9l�b�-,�K� ��ݲ�USSH�:q�R��`��Pe���C��w����B���O�]%�0hx}M�/qv�x	K��Π���,�MĪ�R�Au�|A�!�G��P@r�x����H�ȇͤI�#�neA,��#Q��py�O�F=�^}hؘ����#������_��<=q�%�v���������ed ߅�"�y7��WEp��t�Q����ΰy���Hc��P&! ׹�jv��.s sŌ+[�oĆ֪�Мq��,���Lq��d��RRO�nI5�-f�|g�&X���m�k��:��/�/Z��."[k�m� �FN�j����M����c�9l��/!{YL7׈��8�3�L��9q Vܒ1�IN���t)S��'��K2��}��˳*W8I��/�ssZG;T����6�@(�hM( �G�5�(��]B0W��5�*��Y
	8��|��d���0��A7���������$-ϵ2:vHvEa3y&I�����:P�1.me����O��4l��	Pi�ў�@�4�Kq�~�K?�
5VB�\i����CQa|�\�^M[��T~��i/)A�B����f���s���n��7%%n�ɸ�,��׀xX��+Pd��>-�uZ|mE�*��������a�V��k�_��l �0k��Z���Fu'P.�-'D�Ku���aU�]�Q	t���M�@]���{$��;
�U�D�m�t���j����PJT��u�/G�	I�q���tnn��)$.N7��BZe@ŷ !ާp��SK��]�9�R�[)���M ������҅`�W�ˎ�SS�2��C�gð����ebc�rc-�*^
�J��ꈜjyP�6W���U����!Bٛ)�D�B� ;U7x�Z&�ek���h.��p�X�x���GE�ps�J}ᶼ���Z٪v�ԽE�Q
e�I���%}�V^)W�2A��]���:�D��������X���Cb�6�ά�Ϣ�
�\Q}lXd�H�r����b���-x�v�gB�st�ߐ~�DϗT���l~Z<�7	��aQ|����5���>\��q-k���j}�\����A���H�f�d���w��;Ԑ�^���-]��Z�'
K��7��	�I.��r�-o�`$�m�#��Q��/��텚�7�k�2>��|/�e+Dy_�?V])`�m�aq�(P�o�CII<� ��E��m��ݶ�H��������t�]9�n������<m�% *חR�v��<��̏�v�.�C�H����Dv+u�Wr��|�Ţ���F���� ��9���ǟ��2n�DC�̶t�r���Z�q]���9r' � �^��^.�M��ϵS�+L�[RI�����S�:�6�Yz�9���o���ѡ��;�*I]}H�AUzC��7J��#�E�֐��3)��x��'
�O
���Jɰ�ntJO����1�H�:�7 8ߦF�m��ڿE^�����XQ#1�׀~�L~��� �]k$V��$��i� �V\��q}�����$t��2�G����m���_	��$��\M����F�8Ü�"v�K<8#&9�vKǅ�}��⺃�vj;�:��P�f�����~Bޝ�-��
�PӐй�O*�u�7�@�d�
�QGJ��߉�ʐ(�������p��P����ϩ��W$��M+bz��j.2Ug�%ب\� I�rIT�ĬjRۭ�mn��	u8�t���0��$�x��b�@7�un�Q!��y��Ӷ�]�bܘE]9LN&T﫶4�Z��qʋ�w���6؇�%j�vY��o���5�4�Y�^,LSU%�!j���>���R�!j�0���i֦?�_N�+��m���@JA���9�Y�{X���Ws����9�)c�u��'�|Pu/�f��I8�xiF[���=&�X�$�l&�`��
ww������[Mwܒ7��G����-?��1�R�)&;L���:�'Wȕ�	�sŻ3}�Dg��R���~�e��f�.h�6ѝh����}T}��=1Hs$����5�g��J���4n��]�w����)x�uࢠj�u��O��j�w����?����\X�QF��4_��H�ٷ�on)bp.ǭ�armws���Q"����"Y}�itE�i�QY@:��J�7,N���_.mb��}� +��'j\9G��Y��i��8Z�gF_E0�Ú����i�/'�e�l�]}*��&3Mƴ�io��{L��������v��[�7��Z@�t+0�Zr��~�f"�m�Ni5�k:�}�V<��MC1MWh2����<(X�
���%��h�V�>"w!?A.9���ԩ��(��~ߥ�ٺ�,����Tl��;�k\H�)ٗ�l����zcB[A��ֆ���̡�*B*��H�
�sv�N'�*8����3��q���C$8��D��q�|�������<ӌ P��s/��^�(Z?;���v����ľ���ݵ��t���ۓMy�CU��2�:a��g�C�*~Fھ�vPz5*�,����ޚ���j�����sfH�m���j��ژl �0�3��;�+�Ő����9����?����!r{�+����+G�τf}A^��К��}�QKp�S�����D�X�
���<b�7�c�?�}8] �|V��-�h�>�Q��YI�ٕ�5a�ack�Q#�gnFf�_���2�]L&��j��m���#��Q�P˽��{�~&���̕~�y�,��3V_�y�<�X���T��6���6O����OKM��ZX��8zq���9&�r�$E˿�"�`��Z	���Ŝ�Vx��X+Py��30���]��z[�L�^�9��M7����$��t�Q.�O\�M��յ��pX)�2_�&b�� �4I*	ԓ<�  �<�dv�"��H��	��7 \O����7�h��0��ދ!�K��[!��.K�#����K	gR��R^ �F�t��(#<�5�"b�xމ���)u�vT����3!����#h�@���K5�|���@����!s��}�?�^��mԃWc��Һ���8*d�Gy&�MD4 �"��}v\�啍f&9������X=e�BN��� �}��ST���K�� �h����OO�՗�~��c�~m*�GTr���$���f�!ez�_4_M�A�� ����j��
<����Qt�z!��N��%�`�ߧ�����m�^��������Q���P'��U7�F_�����4=��N�>s�f����Q_��j�][�L���n���g�b�X���t���EB�btyh	��{΅��x������w#)�ٞ�W�`��-�6�{"��\L!���˗�d��{�,��H���N�B�	O�3a�Y:�a�y5�ф������+���}\�%�b/���W�C�3J�E\EV����ƫ�w+ֱ�7�O�����[v	�@Ҷ�/M�Q)�̈���_�{'�$����l�?�����:�b��#ֱ#`��.nSx�`����כ�Z!��̔���sN��$�N�.8(����wx0�KP�"�J���
t4a$]�$���x��g��u�Fw�v~Z����E�u��J�B� jF ��e��Ip��H:~լG���\R%���Z��+���<p��ӣ����[�vP�c@�g=L,�-_DO�9�e>R���n��Ɓ������r?ݝj�Ob�bÓ V�ݞ�$F��6���K�'�ɳ��`ŋ�Ν��ͫ�s�/'�ZG���%!~���Q�Z���3Ŵc.�/�����)U��Q��%)���1�aOiNJN��?ZY��͙����� �y�U�'� ��M�Yκ y`�l�K�`ݘ:�����ڦdA�{I^�	~���aod&��;RD��>/��_X��k��[UA���8�Ey3����۪i����z-�?S����MH�;=�0������+y��^�f��^�!V��o��� \�x�__Fi�LF
S���nK��$��ECM�/�^Ey���\��e�V��c68�$�k5k�k�Z��;��Z�0 u+r�<	�kڠ��-�=[I�{:��~��w��j5������6���hd��"�Pp��}jA��x)��t+D�`V*5h�b���s�a�jc�u5�,
��,Ɋi:�H����>�?���KRX��CH�:��"��o���b�:����P��5�!�I�����M�gaKͻ#l��TM����&ږ����ݐ.�A�n4�#""���;��$�?����]��-J<��D���F�L�L�쭿���i��-�z�/"��x���	T�����}zܪ	sM�7b���c2ʘfz��X��Y|�O&��	��_��K��hu�!�`�!ҟ�s��qq?]�/����P�v&����jj��N05D�db�>Dk��z�E���]�����#��㚞�-���و�f�,�3q�b��;\Y����ddr~���x�b.~n$��a�ܫY�{3�à#�jkqg�1�����
+?�>�?خUU3�?'���Ru�a�c�8o. ��]M���s+�H	R����<�)����c"��I���x?�*�;��鳹a3����Y��La�ua �zn-���XI�Jڴa���fG�q�����_��1`���`p:��!����3�����(�&L��X��,ξo-��pe��p���w)̏xh	k �J�3��r�U�zu����*�3��?�-WG�?�թ���Ⱎ{�J���џ'j�!tUz.�G�riua&�r����� �=���얁� �����U�B9�ޙ٥�-��Jr�D�
�g*!5�|��^�ozh��>��T�<��l��?L:j�5�X�Ɲ��}��w_|�F��E���5H�
"`��Z�v�SXi�36�W����q�=ޅ
y�H��f�⠵ ��y��`	�\O��2$j(���N�������ַ��5�Zx��rE�����O�%���@r+vi��vg��k�:*5���M\��%s�3	7��8
^Se���r2�Ei^ts����x����1<����-���1�T\���2���A,�dP��[Ő@��n�!)���-%�.a���W S�ê�Z�<;���+�uUz�Q��hF���Ċ��L]uc3т�n�o��-��om�f���y��.�F<�d~��)q��co��AI�0�q��k��7}r�G��ە���oSi͠
�8hz�5��\���?��2�僩�&1��(]�A8�^�,�	hE��&����w�疊�f@��WҰ�h;�c|�M��0��s�/�1ji,�����Q��+��@U%�!t��x�q�@�!p�b)������GX������7o*]�;c�zi4�^f|pK���pEK��?���B(��tQn��5sZ���Av�{|QDqˀt�֙�o�1���Z��(!��8oD�a zo�%U��� U�]��E�XE �F���k�u �����h�?yN	�t�:�ݤ\�]k�Z���޷���83�U�Ge�$k�Z\�x�4[�`]H��q�3���Џ���"�D�9�.�!׫��-�\:�	������.��ž��~�v���i�S?
���K�lP�i��%��0A7|3x�52�@2(J	M�g�7��l�Hk�{|��*�W��U�� �xC
k��}��[J�hN;y]�j[�{v�4�Ш�{G���C��3�I��6�~�XU-��&�C�
%�!�����&M�\�{��Wa }�|R7�2��k��79�mY1A�" H�R�@�3轆M[�$Q������'[�z��[k�Y�L�ī��z)G�1��9�T��
�rܩ�љ��t+��l0���*�_��F˒�
lH��r��~����j=��Tf$��M�3�������D�S�#�$k��`TbЬ@+q���!�G��k����p�v,n����:5�4��YR�ޔq��+�\v��Y%I���?"��;M�:Pm�+G+ׄK|k@�%���/
Gf����4ڔ�q��%�C��������sr�������ָ�ڝk!vC\g顎�(WEX*td����]�>� F�s&��l�_�V�n
4��n)��� Ϊ�+�D�Yj���V�KT?���+�����H%X����I)��as6)�Y����E�K}4;��3�i�V߇�(0Z9>�)�� �Z"
hh�4+���$#A�f@�=!RH�x�/�:Mj�
�#8i�q(�o��g����68i�(�ub���&��M��c:6��8eb���u�ߠ�T<�k�>o���;��?�b�g���%8�G�`/�T@2u+��&t�pZ�)�=gb�����j�+��9�ݡ����t�Z-��h��a��^K��a1dAX��q�M$5+)�*�aZ�x�>�(�H�O��U�,;�n�LY�:ѧ�;�nA�VA�N�M��S��ˮ�42T�� S�C6BrJ����������;�>۵����Z�~\cE6�w
t��~>��l@s�m��G �|o��@ ,��ξM�)o�j�Z�J��DK�cƃ��� @�(�D���T�IZ.�	�?�Ǻc��	h��?�ˉȵ�Ɏ��}LO����Ȥ�ny�ڊj����,����)�&���ZV����D�46ޟ�i+�A)�
����ͳ+��C�#�>a�G��r��p��$�'�:c�l��w���T�_�O���60N�a��/B�'\{LOM��mK'��^/.����G�e�OX*D�� s	#J�Tv}9�<��������x���2L�޻Ad� �C� ��rpA�sw���C;���4�3�8t��o2D���WY��q�#�U�RӾ9��Ӕ8��l���?�:ǔ�Ȑ����x�`?���w�3FV�F�9�	��R�=jN�/ʢY�:1:9]r����{��g:�l7�?�������1U�@T��WM�M��Ju���7y�љIc\'�2�����<҇�B"�r�ג�F�zF�ˍ�־^R�-z�d���g�p�>�A�+�xc�@@�i����ģw��<9l����Y�$�; &����?�� a����>���7��<h���Zo���]�f�I�'l#�D �>���§����e�l��Q5�J�I��=˰yV�2�~��{!�t��	��ꆩ�~MG�c�PKl�o1
�KY�e�4��@(�)�N~�L�QYX���-j$�����#����A�*j�RG��tm�"��E� �Y}�	���K�����*��[���-Y�[�b�KB.�������x����/�0դ�*������]��&��M��Ne�}�W��!],.|�벅�����/T�jM�v*х	L_���z�Pd_x)��?AL��v�5F�|�����{&�Y�V�� }~:�P{��$�t��K�rE9m�l����Y'jo؁t4<�'	|\�0�+�J���Њ�AK��Zϲ��m�?�ZTu$ݶr3�2��!�%�S�?3�P�.$iBa]L�.Ļ3�Z�Ҕ�����Y��[+���r���]�̯�^@�&�2�vW�,� �yg腄��1��Ѫ|�Z(�#R�3��������������IuN�TD��w4���6��r�1+��
����ۼ]g�M5\��q��W6[�.A#@g���pt�ag�B��1��I�ŧ?
�w������U��;��`Q2�lJ����:[�zXh3�^&-��4�(���di-��ll�3�tC����D-���j��h/
�A���xAF�����\�N�y�,��3������U���fqϊ��k�h@;x�J�yk�-���_Py�m�� ����� �i{Y<�c��F�f8�����6y˸N�L�N���lj3�i����[Е1�I���d����+�-��k�L��Z�ْ��������K�}y�`�)n����F�isR���3�
�ę%� k�44ҕn���h^8|����ן��g���҈X�鉌�M?YE����0O�<��eau<�n�}ŏ���
�O��i8M�t=�������L�D�K�$Dh�����Z��r��R��ag�gl0� �q���Z8߇C�LT�4�[.�Li�4��:��K,?�P	�+���9��WmRҸ7-����z���t�o�u���tp=�e������qԡ�-#)����F9i�ҁ�6~XWYT;U �N��d�ڑ�$z�|��r�*��+�lKȺ�:~�%j�hH&���Ҩ�_1I�jۚ��@뵽��&�����}(X��t���)p��>�9�ǂ������mI��t�?�'���n�4�'��5�M�� �$Q�k:�|�FDM�Gk�]���%�3�1 a�v��D⏭L�_�9�{��G�XZ����������#T�TE\�A� �'Q0��TV��_�un5��CP:���"�B��.� ���ZrJ,mc�e||s��n���e�+�f_ٲ���A�c�j��)��!����OG]���0A񰐣�߶��A��+�ˣ₢�𖼈P#��lV�Ne23�;b=s���']Z_ba3O�s��NV�Y�'S�8f��������~ln��,J��ZN���ž�����ls(y��2d�K�h�~���h�H�/��	>+ ��Fέw�{���,�m6Ɂ���<�7��8�͐��3��s���#�0j��#z�EL��X���h)xJcU��� ńW���ߙ_����D��J� ��VVH�XO-��S�ݡou��U��6�Z�	B��|�q���-�TѨ���5iN�ꈉ�H�Hf���\W��40Y0Ūv���իins�|T�S7�Ib�g2&ûhe�nM�,�7��/\���S�Wj��L���G�Z����\�4�yr���҆
;��+��ӫ���]OBi��r���z_� pˤ��`����&���5�\l���v�-��^2��P�ߥ+��񦪲P��ڒV�aU��)rY-V0��8�r���4ewb�67	x�	�-*�jl*�M�=�+�B1n�Mz��ZMZ���u^e�����`�&M
�Dὴ���g(����y��z�?3n3kX?���+�B��̈́�X�e���;�!)�-֩�������	�ձ�f�9�M�;L���=������e��P|e᳡�J(�߈VL�S(�/�3����Uv[!��gat����J��.�1�z4��*s�{���d�<�����S~+a�Z��5�A�8���WLM&��?:��XU���٭RR���;C�v�����B�/9�v�E���$�������f;j%���L �љ�SAà�=w�
���[ܑ��/6 aE�D��S��^��H,���A/�5}��/^ݧ�y���0\�J0���"a1����`�+�iex�"\W E7T��� ���8�t�jz���|`���)���kϡ���:��^0��<��Tcx	��d�ZPr\�e�� �!4��M���T�ￒ]�~�h��6V�m�������i�'.�D��F�0�0�NږS�B� X�ݜ%�w����D8rP��	!�s���y�U�2��B�����s����4�a�*����{v�� lh4���?{��d�6x�r���X���)K!��n7K#�&HV�!�t�TE5���c8�Z�RQ�ئ�Uզ��
.S	��_� ����0����E�e>
Z[Φ]�+�@�D���5ְ_�Tn�!v�%Z��P��3	F������/�܌<3N2�q`���9Η>�«6샇����"����I]�d^���l��{e�Z��tx1�n�!��<�q�qʫn�@���1^�����r�1�k�K���ן�i��b?,R��b�`k]���f����������H����$��k��כ�u2�:3���%(_�6cc�0EGU�M��|���3}S�X��$D�4μ3�*G�������LUc⛒��i�'j���־#d�ڟV�ZCXGF�J��éi )%Ќ�~ا�(��ӬV�x)2i���B�/49ɷ
ۈ�}�32ĥ6FµZ#��g0r��р�ل�C�s,I!>��'@v�V�E��ƃ�p�ų��o��I��iY��mf�zz�� dc���:�Dv�yC�pQ`��3I���?E2�wi1�ϡ�v��?~�#�#�����V'�{6NӒ�W�#�Z���׼��)��ks�a��aMX+�Z�i�q�Teo&#��m��Az��3�=�Q�˗c>e�9��H�A銺5< ��8����b}��ǚ*�95��+;_��o�����){�̍��_c����LO��k� HK�Bt��O�J!kq ��3�йOw� (o�};���}�p��7˛ɅG�<sz}j�{�sa�����U�P�ťJ�9:UQ��$^��U��-N� ��Q[�`i��X�4��`��Rb�AF*m�vj�w��\�-2O9��/�<�_��I���V����L3Pڸ*��ڨ��o�Wj��GlUv쉅|ѭ�y~w"�%<�[�5�Ym���<C��RI��i�� `RC��W���\o���Tw	s�0�(=��&��?�{��-�2a-5s����u�ZQ��R����g�k6�p�-��n��������Z�Y,IY�vY}��K)E�_� ��f�J��7�~5��0�Y�%Ǉ���N�p#�;�\�~G�{ͥ�=���k��L
�b?K
5}��P���i7/F:�R�e5�LG{JL���m�9x_�-�ЭJieW�g��rÞ%���_���;	���7��Jشo��v�SI�:D��j~}�d�ou�,pXU���
��V�^��>��}2�>ulω샨�)T��EO�?���o+f�c���`���?���/�x����`�;�v�3���c��Ԋ�b�_:�U���M�f�u) ՋȀ�����N��ͦш�c�@����]w@����]t�~��,��½���|��1w���	|�چ�hcЌ����7g|o��~�H*����9�zA*~S0|[f�Y�O�Q�MU$8���j7R|L㇄�i��7��a՜�
��������H@f-=|���ȇ���`!O<��A�sϽQx�7R��PL̥tӏS	"�	��j�5m�����gk��cj����b��$�b�&�%ذB+u�� o4�Y�dzeTH�HtL�7S[w��p�8���}�?`V�j�����F�_�58��&��t�ύ�Ǥ0)a�\�F�ly���1������c?�c�⺥C:�D<y�J&��e�M�"��~�l��qɤ���6�ے�|	��-�Q��M�����#x�$��E5/���n0����6N�S#q1q.��Y��m褓��#p��^�W�=�(�ꠄ1�ť��4<9c�#�ٚQ�#`j:��Vd��8��nD�����Ư����[���QӁ^�S���:b.���З���Y���3�$������y6�N�=�}f��LH/,5>ᵔ)'a���"�0�m��M���4ʒ��rrP"�|�A5�9�n�� Lt}&%a����Ӄ^�W^����������ǟH^�P�[�]��~�����!h|�.�\���c%��z욺rZJK	��Y(r�1>kN1m�'�d�2܅F����  /���9/I-�q��6�]O!��;�4u%�oǗ��nIvjx~{�[�FROy v��"�")�T�w������I�a�FA-ݥ�e�c����8��6���Uh~���_F���0s}�8�\3��YTL��=�����nɰ���1v�b��@j�B�T���3WD=�tT�w俬���������N�AJ�0��JqθP���]S�ЬqOz^7XDp��y��a���婩�~�J]!�ߒ�D��S�;�MM4�98q�Դ���]��"j�!�j��>�rQ��h{Q̗4N��
zc{E
�z��I>VǤ��؉�0������2������e~���F���#��ҕ�@���Ae�̱�˦�
��W���@�eq`V��׮����E�?Ֆ�~��9��ܽ����G�p�QQ$������I�}?f��'��D}Aԙ��Ї�i��,�E����G����6��/�O7}����-��!�1&�t.�*`�MJ)wF�����h���SX��`[=�F��`�����W	���]v�O���_o(�<WsM�wqLU�P�P�������yl\6����&��D�ʬ���K~�.;�w�{�m��r>Ϡ�h�Y�?������1��f	��'w"͛�R���帰�=��i���Č�8~ĳ������d�]k��~r`A�ߺ�-�2��R`-.��s:�����+c�0��6�؄gsx�����2H��x;,~�ǐX+D�|]m�w��I� �r�h�IPX����^�X���Y�W��Q���W˱�[}�j�6�(=��՛
-�$	f,���qV�f����O�e�|W��O����y�K�<�w�|��}eA��8Y�ص��w���;!�+*)���:��k��ޣA�{e̬+�CΥ��;�G��g���q='�����p��L��X��ζ�[�oجuȒ�h�sG9.��^��C��l �3��DD���W�\�vqmq�د*=�z�~�v
ݪ.)�Y��*��b�-��LW�iه�cG����I��ü/rΐ�P3��i��F	���t�w6�o�0	1��J�9}��0�����+
�} O�5EUC��s�\��=����4lL����q8���7P�9&�\�ڴ��У�����Z����}0��<>��9e{S@ܼGl�'`�D�r�N3�ŤCu��F�i��2R�^�����0Er�5�Ǧ�ds����x��a����U���n���+��E(.�?)���*�),N(4P����]R0[z�=
�*��Hy�o�<�W�4��u��L+�	��S>����H"[)�.�{���.�ui�5�Z���:�mG	l-aZoѵ�����s��"����G$��迲M#�3�ý	��Z<=7�����+���ϑ��Xr�"���#��̋̿R��4}0FW���3���=�ҪI��b����Be��n �|��(��b�b����4�8[�R�� �9��~[q��~F�1�7{�v�B"�5H��L���=�ӀU����?�3�)�ն�\6Qx92�Ua/k,m7��ՉR��"���X�����WXY`Rn	�⟊:�.�����'G�X>;���t�y/�C�;�K�!ځ	�޻r�t��y9ӐK�g�V� ;�m�O!�{*���DA�T���[�e�A��:+g	֥7�o
�TćQ��t��J�Pj
�vݩ�6�t:�p�ԟ��r�Є�h�o ΍ƉW�V�9n*�@����-��.�7�j(.o��*�A��b��-�Y��{�	�B��ia����WC�6*�a�e�IK���ު�W�G�y����~���t��*n��lbN����|�����i*��ǌ��v�tو�s�-`���C���R�r�����#wX�s�����oB�f�)��c��Rf]э�ĳ)�`��7G�k����s�UX�@�jv�P̗_�=a�	 ٰQ�3#-��4�"��eYy�P�qa55�Ԯ6��.�ʕC};�$�H}���!P���a����h�.���+�>GZ�
Ow�3�܎ʔ�3�6�Q$����.�V7�{�%���P�1��Q��!�Ź��.�A1��eW�}�
�bԎ�w3��K�#!��m�b��܄�L�_�n��:�7��B|��A� �9u�4]�>7�~>k6�o��*}շ-j���}٨�W���3'���?N:�uR�~F�gV�e�T��QZ�~��]:�a�L� �սK� �E���p"��4zK����Z�q�eQa�I�sߟ�H���$ҥ�h��"zm�+ ��|��"�^�i<�R��&U��Uә��������xf ��pHr�O�ƹ�e���%��[��u�BA��y"� �@A�<2�CE�䞻��S��R6p��3�� �6��T'�:��7�{+2L��e��
�Er��3l~�|���<\9��!N>ɾ�s��؋�~�c�8q�8��%%����[�o�����V�np#��E($�9Q�A5��,����b�����}A%ƭ\�rjj�3��ƺ>���.����AA$���x���!K�5�|�Ɩ���Z>t���`s��5pE����gön���h�����ɔ���J�� ���e��F�
��L{%>7Z��eG���
��F�ZzϠw���
����.���L��_�C��-�!MuH�?&�oc_�C�&:�dt��Q��E[�W5n���*�2��$�e,�@���O�H���cݒ�����[31���~�"go�d3�(I?�׀7�)}!��V���j��z
t<A5���h�8�-�PP�5M���W@�cM5�h�`��2�>�	z|�I���ûaH��ֆFV>ih�9���z��ms7��Vu�ۉ��/�6����=��9r;u������`3���>�b	�b���u�٬F}�J�ĳ�����]ɒ��<��M�l��������gu	�tN�uj�yF.���l��z6����r�Hm_1 �	�q���M���z]aP��~.AR�?z��!'*#��+Sl�"�T��27dJ��g?�@�IQ���hc84����_����sR4���V[D��Ft��uCT��j�W쁋ը��Q��jӬ��H�]�8�
�����a��R��>`S<�8La!D�:]+�e�w׆�X����|}^�۞�����AZ1�6�5K	�N^ډ�����b�	o7ҏ���]:��R���B�]�<�H���y��=g�U��϶���8�/��j���G�L�Q��Mh��Ft��Z�4�G"�9����H��h��}��v��[���Q
)�) ��@�_hd���N0S�HT#���y�_�R�+��$��R��R�R�|�Q&9�� �����#�WRg�6y��� ��u	���ϻw.�Z3r�wQ(�^>�VC=jk�ьV1C�+~��Jt���s�:�޲QBD����S�9����-��8����G6��ݩ*u=�֓���k��?��N�,�V���4]v��~m zN7%�wҶ�5 ��a�r%���1����g�ǆ�R-
E���{�;��
r��_M>������}�b[Go�BO�0��+�^�F���wN�"�PNyi6���;�Mf��.3���}n�~���.����|TZe�N s���\��$�?�ʰ�tF���4l�HQt�ds˜"<g|]λmG��_@M�����`�<�q硴kR��>8���g�n�"t�������0�}�77)�����܎� y�C�@;�늶p�Ưa ���sEO����Twy��:@�OW'�,[A����G�G[��i_�N��{w�)[n�U/�yJ�~���t��@�N���a�Qi�3rXZ�G�R�#�~��-[�Eqy��,%�=��aƱ�o����@�kO7�����#W�JJ:w�ާ�e��s���ƾ���h����A������9�F<qe�<&ܳ��L��>��U|��7�v�^�=3�M��U �L;-���"9\t粆���q�P4g~��Z��0���W4R܃c�������E:ϳ��s����w�M�sJ&!�����j�nV'DI ���c�͔��ڪ=@]mR�V�.R��p�lY����)X�6�c��i� �"줞w��n_�59{�:G.��@�tU��E��3$�X�
a�]�H�ƛU���h�������W�zZ����#����Õ<<ৱV�Da̫g���D�џ��M���
��������}��\���=莄��"��i[S):Ma�NV�c�F���07�<p�e6�S�D\�F�[]K�)�DU��/�U?�����Ͷ]�5�� ����/�B�6�-���)!C�Љ!�̓Imso�e�*$�ɱ�-����Y|-�^�wN�&?j��*�$!��Zpj�q��g�����T�̸2��@[w�)�h[�D�~x���(+��$�6���A��N6H�3� z4?A蓙���[�E��E@F����ޓ��++�]Ft��n��]��]���� �KRX/f����y~K�Jt̓��3������
�{�8�<H�
.�%��w��;I(��9<H�#��H3	(g�����R��(䑭��S'�j;$�H���#pM������S'��/q#��������^^{���B�+X�@����o����ˢ)[����T��?C��m 2�M��XdEi.�й����,�=KX�c�AKy�r��@ـ³�i�Zs�jlc��(s3!Cw4#IH�8���a){7t,�� >���
Ē�+Ü����x�`Hݧ:W"V��
�"����9F�fO�ݭq���*�#�Nܔ�"�{�#��RI]��'�ܗ_���u/���:D_a�&��𖱶�Z.��E�%�=c�0���Z�ugJ��߶]E�t��[�od^�d���P��J��ć��M�d�g�����|���"Z��#�eB+��*�k��C``��&�/4H�h����ܫ��6|�B��@
h�z!�O07qaa8�]��:�oL}ӑ#���kv|'�-��f��V`��lz����W^J(���Z�O�,�����Ε���E$ܠO�`g,�ө�	��T�Z �o=�!�� �ǣ��L��[q���'[�pB�V(�0�[E5�#q�<�H�����"�@G��{��c��MH�tU�0�{�Xss�|r��[Leդ?�M�eD�ѕ�hIv����M���+ϒ}��d��ַ��
Ԙ󘶟�E<Z���T���b�6��iн����M�1��6�Nl�7��	���pV
(�1�2�]��z45��}���R*�fU�|n�|�U*`^X�.��:Y�|dMM�k�O;?O��"w���Uю���y�f�C�!�����_x}�Լ�� �ds9y���n}�����DM�5�}6�Bs`��kQ�5֖ l�-[�NL�wx���"�E��\���<NV �	1׻A������@D2Cfuh��(�j�&O_*G�unu�g�����Ŋ�2�/�<$:/1b��#��(A����:|~|@��{�LX��2.nd�u3�	�ڗ��"�O�;T�~��Y1�5{�F�4���	`>
�t�x����j�Z'"$N��t&GX��jZ�7�n��XRM�Z��q<S�e�0��js�9�ج��x��-	X �/��m|=�R��2�T�M��I�$�OB2�@1�s����C�.�,����fͅà�5s@Nt��#�y����_b�X$%F�ҠOa��F��
m[����O�i�ű�]�w'�91br��e ��7�t����k`Ks9��g8�ڽHA�H��۔Od�;��7ǚ)�ܣ�2%ݸ]�	�:�(2q���q���,�y^�b4CY�c<��8V�Cq��T�%��w�|Fm��#羡�2�6����!$Lg_�#��e�w2{�0qP��[����y�ci��ݭ�;�R/��s����&[��3�@��W}G�_�/��GA��D�4��o�\מ5�8\ ���s��v��|�@����o�j�u\E=�>��Ti2.�� �Mю��|�[����Їp�x�ǀ}Y�\�����W���b�n�Yl	�i���Y2r{�{IQ�9����5q)�l�K���{/��Z<t��SO'#��|_�{&5�Y?�=�pڨ�	��=���գ�#��ݴ�g.��wd��I�O��[xK`��8���1��f�,�`̿d��{�5��>	@�	Sܾ���z�P�.>n���UU0ʰ~���)-v�vm��C;,�:�����߸��c�N`�<��MY���ψ��F�)j؊���:5�P-+������K��i]�n�A�_0��v���J��z�	�'#dM�2l��Ы:��1EB~>Qk��)�v��W� +y����b��5�ۖ�TvX�Z��=��%��Ե�]�x�B���A!�m�L< ~hu�K��V�I#��� =�����
�E��Q�� ��i���M�ؤ��L؏^�̳/������V7""e��5pD�a$+�Y���%�I-�d#�^L&ZfL��!�0�_X9@l[�k�I���)�w��h]+����fs�d���_�\�寗�$T����O�|�K��b����'����l��D�����H@^�����P�[̷�w�T�hz�wxPB��Vǌ2[զ�ϲ	o�Jq���kG{��1r�6���&fE�4/�A������"�p����>�Q���B�����U"R��3�?�4�^�f#���FZ���RB�4K��!k썮���c+2��Έ^��׾H�or��&V����:4!��T�kF�P����n�Fy�[����"�D`~!c�����Z�dt@��v�(�'�B�u�}�
�,�?�����̄Ʀ��f�~�x��}�=��[��C�����8�
7%�{��Nl�Ԋ̪��z�K�r�kG�P�sǣ���Ezh7j�m�Fˈ������Φ#}�Ach�|�7�{~���ߌ�ǉ��WOy+��U۠7�ۥ�ƚ?������5��ê/��)��K�Ƭ6�̒��x@�f:���M�$��	�¾��e��rq���R@�����>���x[EnA���wL��ޘ�4��8��{���Y�0�._7�T2g�2�$t+�$�)���:Z"a��e�d.bXr�l�P��:~|C�����z.���E��O��S�NT\�Z�$ՃOR�����R��iO�8Ь d9�Փ��	TR��m���D۠7�&V���2mu{Y��6{�(�ȒԞ��˥�	�PF]
�n�U��Fq�H� �O�ǜӈd�-�64�4}��O��͘r�b;GªZ�d���5N�y:�:�O-�����Ys��;lג�ZXX{W�A:{Z�8YI��'o,8L�W�\ 6 *�E�MM8K��A�� ���>�� hmm����\�A��t��)���;! E]�1�o���
�s7�q!�FS�?��s��ў�O\Z���Z��
�*.�EE��.�AT�#���Ċu�V����+X����foBw�+�1�y���T�h�U�3
[`�dP��DޟH:g��6�RB���b�ٱy^��y�� �ޙ��#��ж	���\1�v���_�u(�������'���٘+��x�^U��~[�C%(_@'�*�付R!�H�j���՞oJ�q�i �k,�-W/�P�&LxwB��䑿��$���?9eԵ՘��@}B^�z~�V�6�����	!��	����M'��s`g�����QDǰ$~�v%w1od̴ΛC�\p��6�S"�*��`����.®Vw��Em�07�&د��)���9�6n�t��)����-Ґ�`�����^���I�.&b |��'�5;�˝��[���X��	���3�I�Sv6���!6��3�!z��,�E5-���A�����b.>����hxf�<�7��6�ȗ�]���YM���k?ِ�N��jiV�3�Ķ���xY��2H��v�	�����<����Di���mBsegTZ:F��� �#��}4���fN�aS��]�����Jh*���O�/ex:Mho8��Y�ui�^�8�+�߷��4��q�K���)�3��ƞf��2C�t�[@�_RB�|^��%�ʠ�Z��T�=ٸ�ɔ��d���Wt`����N���T0ώF3H�� |�&��	�
��B�p�Q��	N��@���PCKf��HD\}tc�Lzp5q|e{ws@`���
�C��N�HK�VF��X>���T�`+��������KӓhWCGy�i?/=S~�^d��w-�Z���}��=�0E{�������- 10Y���b��}7?��nB��{�+�_�1ސEpo�*����IE����m8�O�;R��XE�?\ ��lEig���?�q'PV�|����E���Q���op�]׽���|w��D�Eޫ�:t���,ȕ��B��W��̿-���=}�ps���."P�*u:R�Idz�{�\��;E�a,!g��N6������܏�{�n�LZԉ�"/`�,5W��û����Z�~Xf4�]�:��r�a�6���U{dے�Zn�f�+�,]�Y_RMN_7_�����͵�i�s�����~Ԟ��m�M�mQ=R�"7,�<y4x�qX�V�
�Ϋ�6�&f[A~�s��0;@���X�g|�];�!�d|Ux�0J{ZY'������Ayn�!�m�d�N䓒ͼ����m
��ڒr�B�p@]�s�����8�_=\��HW�u8�ѹG��{���f3��>�]ۖ���\%����u%Գm�p��-q̱��7@�*a�0}��zq�B�X�Bǿ�Y�m�N��������t�*Nd^�ݫVN�a8�0�2rR���B�0����e\���)<���D����d�]²�]�E��1�>D�4e�	��̞��9Xv���`K��fS0�pɰ4���M�E]�[�X"�P��F����$�g�Ħ����m	�➪����0�*$5D�|�S,׻_�YѪ!Ƭ��T��q���Â�C�=T]o�#d�'�m���&&�S�`KA�n� ;�P���\=�V-��%ZMߙ14����c(��O�ǥD�dБWT&��H5�2�9���~J3���c�����)�t��*����V�L��U%<�7��v�h�w��m��yi��iF24N����v�?c�B�1�bެ�4���wsn >e�o�46��}��]YG�$텓:�;���P�ϒ2`�{̵š�& ���Z��x���װ��
vu��a̣GSi�G��x?��< q�ʇ��f
�PXFS0�_�O���%�2��r�fY�h1�Y��j��|t�$�r5��Wc&��P�iC
o�����m��>t��vG�U�����'�ޗ_md54��O��aC�"z3�.%��oGT��Y�u����xL~��ʃ�"�vd�N���l�F��3}ޜWd1�y���:��P��4N�F�׺���Q}F��o���`J�"��Y� �e��:����I��l쾟�P��>�8G��p��¥�G`{����:�:�?}��N�Gܾ���|o�I�bF�k��Q���1��<�X-Y��H`J�7O']�=�fs�xqW�.rI2i�]���Vi��n�D3���"~,n���P�
���Fx��cN��%���&D���%n���bHC�4v�_]�ժ���]~y�0��9���^�:�\3!�( ��d��D1w��wOE��V9���߰�1b͘���^x�L�Vu�.���V��g�JC,�n-�����'��h�ok��>��3�sH�o� ���yb��n+V5�s�c\��w��xY��ޑGޱ�'ѷ�^O"� Rm��-	Y��s�R�0�%���ć�)�թ._^�gO�7����*ȋ�^��.L=�P� 4�lQ�G�	�1���3�JQEF�D�u�b�8*��4�����3�S�&����rq�0�_jV���c<�2A%�'�y$�,������<&1�VI���}���]�6NR��m7�-�
����F
��]p<�P�pC����;A�YE�&��f
�$���s:��^�!$���3d���ae�@dS<v`���`	~�j/�
ӧl �+'�,�l$L��<�4�i�o�q�*�DW	K �n��R�\)lf���2����قM�U�:j��v�1��;�8��&`�����]�mb�����f3 P��{�Z`��I��Jk�nH 9�o/��N��@.�;�����z��� ԓ k���
O�\N�I�K�x�J�+�c_�
��l̕+�d /\b�[~�Է�G�T�w�sM�ng���W�:%J�T��Ѽ7ċ�'_mGRIT����o����cK� �%G��J��X��<�ܟ�+��e�k���-�d�^�s�qλ�Pl����c�P���y�����p��Q���&����!A`��B���v�R��dD�/�`ũl�x�~Z���|���]i�"�Ru��:~ړ�7���=a���ͺa�6�x�ӳ��Ą�����%���Г�Vn���ɶ�WF�C��1AL��r�۾��iCX�	-�Lgχ6��cf�}� ���k�ΠJh�vR�Ԣpq�8]�H���!Zl�N+n�Ʉ/�>l��!І��h�i�H�YG��hri��D��?Ŏh�n�X���tO��m��n~sQ^�Ժ��k�O
Y��ۥ0�ボI�	`���Q��	W�)�,����[<v7J�q�X�M\�ɵ܎�ݠu0��8N�������9,�٣\qx�B�$��9QR�<�UP����T2��iu�����hL#n��6�F}t�gx�-Jg�qωX�^.�p�C������?`]�����2���;*���l4�^I����b�au�R7��^�6�̈́><�4�Xf'�&����YU�/�W�iP�C_�=b3��F��Ӊu�����q]o�`~������W�-����z�F1���G/̞�t��bT���\�֕B&�A�6�� u��=���U��l�s/_��"ځ6�F4��x�?:��<=�jӻ:Ph� `C똝ǈ��Why����'yN%���S�ו��i����8Q�px�F����Jk���n��'<,����#�"��L�R;�pp��:/��$�⮍�i��q��Ɓ��[�����F��?0�b���鎺T��A�JJ��u�� �2_�P�ƼhA�����u������d���b���~����}?�R�
���8��O�p�X=��`ԊU|���\�Z/�4?�r����A�p�WK�k��(q[�Lt�R��#����V��}���Ϡ�mE��dLj\t��&�L�-�T~�&��f,�W�2$覘<� �9�:�����=�!�Ư2����MOhj�sÐ�PCKR�@�m��(�
��<g�m�BF�.|	��g�s�D��j|��\9���
y`��Ua�eP5ݿۇtX����F$��70�Q�;	îŲb�5vsbCy�r7;ܔʜ�qa*�y�V�iAU�<ك��>ݮ_�Y������JP����<�6�� �~��Td������=g��.�y��L�B!k3j߹�8X�L���'-c�m���!uo_�%瞜�b�������6����rA3.�Q}x�"�Lqg��*����S���n����#2��s�>���e�\8O���|�eyt �fl�g�RWåMsT�u��u!ՄA]�@sɧ��Tl�ׂ�8|Є﹯�
~��#��C�ҹ�!̛���<�a��1�|�,�ͨʶ�wg��;������4���ر9�\���/W�
��d�w/Q%}V��(|�����ؾy'C��M��k3PB��Q*Ů����QI�46��9&�TU2��μZb�=����A��s���>ݺ~��_Q�mЄ�ላ6�aÃI����h��**#��J*6�e�*��I�9����L���nzv8�KX�z��D���k
cS��+��x3 ؔ**l �x�����e�o;�QM�p47GfF��zu�D,b�|�KG0��C�J�,�0�$��S.�����c���u"H�x'P�(6=��ٸ'~���*�?�A�Jx�����߰vs�Q�^%�K#/_�����a��gx��B�3�ȗ���9��#Dj��IQ�x��D�6��fgӆۢ'a�g[�$��H]b��6�K�|Y�dkXZL�q��WtF1�^�,�b?z�����}Y��w�	([2ׂ��1���W tݝ��R3�նJfb�U��SOgJ��f� x�iE�DnX�/��<�v	�wc��K	�μ��ħ�y�§�Ɔns���3��1����/�/Ѣ��I��a�d��4&vL[�V#`.�z���P�7�
ҝ�	�V�����Ö�M���؇e_q��_{z���1y/��neӠI����B��$>�h�t����1�t��E$;�|#�(�V���%jt��BcU?��_-p�_�i����Y,Z���x�(����Bl�`�B���A�����Y}���t���<�U�gv��p���R�uש�h�������ZBL��	a��x?�$Юźr��|�,��]1|JRo�����MG��J���Ŧf6#!��:�Y;	�l�O�SbQ!��;��?��X��E��
�ڪ�EJ)�㽜l�6R��X+<{���hw�kE�Y���:3�Z\�s�c�� �[*�և���9��uy��
�IL�K�9�����P�C�����>.��L��P�K��7�ۗ(����@�*P�'���6�s8]t���P/���O��\���m�4<�u�I�L�x������9W�M��B\�������dw։�#>յϾ�q~]�11L5|���Er%���n�H��϶������rӼ�n��l����"od�(��2.�qS�GZq	��fNo�ѝ>l�~�0����u��B��c��{Y���P���_d�J�zW���c�⑗��8���ԶP-�F�jyVMXg\�8Y�މn�݂�,���;*��δD4Gju+�dt��隅�!F�S���l'-y4��[��;`����e�1���Av��r�ګW ��=!HL�ց��������{
rp�&{��t
���XO����]�X����;DWv�=�cìC�/Y�l-TK�A��b����LƩH� Om�ҤP ߏ��wXfƶ��m��
y��:F�:�m��PC6�[���
>�:�.a�5��ڔ�c�8rh��YX��5q�����/!8�cQ2�M6 ��MƝ,��h?K?vd3o���m��<Y�DJkg9���#�zB
^���\�K�|����: v;���2�$ߺ ���$իμ�w� � ,��5���:�a���
]�ґ(��t^pU2���y��:�F��ͩ�2�=���lX����X-<c`Q6{���H������	���Ps�F�~! ��7SS`�,��%q�;�5�C��/���:�2;NJ��R��ɑK�a�?�d�\zx��'��˼��u�`�s�d�_o��4��q�F��֤tUDgH#}�y��"�񉵗몢^NY�ׯ-�}{���ġLk�t�Jj��\�R@'HP�'�N�ǝo�C�N��5����?��)�;�ç�e�����}�O��H[���ľ��vp�^�F]��Q6-�D-*�؆
���#����$����,����$�wi���<��=�L�놴_�G����E�Pk�b�0�׺�X�y��|��g ��B9��X�H,�D�Baf-���u����3l8;pe��P0*k�<�T�:���ˎ@4�g +��phi�B���+В��t��JF�����3q����r¤wIx��,Ǜ���.�Ư<+ Y�hi,[#��� #�&Fb&�	��;�U�a�h����e�<��������҂~k:��Σ
B��X���H��K�="����L���m����� h�	R���Ū��T<��r����h.=n��j'��շ�P���QЃDy��﹙ Eo ��Ǘ�Bɤ��燳�.p���m�����bڅ�h㋠8��L�)\��.�ǋ��0BU��ad�tG?=H{Y5��\�'�PgQ�<�����'j�J���XD[�z�������"��-+��J��_e�I�_7LV?g3X�I+�F�r[��]�k!��xsҳ@Ӎ���*:��Γ���GQ�V3�0�*e&�D3Ia)-��[]��!p�us�3���������f|m�b5U�������f�'��0��Z0����G��s�V��{������1Kg��a�����o�}�}�Y69zm0�]���ʵ�.�q}�z�!��[s����v���,�|H_#� QNl��j�ԅ���^Ƒ�ݻ�G��aZ��`��f�V�I�=�s>�WDq!:]�yow�G<>Oِ�/����!.����2d-����ʸ�(N}��~&:HX����N�$��%9;�4�N�7+��Q��P~����*����v�DF����򠅥d�D�1����FL@�n��M7�0���KE{{��(����7?-��14��w}�}��u�V�HFu9�E)7:0,����LU_�	����fMe�����c%m����H\§��D�b�x��j\/��3�A��m l�dx�-��޽��V��T)�iE��ݾΨ���ҡ���2�I�\�����>w.�4�E���;�?:Zg%T� �}��zf$&�j^�����Pvs*��UY�!�;��\���zc���G�GD�?�p3�d����
(������Q� ��i�	�(�'������QmM���Yh�E�)��d+�O�e^AA�2X��e���kI�K0�+	0���,�8�w����6�E7�F��ƕ��rD{�^.����53�%8?)�x_;o���G���M��]���-��+oF�z�C�&]���J���Ur�;�	{#b����4���݋<�h�/[_��a[�Ը?�wA�ֵp/�h�1!۷�m�K'lX���=�����,�h.e)��!̭#'��7+�w�ɔ{Y,���?��W,�Z�����0� �}x���f,(�/Bԁ������7��ǰ�,�ݘ�a����n��>y� �#r�ʣ�)���t�n�U�����Yy�����i�-~�a��	 �<��w3������5+�� F���	K0�vY9A��B7
�_終c���va�u��ԓV[4E!�N�dtGB]��na;�+��_�bt_A-D|�S���v�ʡӈ���S�?���҈  ��`�V�����r.�8	��9�K6[�&X�"��"AG����yǎ�}�_2�g��X?�D��+&�E� � ��;�litN��5F����E�}Jet��������1��t�c#�9�ۣ�%����ZlB:��ݔJ�qZA��Dc�;*2��O{�<b˂�mt�����Գ� w��\F;Q6v�O1�3$�����W���`;�P���~3u�N@JJ�	�+���+��:R�r�͵k?Y���*+D���V��~BY���'>��	�����bY���)����QG3��ҋ,�7����W���`oO����2g�w@6��|����&O�S��ۉ���G���^�{���r��t���5=�y�}((����LQ�DK0�+�o�ϭ�F��)5`nE�D���n$�P"�*N��/�8_<��!���V�C��O���c��\K�b�/�rd�� kG{��m�H���v�F�M�U�;��R/�`5���r(],�X��xE���9\�]Ҷ�=8_`�>())�t�hp��+GkD�(���J�'��Ok�k[����D�Fn�T���"�^C�R���#���/p�Z������{AK`�L4q�W� ~�r�a���J��{(	�	q��LP;ZJ�_-���|� �(a y�Hg�ǩ��J�5&�*���,I_�Ÿs*m�`�ÉY�|w�6�� HK�s�@�2�b��ф%�:_n�ѱ�)YǝR�$+h��Rۍ*tv��nhB�B��B9t M�S���v:��+�NU��|�����ف(�#���Ō_�h�fp� 4L�w��6��-Rڙ��Gn�5̡$zHL��bz!�n���W:��S����=S��c��pSZ���I-W�`�&�d�_��7���J�)@�Q�!�I���QAg\�n�/�t��`����(5���5��nW7��'_�M����^���=��@�}\G��Q��J��&�W���� ,eP�=V5TC�:U��v(fk�F����uf�c���ؕ��K�uͷR�Wx_ j��7�T��pMxu�(spa�3�ć�zM���L���I�k#z�/G`����-ܰ�ql
Y�� r2�	��@JZ�?4��ޢt�#�]q�T���S.�Ld��b<:Y���M��+l;j�c�L�L�:p�}�����1�_@G�V~�<U�08��;��}=lw��!�#��
�5s\�[��g��-��W0�5T�=�o�z텳Α��(w��"4V)��mK�;0?�~i��{p`���2�T�2o>)�
-iME�����X+e�q�gx�B�o%���F�9��ʕ�b�D��cԺ��(�I�1Ӡ�x�5�ߘ����e#��&W{�z�Wq�RC��/R�l��ܞ�7z��
ל��s}��~�-��y�J2�ʝ%��J0����o��[r��ԥy*ҷ��TPl߇��
Z���I�+O"�_M��8� P ��(�\��F�9[�sf�6���ߘB��L��2{6�
��:T�d�9l��h�7KJ,�u�uh����ԾX�a7Qm�"�Y�~�?*<�E��Q�_�nPZt��n ��d��!�j�`���b"yO7N��n"$��Ll_�!�S���?��-�sV�k|V��0��b�y�U��%�6���wR�����$��{�ѽ�<s���F�~)�fZ2����,/08آ��>\JΆo�6�>���vd�2���?"
�^�!����DF��c=�ISG����B+�f47�u|�]?����!�L2.�����|����Y���V���+�XL�g�89���X;��ƫ�S/W"�.�.:��l��v�Ŷe]U��g҈��qX�g(��ͯ|�ǽr}��R;!7��?^�4/���#��lဎ=ap�!�ҹ�� �3ˉ���6Z;l�������T�@����~)k�,(�l��YV��5Q�P5D�(nx��D_�ʠٝ����L�1�,߰�%�xT>Ff��=��J� �b^.��	,r�(S؈`�E��X�$���)d��tv�y-��B�r7��J�����uP��y"����5!8!����G㑣��S��͚��؉߯��pN�#���@
H���}ѭ���<Wۆ>7]$S�B�����h���Y/f9��s�����
�s�2�`�|1�g@����Ǽ}��4#M^!��;��t�I�R��e�*�a�2Q�ٺD��y�����C)�z�^^(J�{�����Ґl�[�f��"̙$��^5�/t�Lqf�==��8�O�G�5�Տ �v�C㶊�>�'�e
��^�Bg�d��|Q%Q�=��Q:���A��r�3��:bl�_�O=�~�d˲�Z���pi�、��}��l,-�HJYa&~��[g쥃�ij�g7Ӈ.�!K1F��dm�W������M�r�`�X!������2��\���S��q�q�$�>��M��5�Y.b}X�ހ|:�{<�"���B�q�)u?�Wsb*��h�
zf����U�es������'4\2[��l�rCL[)�?�0�ȱ�?���X=�M��?Q�z)��k;�P&�B�]2�D#.��0d��xT�d�g�E���C�T�����mk%�z�r�Q4L p}�����%S��Y9�sY�P��'�q�׋��(� G0�D�Yw#ڇ��J"X$��q�.0��''��Zc��Å�#%�!E���wA����؉0�.��Ṧ��Mp@tF]�tU!���׫�3W&9Y��C"�޲��<5$*�Mw�-f)	ܿ��Q�Z;�Z�h|�ϲ'�*��r�$ޣ�?X�<P<��飳/2魠S�l�}6�~��g{¨y��@���}_
N��B]��!�9 ?�+��p.<b��yZ�CŰ��͹Y���g7P:oE��qm�:8;c��1�2�"�Nlp�ߐ!q��$k��@{3*��69����� ����m/����d4�W�������Xe��z�ƪ�_�m�`Lv�Y�t?���PϏ&R�DJ�k��5'���v������eb�4ưG�x�p�X�YrjN�"���"��a���h^x����������J�"/^�Y���E�F�{x\�x� C�J�^��T��|���/٫n��Z9��Ra"�>�:�\CNm�Y��4�7.e����	R�!���K�Sqdy�XD�#��=�db�V<F[�K�%�������`E��d�M��#I0D� ��D�'_��,����5��Vg�q=�L�n��y�]c��5۱�R�4 8E�h)��1LU��2ȸ�����
������Wz��Hh-�j�Zs��L^Y���?�V`��(�[P+�G����5f��
5D�ϣ�*�X�B%'�0���\�d'�:u���D����`&�1����a�q0��>cY"��M����������z�{]�Ҫ4�2�5��ɝ����n�q����e}�������P��!��kU^F�k�X=J͕e)����J�ѷ�7�A��}��e��R	�͑��rG�uW[�>���d{v�_�'��Z�{��%�qxf����A�tpYG/�q�+
J(����sn�ܻ�7��icr��tv��s�J�v�W��9^Hk��Z�OO��oM��53�x%����b�6�I�-�_�)���a�W`g
>��A���.��E�%Q���Y���6 ����ր�3�U���VHh"� ���9�8�E
,Bi:�\����Tq`E��[ˬ�[{��ynz�˔m�P4&�'0T�z,�=x&Ř�b�+D�PwQx��,��'rD��.%��O�z!��Tf���$�g����!ۮ��M���],����/p$#if�N�p��O��`ɗ,l�k�007���j@v�*�'�$��~m���)�C	������X��~�0KWA	���=:a:��y����
r4��`�Ƒ
�ƺ0��3܍��X�l�{4��I�um]���iZ_�R�(p	`�h@��&�x#k8S�����g�b>�����\�e���	c���;[���X�aB}a��c�Xu��>D���#OԒ����%��F�r����Gn3�����.kh�U/*B��ҮQI�b�@Ϸ� DOsU�%1����i`㋟`���ԉ-��g���fɞ�Nq9D��JK5����S�U���F{� �,��h�mɯ`3�< w��E����wUht�?G��F����q�'1�S�r����:��H�3q�p��?�?� 㮡o<�[����e�0�I� 8������jGu��関~�W��Z?���O���{���5Z���Z ~2.�,f����+3?,j ��Q��V�d��T���8���4��}*�����¢�y�������#�D��8��w�:�ZT���jYj|�ɞ5������9I����|��'���xN���z v��G��,@�|T�.svzu��k�PL�S�6��U� ���O?p?��%��J�߅�MK�POY��_�3sW� �%��>,o�e���w��h��Rp�W"
v��U���;����g�̈́=�a��۪m%�=��Q�[�D�\����c4/ 5�ng�~>W��{:�:� 4uKrlW%��C��'�w�˱w4������������JA��þˋ��-Y1s��\y蛝�c��\Ć�N�]�n_�����1��9t������e��z��`�'�[���J>��ڔW��s`�>�\����Q5Zf�$YM�<�[�����P)���<}�f/��E@�z��:`.B/|���Q����yͻc��Yc��e��q��#ge��5���&��|ģë�'��26C���'Vt!�C���g��&MH��=T	$�W��3�b��%k��q#�B�j���Z?��餅���i0J�UOcb:�re��s�rK.I��R���=�;v������׏M��o0�L���yD���̭
6x�N4ڢpI��I�.�"-��d{P��'���۲2�m�\s�싸���@�*~q���_|��h�Tpo�?��Ƭ��Xa j�B#!���o!��)��h:��;eM�:��Y�����������.����p���/<�)�:Xcg7�)m���t͞Tdq�sDp�D*���B�˺����~�����8� y����������ұ�5�^������4��(�nA	�Z^):iwh��ݘ��8��{79�Ǳ����l�쉠`C�h�"�Ц��7ɂ���[_�Hk��C"n!�-�|z_R��U��X�st/��,�9�����]=67�zf5R��l�� ��'P:��m�N�*���^n'������RRG]�)�E$[����E��"��}�M'1�_#���!$��L�ck����Ї}le˓B�fE��u�B������W��i�'�:�1\@4¨6�a�cv��G��������T��R�P?�	�|D�"��Bנߞ7�i�VK���ۤ/�:�^�J9�YN�����4',�����E��u#�lÒC�a\�`l0�}+��>q��������<��Y4Bꝸ�<�5���L��(a�dU�0�N�K�4UU���hO�O��ܤ�K2)& d��TI��xf��A������dNN_1���wɿp+�~J6(� ѕ�_-Aj�p���
*V�WvRz"���C6�?|�>�śz��ZA�c���Q��֡���p��6W�m\kHe��436�#mP�Rk&&r\�7v�ɷ�S�^��G��`�	�Ɉ�XAf0{���.ia�!��>�c6d��x�ԣ9�	��34{o�����y��d�z�?^d�Q�m�$1M��yN+�����!V�nt�.z���KT��xB��*����kfz|i.\�_�Pѓ�P�p W�q��g��V�P�"�U_�SR�4��.m��)� 
/��'�|[�װ�c�I�gB��fp"��v�H���0JΞ-4��-+���y|~X-��톎�#�604�U���MX<+�MC]����9GK5�5� #�� X�wΐ��8>�+���*��s�^3aM]5CJ�m�{��\�Mw}�^
�`�����|�	�����6����^K��{�N�]P�>�R�9�,}�|ߒq�3��z��aB6�[�`L)����W�p�%��N=����VK�U�m}K2����1��Ş�(�WR�,��*��j�P��Я�~��V��C [��t*���r�5�{�ѼP��"�" ����,(=���Y�K�G�:
�ʭWݜZ��o���}1>'�����Yn���|~��ns��*� u�:r%���\��i3�h���QĖ�{��G�9 ��;l⮮p��:���Q�Аx�6��pB��U��"��v�"���R���Hnҭ�U�5�2Yo%wy ���<#}��B��aCm¯)�2[��J����Ս�#rS]��\�-�(����9��K6_QW�a��o	@�kG�lL��,J|nr(&d���-(��$B�R��L��8����#r��(�%Ub�8<V(��]�0fP6�D.���ž�~Yrś�N�@EKc,�?k�0��Α�xh]qs\�':޲�s
���yu�<
�"�wN!��	~�TO�X�m�8P$@X�E�1;��]4�GG���j9���>c:�SUjrT�>�$]ϙc&j�aߺ�'*��ȴݵǽ�C^���[��:q�Z�5!�Gc�1WP���u�}�����gۺ��煀o�a+1z�¼��O1�W�ʖ�$]�a�f�����|0�70{���o3k��� ���^��s�dU?��{�C�,ox��MrۗL��� ��;�9����}>�嫏�68�;E���~97h!��i���ʭN���fx���K���pv� �i�#Z��՝�Ǌ�9����9F�yA5am�~��بC�\&��I*�j�MǼ�/������}IɀV-���IvW��N3��(�Q;��"���?�'l8}!Q��P�����T��K�������ǴBi���^�l4�u1�o�G��i��8�9�g:���J�V�r?x<;�%�9^��S��Q8�,D����\jo��~2̡ >�6�L�TZ�Ft� fj�9��e�gJ�H�ͼJ2��~U��`����|f�-a���F�_b7�Ů6�i�̎�ScّYw>��W��f?GO3"[*?"�����ZD�[P}��p��	"wC��H��t���c�7t�O㘅Y%������[���f�g��B4[���s�9R�Ɩ���X� ��!^�ظ���t�p�ZK�3�Fe��븩TP	3�K�rڠf��[���%�v) �僄}����.�G^�+��3�Rz����H��d~
�)��F�%\�G�%�ʎ�߮ݝ� f��������6���u({B�k��!	���_�O��|�3^8m����22۽���r�\<�F*}�eJN��g����v�R}9��I�<���r��mNK?���?1��i��C<E�<����� 5�]�T��{��߳���]���CM^:A��w�w~>����0�a�'J=I�d?�����KºC��e�Vٮ�lA��e�:�lL 6ߠ(;�\PA �U��ߋ3��vl��r�r6�C@��?�7��,�.���sAmϭ�?P2q/���\u>[zbKR��qE�?�c/:2�
ie�1P�HA���
�Fd�OE�(n�\����)��p��V /g�2�v�_��z�4w��G��1��(���	�f����b2�c=��Aw�ub+��Sd�-��2����Z�DG��}�%?�+���jB�z*���!�t�Ӡ��<i�����?��yѓ�,F`׵�c�R^­�<�7I���e&-^�Nz�)8��=�K�6�a�2����		C�᷼׼�H�B�
@�%�[O��p|��;�Km�I��lD�� ��A�B�GF�6��?�����H�k��t�8�?=��E�|nH8��f��}�|oo�"f�@Elb�$b5 I�?�ʗ�_��wV2��`�`��C��+bҕ�l��k����zC-^r�M�z�l�j�R7�d��`/��#�tQw$T�� T���6
��^�(�SN;���=,w�efnl؉p,��������Q���@���p�9<�YP�ڛk���5x�Y�~Sqw�&I?N܀��r�L�5U�dvԔM{y��W6��!���$>��A�H��w�\��Y>��9x�U@Z��т�&*�G0!k� W��-������D�K�9�:��CtK3&Xn�$��淖���m���2�p�ء���"��ٚ���o�Ҁʻ�@sB9dY�&ч:%�8V\�`�p���~�������)%�r��
�S�A�(�*��ɞ���£�P�)rܧ�&�	��,�N6a~ֶ��}j#_��Y8!w��|� >�d{��ǭٸ^b�;��ZJ�����+�o�\(������~��?1�5�J� =E�����ߣO|���Hȗcl��C�7T�*���ٗ�ײ¦�x;�#p����^��su��#��R7Ӹ�x��+��y����i*|࿀�@W	K���Pе��=��B�A6OL�P<c�62��9���~���܊��Н�v�$b�����y���m�hYʠC�r_�����<-f�Y�)��hX]�Lp�8��E����t��C��V>Wi!^!� �J��$�ϭ��E��W����	-X$��o��H�2��㙍�㦶��M�]Z�v�k-��n�Eƶ��{���� �V���eߔ���]�5�]
b��MDT��0��W�F@!m3D��b�l'Ü��M�A�_��L���%�&O}r� <�����v����{4��j\6̊��:b��5_�kEd3(��u�-��q�%?6� ����$5��)?a��}�����v�ΈС^�����h86���S�K��*x�r��$Fno
(�%��>����z#U*ϡ�Ҭ� �fK>o�z#�T��	f�ߓ@����w�Y�k��b&:���<��uK�1,42���~����� ��ӷ�VQ�
9L鲸��f~t�o���06�9S��[���uȝq[�Ȱ;Z��.w"Dp(�
�l���u��[�6xw}:C�,�ki�3	��J���f���M�9�=�"(��Qc�6��f�p��|��kC������00����d�`xٕ��ǖKh��c�=F�0V*�\����I6����G�:2 BÄ�Y�N֊�`��r'v$p�^J��_���w�&M(4��,g��΃��v+�B���;�*7!�V�Xq�}���A	#�d�S^��x�< O�t
h�������JkD�X.�i\��w��e�ᎹuY�C�G=U��BO����>;�2��&�h�u��B2���c��v$޷�&z�"Q�gN���Y
�M��S�#�\]&�<�l���l���0���}^ΉدL~�s(�QI<�qn#xt�!�� ��?�w�!d��N��&���H�F��Q�/h�$X�F��C�q�׌2����\M�$@��E� z�S�d����15Ǥ� ���ށ����o�cl1˦oZ�ps0��ծd���k���s?$�zI�n�'iw�Z�+���%]�����̘��_W��D��gvNT��BX�.�l��R��[mD���&�q]Br���ͿI��Y$��n	3�*z<��%x����t�Ka��ٰFx�-�f�¾8	u��~���:�dm��{�9��������"'��$�e� \��AN��m8�>; �g��|ͤ$tY�1ǌ3Ͽ�)���HR��������ycBIh�=�:i<��M����}�eJ�I�~e��ь%1�[�}�)qHA�5BF-���=+a_^�n��8�D��4).��,:l���
���ң����F3�?�^����8��P��ǖñ��[[w�˜�o�U~h�^�m��J�#
`"���+��w.<L�J��Z��}xj��������7�+f5����`�;����X���6�I�ħJ�C�*_6�_Ϛ�_% ��Rb�C���VN�_2f��`@R���9a�,�_�n�c�����y�d*�4��ޮ���ms��Q:+�������߽�	e��ڬ���[����ٰ�򱵺��V�#u�(�X����}�N��9�w�JVc���Y��=L����d	9t�J�'�Z�R��+�Zb`k�[k n۝ߚ���<� r�;��L_�5%%{���"����n�]Hl�?�й��G"��g\w@\�e�l��<�?��pi�����]�;*?��~���05�Y� $�^:�� ���D^���~l��h����������G8�غ9	��ȿZ�Ö�Ѐӷ��0�g�,p���YYU�R��^<�����Z1K<�g�%�00Zu?�Lr�����#��6~@��ɮP]`��Q�x�J��!S.8�{����K�{���Gq�/�3�0�_q��cg����e��
�[��<#p���tT����],�1�h�Wߙg��D�2���L1��V�;-��K�1��,�Y�K9�?t�Q(�Ǽh��a�vng�,�r�H��X���S�����vUG���3�J�4�m!/_��oN������!��0	��(���̨ONc�2�^ڜ�v���d���FV� ���E�����Ѱ8�I>��e��q�f`��29y�;�t�'4�J��w<U̐����i��l�n7��y.@0ʞ��}/�h�@�V��&
��.\<a�����G�8,��.W�'
�����g� M���I/�خ�	`�aپG�*"2u��>/E�	���s`� Y!�v%������>:�*�2�������%�$xp�ؖ�L���
Z����cpQ���ġėቦ�ĳ��1���7+�8k��L�'?�i[���M#�yr,�
qn:Q���Un.�Ŷ|��IM��
�Wx_@ �����AR&�g�*������{���o< g�w�}���9g�㘅�T%��6��w��4i���OsPg������fXh4��Ypڄ�D����M��`D���_S��������M�D�{.)���}_�4�J�w�Z߀��G�S��6(�w����)`�s�����~Sy��遣q�_`b*�ULh%�0Y��B�/11;�8�'��m?3�]^��<W���b�=�ۊ�q�~�ϴ[���;3:������S�hE�[��{f���P-+��'�gVf�}��9�� لh!�͈����j����A��&��hָ�[gh��b�g,�8]�j�E�5�wr7+c�$[p��x#����O���8�F����R���<����'n����jk�6��`ZT��:u�ܻ�����pf�|o5�G\����qU~`���Q��(�У�8V��(8">Z�N�h�z_�-н�>�7����_�s^[f^R��"y����0+�x�K�׬�k�z$��Nl�������%|{����.t
�ūY ���n��P*\k}�A`'Kՙ4��=����-��dx�H2�ebF����Kl0�} s�	����d�,\��%$��H0��_�@�}i�{H�)/��C{��>���8�c�B��s���4�}#f!�_�*���ֻ�Id\:-@���Q ��b�67�\C'�]�5ܫ�b�e=1����"��
9��b��ha�.F��i��ø�`�N�x/��&��@�����4<����H���2���w�>[:f!�8Q/?cW+�l��_��0Y�����(��!�8o��B�ZW#ی��u¡-��$�*[���LL"��x�0���6)�ĩg�y}�i�c+�r���Ms�C}��"�y�4�7϶\\ظ���A�ߔ�&��z�,�ߤΡ�F>�)U��0�Z����4-��أ6��i�������q%�0��s58�WrO�|~yC!N,Vi�Zc����R�[S��e�i�R󅺐S� ��d������Z�eb����#����(�&�0�##����96�$l٭t$�����+K~�(��"*�y ��H�}F���f]!�*\yD�=� �e7H |���Z�lĝ��6����n=�>� �J�Vц���5�,��M>L��+�P�{��r�:�����u��Gm���K�8z�Na|����e��<^B��Hq'hYǊ�3s�-���ȂH����,X��v�9nE�ש��a�B�w�al3n�A }�0�	�����7�d����UQ(��ٽm�^�:�J������r�gC��cq�v�XF�sj�t��rt	̩�7���b3��p��ͧr���Z�m���7}��VL��@ξK��Gը˘������ñ`̊0��拵�ΰ���0bp^O�A4�ZU�����X�Ƥ�n��<<4�y�8/��Ȕ����.�WB�2>Y�?�/}m����Q��j������=m
�
z�R{|nhc͋����$(��ݏ�vO�Dm>�6o6���v�F	���k��R�EI��t1��F��C���5��!��檭�'w/��wޏL2��r�]�J G�BgJaPŪ4���P�3�<��Țo�u��wO��w9?�Y>� ���E�H֧��Ͼ0�,�c�y����	������F����Ud�ςm²��d+��J�C��L��B��Y\�QF\U�C@�Ux����^����kY�̨n^��ZZ�t�����%�Rw#:Փ�������u���?�_�A�?QDp/�n"�qn����e��{��M�A�S���#�oa���MMMP�fl���;�`�?;5�J] P���'CU���ݓh��͔�?�,�Zh�]vD az��2��#HȲ�b�\�������RK����/����D��c�9�ְ79�sk=ë*��1N���R��$�=�����������Aј�8~��F�+��rN0�e�Y�<%��.n��˱���@���*�����X`�9H�f�QG��]�n�v%
�����X�k���i(���+�)�V����L��ߚDqs�.�ޤ��x�#�U3��)����Q�_b��c�>�)τ�b��p,�SD�(����s:��{&z0��82�O�i��]�;rtoM??`̒�.� *ؔN�+��:3�O���w�QN��<B�8�);�� ��~y�ǉ����hby���-�ۿ� ��V��n&X~U�<=��i���P��A�R*�kH)��=�ܜ��PB��U��O�h�R7�M%�^��0�Ҩd����-u���J�խx��	�yQ/�T\Zm�gMɴ�fd<��e����5�-�����Ո���XO���WK�ƺ�R�<�Y7���ج��2b\>=�\w��Oc?����.3����upcj�L���)�G�$�,n�X���4چy"�1?���W��!��%S����JO>��"t��,�~.M���[A�mZB��R$am�Hؙ���+c9�yS6ē�1G<J������~;Uĝ+x�� 	�;/�?_aL(�O��&�i�ƹ�UN�Ť��4�����_�sޖ̇I�E���_Y2����k�i�=W��2���g0	��r��n.5���Je �F�a`�bV���*���%�x����i,�P���VGRb���@vt�5ĵح�`}�V}��m>&w��I1of��sV�����>;*��G�;��Ə ��tF�M�Q�-�N�Z�=ٛ�|k:E'���Gu�.g�0���c���v4��q�����/�����,7�2���u����k_�yG��/�����Q���c���ǔ۾!���$��cg��?g*y�����b�F�#�q[L�?G�BN� N�בs�[W~���T�9)S�S�������J�n����il���J���fA�A���ep�(�a�8�6G��i��Wp�I�#��A��s�T�Z�Zs�ʩ��%����5��[�i�J��Rk�C8Oa����x��C#�.jC��*�ة+����:i��җd����g.]�a�yȤ9�\0��Y%�ʢ<�	�,����Y˪�u-��\��c3YYބ�=��LW�Ӕ��q��q0�L�l�xѺ(�y�M�L���!4Ӧ���g����o�[d;M|o�-��y6��gܧ	�=���2�.a��Ol�ք��Y��>�n�9l���^6��e�������,Pe�1��.�讀��h�`ށq/MQ�E���"��BH���h��%��X?X���Uc�U@�rx��ꂪ�����KK�H���]�8�Nov\������q͛�}�ӳY�T��\��c�Z���Vz�Æ��9^>��� ��ƿz�>�b�Ju}c�:�>{Ꜭ�e>$jm�mj#�Y H�sDF�:S>�l�,���EP����gq&��ȝv!��	��{hd�!𲚎�����Ӵ�wp��LҌc�چ�v|��x��9��@ Agw��L������h�t���>L�t�ĀEl�|��`�������䙵�,�Ʊ"L��0g����������q܍�?����xVϩX��L��G�V,� �9BFf�mD	u��f'M�2��5-ڻ�g�M�!d�zRG�O#6<�[ʉ%�\`J�q��A�g>�%9��?��=�A=��9CY�r��M��7z���hBE`�a�B��o��lv=�ʽ��(~��U��v��� ��n�H�ПUJ%mbQ�QE4��5�RZچ�5~�)�y�zt��݋*���=�5 @�'�����1��˞�n������ѷ���]-z����b�M��a�����Σ���ɬ��e�V��q�����7[����Q��l��&�U��;�����<F�����媳��d\����s^V�GN?0��H^���.m��W�톞�����a���ɷ��q>A^��Լ��+Ѩ�p�L��k+M)����k�'��m�r_�*%s	R$]W≎��7�a���䤗��)����*d�5E&A�v��J"�dOv�����R���'���`�C6������ej��l{p���ϝ�����"na�����ԑF�0ຎ�����B��{��'�;#�s#��5�#G��R�nK�������V֍o��'6v9x�����9?�nNBހX@S70O`����	V���N{]\��HߔD�������R�v����T�����Ao_��d��ob�,C�6���,P���5�.�W��M>u�e@8�MʅG��n�[Oz�I��.�HB;��~�,Z�+�z�~ܸ�~K+A��}�}��,�|�5˗3%����5cs��5���(��s�F�l"���8K���%ȯ:'�	�Ǎ9������;Vi
d���1>b�5��+��Ջ6O�>;�ݺO�M���@����p�vCFg(�,�c�~��|F��Ҏ��
�Rp�����W`0'�B`/W�72Q��2��~t�B+�4�}Eg7����1=E�e�=�1X9M�uB�NZ�1�g/��0�턅���>bm�TT�#�qS_���/��Z6R���kbJAਂ�:�f3+s�y���bH��{����r���:C*����>�.n+�s��K5⮹0�Zb���&󪐉�\�|hl���"��Fj����pl?�{@�C��aN�o��ͻ[C����qIh��*�gv�l��"3��(Ŏ�8�4�`��/�)�K?��^y��D+z��x�1q$��"�;�>b��|��7/C��HטC����i�dM)�/�g5ct�#��nꤔ1꽱!����u�����3@�C�%����w^����Ie�ЃQ~�`F��D]<�s	�����if������M��(t�E剀GZM�4���V��Y	5݇���@�O-A&�d��z淦5H���I�Z��X�Sq���;����4�y����$6Ӆ�r�� � ��HΝ����8g,@h�`M�_�Y.NV)0���Y����;�x!P�:��g۳<>�OH�[�5O�e?\��3?�,j�@l���N]�?�;d��l[S�b\���Ҁ�k�u�];&����_@הlN�(@
D+�R�������H]}:e��Q�ʷ�z�ߎ�c��2ޑԥ���Ε���0�==ǓH�U�Cf�w,�Bx��]��X��ْ�i)�[��\��閔F`sH�����u�l��	��d�S��c�i�rָ�@�;��xR��o��;3�iq���-�/.g<;(�d�{$���}�M�Ǖ��\� ;�����>��?�Mh���Z(�6>#z`��e!w`y��A2B�Q��r#�z1�|����\ݤ=��*�ł���ƚ��0y�-��n�cpoD8�+�5m�Ϝ^u�S���é_�J�KQǈ��(S��lu��̹F��ҿ�����Iӹ�*i{�.b��1c��8�O�P{��xc�Bz��BϚN�C���hg�5�G��� Y�ԝ��u��-���j_P��=&�؟,Y�Ì�_������Z�RZ$U�̋�勉�K��@�<晈��V𗁕���)u*h��]�b�蚄�=�	+��mR;nz!��jj��z��GR�2�H*#��@���f;%�^���rO;k���̍��|1~d�;
s�k���(���X�� ���d!оA6��1I`�
1��)�& ���� ⩐��l��֬����
>�wD2#�vl�#.���~������=7�#~:�
ںp�(|���^�?QT�C ���`��6J�W�$:����N�VrE�7��祗�l��,��@�հ�f&�8�BTz!"jE�n\-�/䚚�e����,{�����J�5Y]r(��E�5}��Up7P�, �&�1D	x��$�-�*�!�Z����h��Q�C��.�)�t���a��}�f���9R0�q);\�S�T#�ιA�c���	��	���.~�Ls��{�m�-�t^����&�雋\��'�{�ʪ̚��ͦ��IBK��ű候�fP_�~�츏�D�&�z:΋��,F��h�JKw�+�����IW֦��:B�����A��N����s�������1��i/�|0��w��]��&�����k9U��+��(���M��cg6V��k�`��6�V)�Dqg�t�c��*38r�ԇ �VȾ����&�%�(�x$�2srR��e�b��e����ؑћ���,�/)�x�/^�$d���i�iSc1P8<9�|cf��pz0�y����2�+��ď��!و�qv�V��3�����E����Z;�gI�!S����s��6QF��SZ"1Z7�'C��B"�#��9v���.b�\���%I����1d�L�39u�.��m��^4��;5�W�#�H;+Jm�i��T�]M��#�&���w�A���Y�[�:A��1�(��Q�.��6� |W9�e��f�&���;�<Dvh�n�Zh��3�g�࿙te ��G���o��J�d�'M�Z�2�F�Eg�����Ecd���5������:Nv�ʳ�"P�W��[�[���+Q~�^ʦ�L n(��KS\쓑�_j�Z����[�FN��s}C(�:�x.۬ugb�΋P,vWY�������/,��� �Td�����p��2���I�,˸g���y[���#j�)sWh�Ӭ 8��:;D��C�ʲe�y�Ss�:&�B���(D���QkT^ޝd�g�0�!�P��[l��2���TT�����