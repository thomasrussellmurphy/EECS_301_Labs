��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�i��a
Α1S%� �uj?�L�3��TLei-3^5]E�$��f�A��m����-uOɰ����3�nn.��Y:z�
ٖ��]so����(���5��]��[�H�8U~8�	��	7�&L%A��h�*cV#��ʋ`z>i8����j�-��=� $��f(��%��.ޛ�yU-��1q��0�Z���"^Җ���q��Z�(�Pׄ8ٯ��[��}l:���c��;R�ܯ+d�^�ga�r�R�?y>�oKƦK��d+�K�#D�1���$���UỊ":���TV'��l�E�	t0ޡ��SY&��Ge������K�!
�Zm��`�/��>u��*OE+�y�-�9��>]Z�ā���)p���duq�̒�	�`p ��kko��
�q`6���� `�n��[�R�PT�A��y�u�5�����A��c�a!�-GD�5!	Ϊt���Ebo��q�e���C�;�g���}�B�k4���ǔ`��`߰��?h,��h��b�r瀞��ƫy���4��n�o5�c^�x�e�Hm�6�}p;(;�� �	�z�_�����g�J*J�_\�-
#�VEwK�N~;
��K]$c�\����rꂤmf�P�r�A3�,�����kڳ��wty����Q�#TЀ�(�f���	@�-��P�X�&e��gθ�`�0���ҿ�*j�VUئ��v̢2�W.3��y�w��z�z�<�Έ
$��yX:�ʈ"���e����a� �B�H�B#�NyF ���^�q�{�:��d��y/�'�?����s^�Y�)fm�:�MȲ�^�ۑ�a������i��0�&O>>�{"jYG�1�\S�V�[�36�<�%`1��=���e�mp_��V�e�/��xu��M�E�D�ME��~m�K���J�oZ�����6�:,=9�`0�CF���h�εޗ(��X����E~S��f�0P�-ʕ���L6�AH`g�5q����z�Db̸��tf���ޑ8�>I!�-PI��5CR���%�5]����Ri ,�� B��]�J�e��H�%q�+�>��|������AG$�!�b�\Y��XF�J%܏�Z|�ɸ��Ҳ3r�g𢈴6�s*�<�����I�R8K�Ȧ�گ��S`i$�I�95�䴠��3wz�"W�8D.��<I0�<��aӇ��<����
n���X����v;�O3�/#����(?�+'��3�����z��ΪK�q��V�y�W�Zs��ѯVOӞd�(X��̤b���'N ��;������h�a�ϖ�3����P�"��/�h��?Q��yX�ڷ�$+y�`��R"6��'Rj�"�6� Af���4T�x'� ?��'�|�28O�L���N���6+.�=��5�3dp&�!a�؝X�`Ǡc�,�T̻��`9�
̘��5��m���/2���1���0Le�̲��X(����%��z��J]~��a%�%9蠁��?e�S��7���[�.�@
�k�2"
�f�J�ey�Y��� (ɋ��W�i!��{�[�����0��w��T>���N92�$�K@�ۊo�Bv����D'B�����Um��{{vؚ�����XQF�?H��� ݟ���͕"��oX���"u�_�[�\����C��w�M,9���!�L�d?��{���΋�$ �u�:t����|E�n`�
�PX����U�.|�gv�q�rʹ��=c~5����A˥}2�vǌ|�32/���Ĉ(h�5 �!* t|�;�m'a����K�$o{YIL�w�3�L�o�J�Rn�U"�?ji��@�.��5pP���-q�h�b���On����	X��DV+�[C�Rʮ��S{_���v��q�j���-5�f�{6�8!b�ߟ�f���ީ�b�[hJJ�3@u��]ϐ��������s��QR�׍(����Nsj�.�I9�l�3��ܔP]�!��k����
�]Swd��~̢�����;��R�z�B�O�1����' RFn���?� bw(�B�IDg~� ��f�hR�U�7|�~,<u�q�o�G��Y�T`;�B]]x�󴁼���X�6��2�Lz�
:̈́LqM�=�����!u�o���GT~�Y�:tC�.`��8v2ꇩ16��cbk�i�W�͆s8�K)�[��n�ߔ�I���{e�.��AF�c�z seJ�B�wn
�^μ7:�b�!�kD5�1���lև�ؖ���-3ɻ�j7(Ew�n��eH�<��*��%@!�k�K ���1n�\?Ⱦ�m�;C���8�M�`��E��8���2/�2���u�cG���$� �Dg�K}��D.��"���C��Qp[�h'pv�!��j��* ���h��^B8�Z�N��֯it =W�J�j���'��~L�_N+�$��^^eP����K������)i���w��ȕq�����x��g��Jc<emM4d�FM���Ig��b�r_(D�B����3�|(\�ʐĝ���7u��?���Jp�X�KX�j@�l��4����g�oç��`��.d�(���v�n0�{�Us��Ux��|��]��,|��;��j�@c�o�[�:����
�(7�8��^}|�5�l�bG�׫z��4h,6@�%i��L����ܿ��2R�!�"rI+���Ȕ�������_34R���<n��K��'!�sxUng�2$(�>�T՝}��@s�H'���*& o-�C4��O�+���#n]j�ra�뷮H���L�}�D����L�5NJGfC|��ߥs��SE76_Hv��5{�g�0 �=�'K4�?,�#��uN��gI� Jԛ���B� Ҩ�0g�6����0��kJ5�T�'ozO�б�6�L�?���.�9�W��u�l_a�#�Cw��qZ/T>S���κW����g柸���"�GvF�/�O{;�їg�2'�-<�c�R�H�N�NN����.���Vr��J�t.y��Jr�$�b,�[ρ5�H
MA;��q-}{yLV#�n��o{Řju֒��ثj�Y/Ծ���M��ߎ�-�s+W`	�����\PWb��e�|�>�>, Lꍀ�����	��Ʃ� >���ިF	RPd�2����u���N#呅Y��◺�<ֹޣ B�d�����N���=�źB����W��Tf>ν<����څw5r��T�Jj��L�R\h���N>V]��T��j��������H�A�Jk�?�}`��4/���aF$�]T�蓯��PW���ph)������gz�����*��Nwd۠���}=]LN[{�&�4`��a*Lp�XO$�`1���f�fTj��ps{g����}A���.&z�n�{J�/��r��.�;y,'].�����0���X1Nr��~����%�I�/Bf~�M��s5{��uA��L��v�=��8Q�dJ󘑝��7�c��jEt�����.�+�G�)��|x>2ZP�g�R��R�����כ�VR	iHG^h�15�E��~���uX�w�9�~)�*2D�c�Z$���j�:�5���Sx��L7�z�&2r#y:��8}�$E�������ӫ/G�D��x@Ic�bU�����v��Gg����2�G�gM�4�Tқ<��])��f�A%m�ZG�B��� �<�g�!�I4qr�����dJmٱ����^l����*���؉i-o�f��c~�֛�I������y\�7�#G���k�0���'�U����dW$�J4"�i�{jK��	�p�Ȓ`[���1�Ñݑ<F)�x�=v8��'�5���V�x-����3���|�*�Ƚ����}�߽m�᫗reu����������0Ǔ}�z�!�s6����2�i�s'�>9T �n��
��7w� ��HfiQ�E�V`�6�ZE�j�3�xBI��t�aH��N(v��{6��Bav6t��y�=�1}\ ,;c��^D�Fԃ�7�IG*N����ɍ�w��)�q\3x�8R"����X��7�vHtT�cu���g*��#oq~�?w+
����>�t�`o�B�!��\�����f����n\<g1�%��~pћ�SɂO�O�rxGl���\4�C7�2����C>6�4f�Xrm��l���b�O�p��rx�s�R�;_/�J�|�Z�zg�c��˻�oy�x|,���d{>�u��S�;MV��z���xK��2X��l���[�h��R�]��,N��zQ*s�,b�3.�kfq嚡��[/^�����NW�0yë��OJ����x��ڍq�����ڥ�:U��He*!�	�T�*�ߊT�����*t
�'zsZϢQ��e��7��0�E�(tjޒ䓬��8�5ѓ� p	;��	���ۼ�x�8�9������˃��,�P�	F���� 5M]���3�Q���hyӢ�?l\�F	�x��Z÷,���kl3�	Ɋ
*N���F+W���W�����{��ge��W>Rd��:R[i�y����X���Y�̟�^=�b��>��b�}V�m"�W�I�MJ�x�`Ѻ�F��#5`(޲GN��4SF�_X��O�ج�JKu���?x>�jO�'�&08�d7�we]�3L�9v�����Fb��FJ�1�?�{��Y2z�w��B�qU1_�_�՜��N^��yb�`��C�����!�i3�j\D}�].�b"6C����g��Y� ���4�HS�k�$�)��e��̓a{�rX8�&r ��*��c栕}7�H@m�L�iFn[�����O����:X݇�G��}Qi}w!��h��v7<�zz��$&�%Oڏ�+�ew��1&&���$j�͐�2��?��r��<�o����i$<P<��չ_�^6��K@[U��������W뮴BƐ��؅�51��H��j�F���zJ���1ﳽ��ڨ�m�9HB����K��v������yf�I0=v,;�I�5��ݿϐzל�Bkh��g}4�8y���J��'��G�B><����x��1�sj���H�E{��x���� *t���d:��j�/�{eD�s!��7�qĵ�	L��GzY�n�"=n�G�@|O�k�k�k�` �sV;޿��U��`,7|���q�Z�(�C��m���/LRR����]y�J)_����=XƝ\ǿ���h�Ÿ�.4+l�E��Q+]��?�����!�e��5_t'[䥈�Ի~	&��+X�Ah*g?��^9C�>ja�lu���R�_�-�n؞���<�`��ho+m�8� �P������R���D���
<v=w5]���j��9i]��%6����k�f��G H��@U���J�L�ը֞Q�\�#��~1��4�C����n��!ΠPmng�"��A�ɫ�cu����e�;�n}[�Z
�"���Y�g�~�B���2�)��ɉI^'����3j����3ٗI��%/�k��R��y?I9ff��'�l�r�zN����J�{W����g���A��Tl�-~��Ry�\��=���a {O�F���g<W������������=���i-��ow��!`mz�&�z�������!��ְL��:_��)�U	J����(P�:��PYC	�mxR��5w�($쒗~�vt+��$���]w�*.+Tq��i���"�j�[���a�f��U1���i�R�?�����Mޔ�y�C>�o��+�E����?C�[%����xCq< �U��سR4L ��A#ԑ�:�!Vn ��{�6���c�k.�x.��o����F��Fe�ʬs��Ťa�:zY�>!:��ʣ���� M�Z�x�U��X	��Z!�O��ag���aU��'gNCy̬o���<��E| �2�Y�[L�~�g������4@�;-+��/�غ"���>(�_�{G��� 
1�!�굱+�ۺ$�H2����d=�����6�5%����3�w�U�m�
r�t��ֳ/���m>�$Ư��oB�V��{�m�NAi=�^�� <��.g�u_Z�$t�_D�-ǧ2��D<I�h	�Xy���,ߞ�`)̚W݇xa6-Z�u� #�6�d��f;���T�4���2��Z�s�Cgd�(���~\n�	�\�iO�l����Pnn|�L�,�z�%�|p�=W6�s��6��Kcz���1 �$Q��WԼ\�\���Z	2Nȹ�?E�Y�4���L�뇔��؎���� Y#�A��Q[ߕ����Pu�F(;;���Y8WA�j�".L��V!p�>k�˴]�����)U\�G��
U�T4�4���T��J�I��;�ՎFY�␴af�\�u84W�+t���� �����/¥�%G �
�)ύ�dm�$�n�@з�ޔp�k�v�^~C���(�Au��W������g�N�"@Cғ�4jRT7��cx	�� �F�5 ��r�&r�P<��b�.}���P����=i;��d�T�M2��~�����mP|2��HN�G�"�T9~�M&�IY<ľD19� �R�2	B�b��ܞ�8i��ϝ�*N2�X�߀�;@�%(6�l�^J���sa M�`�=#}�Nk[D'�)Z����-�~I��40���Lht��*2V���Z٠nj�ʹi�8����< v�=�ͳ���Ab��٤\��s�l\{S�u�6���^
�C�h�9Uդ��{�w�T��1ؑ�L�D�Ϯ��X%9%O2�ÕN��eG�����.��Dw��-w�[��Z�F��؃!钾NVX��(\��J9��gW�HLT吨�
Y�8�џ�e�A�4�x�[�2t�9�L�{�ct �±W_�Ѳ���0G��E@ �;"�|���2F��:�hf����|<]͋�+��A0AǊ�ǳ�a?�{��xῡ�؁v{���>��N�)��.�h�~�w'f�z�~�ѐ�o��۸;��1�;��]p�$�e\�ӕ$jM�(s��Bs��>;�Aum��E�=����Q^LӀ��C�v����Σ6��8��>��?�Ll|~�e$�z��]?�s�m,pTN*@�j§8L# ��!B,�T��79��sj�9��
W7������n"l����UZ��k �\����^�x���X�_�|6گ�M���N7�l���5�+���n2�u?j� _y�:!5ST���m4p��V�qj��ԦO�*:]�=��SuD�ר[̵�!\%���en(����7��T�x*}��/�5����W��^��o%�~K�.�z�͡�W�T�M�;���⚲h`qߡ˅�׺P1����i�K��X�g�x� M���hJ�6z#;G�H݁�攠�:e�#�	J�A9vG�H���
M�Ju�U�3��NpOZ�-6��G���E9���X�b]r������
�i
�+U睋oH�t�m�in����(�(�q1�sY*=>���9F�f(���[`*�0y�\N�1�QN���Yߖ�L�?4'h���_�6�6G���Ԫ�g_�L#�\���X���}�V�3Ä�X�A@1pn����~L������$�ȫ�?��=rG��#e�P#ӓS�T̫@9�V��~?��""�d��هq�,4����0����f|=�(Ïw8��t:?jL��kyL���o�B���#D�S}��֖�e	�UݫG�ye"�I�J�\�*>w�1c�?��X���'Lg�Oi�1��	���JQ����d��u��+�������DZ�͔�^�����-#Y�+ �N$'���{(�i@�j�;�g�$7�a|7hH��!D�X!�`�t� �zv������.X�jZ���~�
w�XO/���ß�4x{���	 �!3./�!$�0�׃02R4/��/�(�-��\t��3[�;�:��_�fk�Ȇ���#�i6��ˀ(r(!�{0Y�y��F��.�������/�X,R���>�m]�W� u?�a#ڗ���ּ�y~�ZR&�J�[�jsC�V��@Z��A�/��J���|s�V��b,�9�2,�%��������<l��r��)n��^��T���H%�[h�z�1�h}���p�N��7��BOb�y��(ݚ���I�0O�p�<lŬE�`LVa�UmX~Qeq�� Y~گ]�n'�"��o��8�M�9o!�BGh\LKy�� ����p����c v9y�>k�,�q�~�ݜ!F���� �':,r4�R�h�4��D�?,��������k{[R��A|��b
xcҷ�}��N�
�#����cQ��E�	� k���}�5�LN>�� D��zX��44��� '�'?o+j��"���U!�B]`X>u����{{P�����L�|%����)�����6��g]� ����`y׌�"��ӛ��=Ż*�@�P�cP���j�o�|���ѿ}E؎7
D�B����j��kH�}�vwN%a�pbr3�ɘH�9d'-i^tЀ�=��?��cAn7|`�k�I�>�2d� �}�![���t���F���r|gh��@�N��!�Df���X�a��RuR�<��ޔ�/�5�c�g���&/X��c�K����R"ł�N$�|�PnJ��,����z1:���=V:�d�q, ����8�1`