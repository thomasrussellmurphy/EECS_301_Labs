��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv �|�
����)���R0j��3I[���Q*������[�X��D"ԏ6d��{�0I���}@�J��1�^������W�Ex�i���)w�kN�n^����o1�B�1�����|��ȕ��,�3�[OU��F�- �[�� �o!������*�?>��i��3������#�P}k�1���ٻ��>\�t�Ʋ:&���/��C�o�%�q:��o��G��$Q�m��8�r��,����E��@�I�V�k���A�.�T��Tv�)�~�a��y�I��5�#�tK��=�Y:}��2�t�:H�Q��(�Z:����Γ��2mË�Ӎ�T{�/n��3Ң��o�2=�7�����w���`�����pcWSK��lfI7 �A�֠(���į�$n<�F���JT�������O�l���>�|��d�v�wo��_7
eSI{3Ch�M?6�1k�{Z��u����W��S��&A��(�ba��h���	��ߎ��(��V]�Vk�E��)��.�X���-!H=���9�F�V�9w�i�P?r����zȐ,e��+����)�qh��ܪ��4�[/J2t�WM�B
6�A��{��QU�Ŵ����~5M^%��w�$���2��9h��?��p���Vy3An�#�lK��z�e��xz�x�b&kM�2�����-�]��	V��v�,i�W�%�ƾ�&ϬcR���WK�X�|�B�;�e�3�$Tj^V�y�u��!�q3y��V�.�����vM��T@P���3sJͷmb�"-�Go�#7�]Q��~<��x2��9
�x6��G������Z)�����/�5�M���!�����u	u��@�Ą����&�Ă�	��7)��g�o�bu�k��m������S��i ]�_H!�ս�]�:V�gc��n�?�`�;��1�>/8g_����-K�>J�[<Ք��DIÁF�S66�Z�}�B?�O�%|��0�F��b�h��4���g�B�@~���[Q4��쥄T�x�רʹD�=�Q_fB��QE������,�^蓖�ƾ3Mb�H2�����Y�9�5���5l<0Nh�� Y��;���6ɮ���c�%�4��84+�:b���Rdg��}�oڙ�iy?hc��1���o�T�� ��Xma]0�b=yo˔6�y;#����b)��O.W[��b�"�h{������YJ��(����骓�d�����C��>���Yڌ���d�w�v㹝2�tr}q#�f�-��Vpy��Ǝ �I��/�U�QO}��z��YW�JD��N���
��p?ʔ��ސv�n���'�"��H����:����h�h������+[Y2�����,���g@*MsR7���l����i���}7Χq	0�v�W����0����
��E=��.��v F��V�R�T�7Qmp�R"�UPOr�)��3"�'�}�!�z��Q�q� o枷f��a�������̵J�����Ѹ3IGՒ�1����1��Qm��9~k+�3I�i^� M�f{醛��*_dw�-|�~��H���i�����8	�%�<o2�ܿ,��4�=!�
8�T�����+��^tRQ@������0�H���l�s^���M�r�Ve��27�wu8�[���>���[�$i�)Cs�9;�#�ρ[�����짙� b���l���Dsס!T�DM1�(�#��cy��7u�ٗ����4��'�7j�b���p�[���4q��s�����Bk<��-���T'S�i7KR��	�������ӃV�T��NF��j~�iא���ꑴ}��f��g���-�L%�7l�Jpۅ�s��\U�󇲣�� ����H�Y�U�߶X��6��*�' ,� �U$���i�C�t�xN�+/������O� ����}��=���Q|" <��	_d�E�INs#V��쎊XS�٧�U<���П��1,;t���Q99g�<6D��e�=�l�́��; H�wQ��EZ��G����T�oh�5W�.U�v����Fx���(#e��^0�@�f�u*{W�ֺ�i�2��������1<�v�G���<*���,�a�x�?->I$�����!@�Kqd�M�=pVr��b8�mS��X\>�Z�X�t?.fE����m�ʺh$���U6�ky3=i b5W�dp�]�H԰���k�I|e�t�e�B����uU�L:���]���/�����+��v۲�����5�:J��6�p�=��4��iV�+�Ve� ��{�����)���HC��D#c��O�洁T�\���hA�{7+|��s�@�VL�T|����UFH��5z	�舙��7u���\Hۏ8�Q�92���X�`t�k��n�X����&���	�o�l����U��P��ӵ�0s̀sa}����E�`�in�2W+*��笈�廫&�-��x�������z
<y���|��}��?�Q�`�ĥ�@��{/�M��ǈ{�E��iK��[Od���?<�f��{��u������oy +�F��"9Yd��(!��
���c�c6���q>yS��Q,|@T�~��p���-�X�g����:1ݢe�R���B�����RG���_�|Z�nIsj]������ݵ]+��jFG�R%ɮ��L;��PyHŠ�}���͓�mF��4UM7�gV7�*���qi�n3^�/M!�v"� ��a�I"=m�QJ��וa �w'��qѵ^V��T�lKG�g0������	������ҒRC��T����2OȕO��0Gti�v��-��R�=��V�aT^t�+��P���r�hiH���[�b+'�j��3q�s��p�
�__���6�<���ڦ�1资`�b��*|GA�q�c�d����͜������HfT^����SB����{b�ǫB�i�#މ�%��V4*~s�`�H`��:O��R?�[�|�]�$�?�-�2H�!����A�qq�K�U����>虭��q��΅�݄u���S
o�v�G��WKYC>�G���A��L:�v>,�4�����p!�G:�Aa8_��~�Hl�wN#���^��3�DW�[z��l���^Fɦfǯ
Q	�)�B|	F��Ւ6�&te�Ԋ&^26�1Nt��Ǭ"��6��/(�9m.�&�?�rJ�!f���b�˦��$�ʬ����Ƿ�B��"���+8HI�l���ѡ�뢲a���E��4R��w,�zRx,��˖c��F���꒥�]Q�\㰅����&]l�\�=Fn�\gϻS5��.2�_��Eͥ���"�Ya��=ema/'%9��oW������X��&��0�έ��5٬�D	���5R��5�D�x�6 Q�XO�� �<�~�I���0��;�E�PY,��C	�65�nQp��� ̠�ͬ��t7�	 d�&�_л���r���R��E��Y���ͺ�?���5`��{EC&obi��$��%Ձjk;�zp�X��_0�Mn9�C��X�������V��2�1P�ؕ�9�5�>�:���� �H�G"�w0�)���Ι���'�ɠ�@�;ki�c�/�S���1�s�ӡW�rkY�M0-����M���^/�#�IV�p��3���}�9(ي/4�In���N~:����̯M���차��!���1�C8栦�֢���䋁��(�-/��t�����N3�5Z���0�_�T�=0�CʍBk .�```Bܾd�4�=-��|z�>��+���ʂr�Hيt�������"�G�+u;�b�9d����y3j����2q���q����N^)g{z;�<pJ��;�@m���ҹ�(D��`�]ہ��KL��r;O�����}���r����������f����H�v��>Rj�CO�*"lr��!�H�v�n�(GW�L�k6�["�!��G���G�:�#/��G4h�����������[�K�&��p�_u�o\ڂ�v��I4Zg%�읾���5
DRX��Y�� fx�~��g3�!\�_L柉���=��.�L"=�%�chޘ�i.�u�мMM��r��$��&��us��J��}Ɗm@��1H�W����ާM�%WV��.��Ǹ�c�y��S�D�����s�ZP�دƃE�r�G�F]��Op "Å��Pۅ7��l>����e^L0����ΙŗBk�x��A�j�%.9�n"��p�,��$�S>�"t��D=X!\2N0����3�Gܢ��U�����'Nɔ&�FA오�ǒ'X#����
��@�(�'(4�w*�=σ�v%=������ΐ��(E�����V�R+��0x[����Y²s���D��_�M�*�ql��N�t���������X"9%�'��ȡMKK;
�HG�7R�T���
�q����/�ԛ -Np�����<��u����KS���
���l6K�_I���s��D ��'�ǿ��"�uaknx���~ߪ�aa�_�tn��1@i-�Ãm『�SP 4l7�W?��t��=A�u9l�P�*�ּ�f���{o�;<Q�_��w9�U�����L
�'afJvS���n;��		���Őў�f��-	<�* b-�����Z�j=Qr�"����4|����Vpu�ɚ��'�j��_-b������'W[�S$�@S�\�P�pa[X��Rȟ���A��#)�S�`��- �GѾ�E���DO,����MlC�s}�R�%0�1j숓"�����~�����e���.�m�� �@6��-��
�`���H�.�$�q�c�7�918ߌ�R��/�5]�dT�]M�;���m�R��PY)�O,P\i��}G�Ͻ9��:2ޞFh�y�{MS
K��{o-�^���@B����P*cd�����GjVNnU<�zU �he� �z)�p>�>) �?��_�|*�� ��\�0�w������A�-~���Qig��9|�?�=!J��X\1��Vȗ|Tf� l&/x^%�m�Y�X��; �ʻ�.pя��zE�1�C�:��P��w�,��ei+bgp���Y���e�h]�v!��cb9й�.X�g��rP�AkZ_s��Ӏ�^���9�&�xR?&[�ɫO4;�3����c!5���k{$Ȇ�\�W	�^��P���_.#�Ň&/�����n�4Ƅ:|=������Fχ�F/`ee|�F)`�^��'b�G�NN�gËH��Lp�V�m���7kH{ig�aa�OԀW�|v��O�'�7{�k�q�<<lxl�sE}Ϳ��,r�^ߞ��;����M�#�|��?tTr��D*��%�3=���k��T����_˪N#Z;�(0̆ʷ�%��'���{��8�'taͦ��1=�i�UD����y�m���&T�Q
�ӣ���m,���,Z���e�����F��?K��/ !�6ja{W��~�
f�E��K���7����2a��p�T�`�Ŵ7��I�"p1�t������eC���}��X$��Ļm���,I�
&rCb��^�����ľ�nm�F�H2,;�I���]v�� ���;=�����E e��?/�pt�PrL�s/��éu$��yXq��'cQAb��t�4�R�=��
���w�FNO�t���Uk?)Z�QX�<�>�X@��%��[3�g/�S����j�u����Q�Q_�E�>u�1�@4�;����{�Y���SR��l��+�$�=%�1�@���^U�vcK���5��`>���h�jlZ�'.�VԑC�#Jc���3�����A�A���A�R��s�����n�U�"�U"��W��o1i���W%u��i&G�AT���2��Q�Y��}"t��W�f�����p�K��_8���uy��!�<���ɩ�य़��J���S�����t���9EWQd�l�\Iug�c�'��$;;c��1 $7� ��l�~A�a@pEM �N[���Jʋ�݅�AD����Y�f�I���ɘ���-F�dJ̳W��آ.���q����}
G��1���/�99��0szr�~�OB8C���I��}O�
dC�7n2w�}�a�}������
�\Pj~�,���4 �jW�S�.}�>��T�@ݠPs�܍�R�w�{tMY��FЩ(t��*��z.(&L�Y�&��#�^{f��h�֤)	`��͠�;��%�- )��\�����0o�-�1èR��d��U��:�=�&%�a*;�C]�)��a�$�3�'ŗ>��i����~�ό�V$F��|I��J��y������}� g'�	�f��PL^E�o�����+��QA���*��[��O/�	���y�x�>��y�vl��-�X��w�F����
ݕ���������b	�~�q^��ܚY^�Z7^9����.TSߘ2��S%h�{����3S,���`ǩ��: ˗��yGb�>��&��q�$ȍ��L�L��;6l-R�J�{����~�Q(Ĩu�?�yN�m�V�f��ҡKaS"�7`��f��3�B�+�&3���{8�-,uUPq�<��52�Gh�S�d�pF��1id�r�������E�m� ���$pڧ��$��CN�Ak(�}����aC�>!�j�G��?к��֕�z�l�U�M!��u�����MW�<��e*�I��`, �s��i��L
`'�@y a��	"$�9��d�J�.�b�0��Vw��y�hs]XD_�=y�6Z����W�Yn��'�v�*�<�F��|����K1X5�'͟�ܖ�=-��h!����L�����c�@Q���b��Z�-����'?��BS��\��T�W,zar$��������s߆.��q9Y%�V� ���ֿ5�'Z}�~�`�Q�Z�n��㉕�Vw��n�6#p	���P��3�7z,r��L�B�~D�n�i�û��rT �E?��t���� ĔD��^уj�����'(�ոS��T���t�Ŕ���Tn-p>�.��ҡ9	ԟ�� �;?ǝ�C]�m؁� A9EN��?�| '�@�i�J��K�$4���*b��e�y���{�x�p���Ǖ��
�|>c�O�	Y.��1�}/��4�Fu�U3M0\���֞j��cL�W\�܁�|����[Gko#	;<*��,�)[&��GՅu<^!�>�L�)IS!�����z�]��NLǏ���W�'�s$P=jaA2�E�uYx��Cc�p}I�E􊝈�wk#*C�o|b~E�ˎ��V�ν���\8m�]���������bc�OM 1����E���	���lgR�֞@�5ށƖ �@�cs�a=�k��$Z����k�C��c �K�~?t2�:V�C��+ Ġ��"�PX�����Ĵ�@��Qߤ�Fi*'��"��.��ьe�:�!����r+���a�T������0IW "��N������@��QԜ�h��l�C��
���6CB�����շGڻ���ѹHk�"YU-}o�hN�u@"��0)��7���Y��B]�VM��:S�0�#r��9|���>�S��=UT�����i+"���d2�>��Z���c�[�Qgb�L�G��{���/~�m���������DU�W"-4�ɮ�#��:��J��W0VJ~v�����4���:AC�R����������d�Qs»L�_�+����C�rq@%Aӹv$����B|3c�OׂY#��3)y�S����"2f�O��V?q�>=n�W���4)���.�/���+����8 |܈�HC�px�d6-6tN#�Ω^��N���Ϟ�@��[���*���t|�#m�ာ�L�8���3�seNV<� #'~�^ص�l�䂐MM�4�g�I�2A)�ef����{�&`��R��I��%�"� �V]�G䁈��)��]!�����{�L���Դ!<?���c'���Dvo���;I��@�N�"���=!���p��U`'��SQ�E�:.8��y�G5j
�t���Y�v�r�1�{�% �[ő�L����ͿR���`ܩ�&�����B����W�9�aE|:L5;����u���S���9��o1���b1���3�f&�jcŨo���N�VU�����L�9�(�/��:@VD�Wm;�����w�M~ུt3�����q�6E�̥8?4�䇽�T�V|+c,��n���mͭ_��ss�\��$�Kz�r�o��J�/�HI��,/4	�7`)�Ðw�a%���{l�k$���;c�Q|tq�Λ�y����G��xp_���x��9��w߳C�￸}�O�#�O���mٺ�O��ҋi\SյD��u~�xNs���y2�}�].��y;:��obH4e�"��2�
P�Jڷ�^�&�3��y�: ת�ᅻ����j6Y��f�7=��'�\܄���X��o����z�qkB�58;�h]����EI��9�n$���R���ɯ�s,����LYV ޲���;�E��\&��_��@83����g$�`*�6f���P�.�-/��a��v#����"�& ���[pT�N��MLl��w����o��l��*0�H��l{��^��|y��\0ڟ�;��(�3$
O4�-���ț��ѥW	_B�	��2UD�u�p�R_�u9�
�w���E*=H�{�7.�mb�0����ķ�����#���q`[��篤w"�s�;�S�w�l"A��XM�]�����y� ���s渵�����K��I���4I5��֦�f�UY��p�g'� q�o��k��7��y���E#�t��I���c,�~J6$���um%C�Y�pc�u�h��b��S}K�}MkZ�곥l���ɷ[	�Cm8i��FC��'䀏����0�쏁x3�F���n�c��k���nm?� �����2W�s*��:�dR1_��U�Ȝ)	��6��r4F}�j�S�.��#R�?�91��z�N���ق^�y`���_�����{�g��Q7�\����@F�`PX�Ȃ}4I�E��ω>/�ŗa$�c�g�,I�e-�ޙ��w�|�Y8�Hnڛ�3F���R��њ�2�⫪��Ż��mPuˬ9?�$�.)��.W�_��#�9�֕������n�>�QCO3܏�p�YL��v�B����>ÎKf|hɋ��C/���;��j�*0�x��O��坄�^�wNjYǏ�R8-��ѧ�$���$������Td\��<�Ѱt4"՞�G�>�܅��0r��4���VeN]�a� �(���$1,�i$RԆIN��>RO!j���5�Dj������Km����cjY�ق������wl�i񮁝j��&�������#�|�t�3�>�_%�̶)���{Ug~�C�2�3���㈌�>��%�)�Lg�"����1���a���?��L��o%O�~<%º��'��@�ڋp�"1/Bכ����wλ��k�8+�$��cID`���% o�\ۛ�)�rA�C{d3��r�A�k�@y(B��
��Qg �B^ӌ��f���e�q�!!�g�ݍ�V��d���]��A��?��`��� r?}!��^�O��֗�~0�[j��r�86;|��ȭ�=	���E\3bI������x�33���k�t1����w@}>�
)�|K	�HҒ�O�~�p$`���!�uaFk$�2&�>��Ӟl��8���޽�W3?D&kמ���(�C��שj~�VID���G��^�G�@Z�`jXf��7�����Z:��C�pUk�����U6�)�]y��Q�aD��ُ%�§�
�--j��H�UY����hg�_��a�@rq2�~*(ң�>�����$U��U�$֦�~�A���P�竮��/�~�~����=��e�ȣ�;8�{�i|Ɗ�j~F��˰��-et���ZT��9�oEhW���ʐ��i2�,����xL�y��FT+�?� �_r�m�@���u���h+Swpo;Â춱�H�]NM#�o8�'A�Q_�'���f����e���)V�s~S�)uI��u��j��4*��'�v��)zܒ�G��KJ����̒s�|�l���Kj��g�|����1���</	����K�;Qg@����I�)V��F#����,��+I}�:�I ��0g�����/#�;�*}t����K�Ƚ50ـ��5u���[
�fU���RK��C�P���oL���T�:�|@�`�ev�@�*�˝${Em筮�v�t��W"���	a���j�᠉�[�#�L�8:�
R�
�@���g�;����2C^��Gɹ6�"bjĥX}D̴�����n�#%lX�7���B�%u�>�ӷ��0�HBJ�pd �I��i�����ֹ�������]y��-�)�S����U�v#��Ȣ���{/�' Y+d�s�GS�SuҘ��Ŕi +}�/yR5H����!������'<v����j�J�_��t%ą��諶�n3�x�~�q;f��W"�I���}���M�Z��rZ���%$B䑜���2��g���3����M��a���EK���!T�������Pe_���Ck2R'4���윦�Rt��vѳ�kH!qI6T��Y�{S����7!�Ձ����������bR�sr�����T��oԚ����8wi�ۀY�cК���c�m�ijc�n��8���l�}}�(�@�<9�xn#������L����
&�k-�s�K��Ց�����]���_�eP2��V���}���`Z]To��P+~�֫Z�Q?�HJ��*.��
�D�w�PF8i����?Gf��<�XӍ���9�����x'�U0q�Ί�[�s`���Ѹ�N\m[���Т<��Y+���w�T�E뿀�~>�,ع�W�%���ǧ�z\���E�MNb��+�TQ}߮<��b��.��� ;����d��k^"X���/�+��p�l���,�cD�k�Ԋ��S>���jJ�I�"^m���>.):�M����+�M�wMX���4�F�;������V�h�B��{lDF�t��~Q���YU�L���s*ޔ��<���C�)E�ѢĬ�h�f�y��{y�7*>���g��v��s�O˽�ك���g�v+��HuY�9���$�M���(3����gce 'Ả��4�j����c��s+�1̃0[���q�I@mYi���ؚ�TP5���E�x' ���73_ۄ�D4D�zP�vGπ����x�:���c#�|���l?&��찃]��ᩤy��u�"�N��!��ÑO�W�����E��`t~�6�����]&.�)�D��(��BF0�ۇ�/��2i¼vq����$��c"��Lě��(���$�(���-�OBoX���{�"�\�,�g�� m�_f��;�a�˓>W:�ATm��_�8�!�{z1�6ߦn2&M��0����<ފ��Q]���I�1�[�@���<HG��^}L�K2-A��4t�꿥�OpP0�FW� h����f�[���<��ZUlԩջ�/�b�X%]�T�%��Sބ��U{pB����T�i��*M��B����Ӕ[�㒒q�V �G��"]�Е��k���Չ;',w���8���8)cZz�M$r���a�S��Mk�� x6�������Q�W�Ÿ���ܻ��>�����.jº(��ZtV'O�� 0�;������T�g���(�̓���Е�������)aH�Q�Z�m��ۍr�9�)�[�:�m2���!a7�����Z����j���~GC��}\����'U�����u�G*���\��-s���L����Y��W�ó�!�	�#��2��~�Jp��W�C-�\�ePƹr��.s�X��NP$Z:؟��5��$���݊���GM�#X��0�����m������f+y���T0�?���)9�dަz@��/���y���$��ў��4����,2�b�sM?�MUO�R9�1[�%B���3��G���k���V�g��w�*�ߊ���;�hJ2���	�5�L�E�ň����@��X˺����`~��)Q�������Q7fP#�|mx�ߝż��%s0!_�c����>����dk��j_kNp���{���G�v�)���d��i��v�z�������E�bv(4��c�X����z:��i�V�D�ka����¾�s�=�>��{%|?�.� L �{A�~�pD�����%>�2ϣHhJ&�/B7���F��s�����\Nm�&�>_����ݙ��`�>-JV�K��-�`b�W�4|��B��)2F��j��n0zC�����51�4�Fì�����8z<��߈�S�����.Fm��3�Mg�VD/�������?82�KY����N�-b��{Бc��@���v7*�Xb�I�Yw��T�¬��P�u�� �b����
����Z�xҝꚢ�d��j�d��%���/8�L־C£�o�@&�K���145�$�?���H��j	���	��e���F��E�OG�����0?���g2��PW��O����cO������|D$ne4?�\�Sh�����?,B)ӑ��1�:<���&Nm���`G/?Cruc2��ams/y���s+C��1�1}G�������K�>Z�C�~=e���i�>�8{�{�s��K*���;�	��۫k�w��gS���_�����΀��N�N���oC�e�7�����\b����~N����ne�C|�R8��V-HS�*�e���F�'���l��S����P��%�ɮq	��@j�s�Κ�<��Ո�~	�9��kzO�U0斲��zܐ�}2_�qv��T�E+�����R�p��s�C_�A�k��;�J�x�0`�BV��pԬ�w���JP�@M�K��l��r9�nR��ܺ�uT���3���D����a���u��܋�4��nh/Ⱦ)���c���s(�G�I��珰�ɒ����$(�In�#K%2�K_TZ�g����N"�U���!�4���a��WE�?Ξ�c���6�$pg��LqA���+߅mn֔�=�VB��;�r�{���@�y�j����� ؂v�b˪��%�0!��m���BM"�\YQ���p�@�I�Z-�^9q�u�}��'��N_�&�~#�9\p��D��4�?ޏ<�E>QNg=<����޴�ئm�B� �3̬R'T)y�^�$��M)ڠ��m'Us���]ZD�࠸D��n@XA�������;:�ԯ�
�M�Av�	�WA���~��,�ԅ�nҝa~9x���2�*لid�o���&��)�mڅ�#j�K����e�W�9������
d��n((&3���
�
9���m�
A����RJ�e��k̎<yٸT(u�cD4��i	2N,���5:�U�ߕe���K�w@b�0�T���g��xt�QCX�  ��.��6�w�ԓ�����[�6�u��!8v�i��po�~�Y|v��yXo�c�!?�~�j��=�''
��~(��N��*�����ˁ�o^#k��|�7�|��J���y
�5ΠM|!��D��0��
�$���X�$_՜�4K�����JRS��ZF�?.`������X7�Ձ�%J� !�m�.��#>�J�<-��>h�r]��!S4��o�\�%9�s�k$o�0�	�m�9��p���WW�&�o��P#����\�̋x�kq4��S��9s�K�Tɍ��@v`��2L�|G����(�����X�Xߓt��80�DO�U�J�7�5Y��9�����X�V�p�Q4��胏釱�uXY�f�S��=t²������;U���l��Fڟ>L��ܝ7���3�f�������[p���^��IbA���x�.���Xg~�����h���?NxN�/�[Q������ޅ����]Tn{C�͎���q�t5s�6G6�jya�X�ۉ�����o`l�^���8�07�t �ٛ�e�b�.�r4We9�i
�R���Sy7I|������O;�'�U�O@��%���+�j�%˫������_��)�=om�G;]/#0�)4%�T�_����.gg�^�,ѓ��I�̠���A6OG�_-�^�G�p������Ȉ��L�L���X�2�i�FFN���E\w�m\4I�^�Z�ъef+��z�(��	;�s�Tj,2�1$�(�	/���>&�Do9�i ��e�)l�&.�:۾Ӛzf?��t2�fLr���-EXT�a	�!v�$��L:ŷ��"������oh��S�+��WaڪNb9��FS�҃��ფ�u�o����Fs;Kx�h����)�:��d$u^3WĘ��9�j���>CdT��q;����0A��a���g���x��:/Msd�k!W�u�,�0E(��H�6yů�!��o�.I���ӳ)G��{�*�~<ܤ(�9�G�b*,ն����)n8���WT����(������(
E�O_z�W(���5�Û�
���M��j��{�$�?R��ᏝC���;J�!������6�'ꠙA�UAӗ�f՗�N��+�E5Bu�aoN�kn����DBba �Ja��Ձ��c/�ަ{�� ��2���(>��[��P|'��z�g<���(�戳s�����<�9Q��,TtJ�dh~�Ɗ��J��i-L����G�ZW��{����.$��� iȠ��v��eX�t{�}��6��K3*�jp�!�
K�����7 �5���c��P|��8<�U��~"@[u�$jP�9m��V�Q���◃��W	�22� �#�L�Uq=r���PV��_��y�B����W|ԧ7RIl7���LA�T<��1A��P���RV�n�rF��Ȣ]й�=$In��k�'��7�`�ܹ>���{�J(uM��rɀ����7P���rO�	}-�楴E����6^☼|K�K��K�6:FC,��C2֎�o3�{L�ᯰo�5p�xyo�i�i	7g��ݾ�KpO��r<�#[=�G�Pa[fv;h]d�0'��d�W����əz"���jw���+�gSj��87>_��Ѡ*FuN���d�F�UBT��.b?��A� Ú/]&zK�ph���1�<�L�'Z@�#M�#`-�Gd�Ɏ3�ӗ��q4�S��>@(T�!��q��>��0Vo~�w�➽Yj�i��R���<��pMy��jIm�V�x�v��V�wu�A���qW�24�X�p����"�G���{�K%q�8�f�����D�>~�H��������#�:�;}���O^h�R���S�hp��g�cDCE�=e�pP)�:wA#NZ�����<4��\�JT�.E��?���ny�q~��?�n��C)�
���C��?9V~rp�'Y�I� �'%��p��lu�:�^=?��r92!a�a�ۇ���Q�]��JL`�
�3�p΁�0�X&�N���k�J�(3��p}z0̤�`�o$�m��1|�U��N��3���H&!�&�,mAc��_� �5�5��l �^踎GJ�W��3��^��<Mp���Fd�lN�Ϋ=�D5ߟ�����@Ж�]���"�x߽�$D���p�w���"��x���u�^˫'*�s7��r����(����hK��o���؜��N�X-t����u����=�@]^��m�&ĳj�pH�����	�$>x2��R����,�J�c"��[l꫍�,�N��bP��@rW��hS��I=?E���$���aubh�%��{�F��]���Z;���W����?�L���n�p4Z�(�b̗�!�&Ϭ�Yr�\�ў��&[c���� a���XzUVE�b%���y�m��G8Lc6�� q�5f#d'UI`�Im7�]u(�,�mаSiѲ�x���C���/�?��xM�j� �Ptk��h#�o�)���+���߮ͽ�nS�l��l𓓙4��#���k�5����y��Z��d�N?7Fqy�Ւ��vb&Z�V�C�m�7���#i`_6��r��.ɴ�N�W����rOF�q���X�ъ���#���z�X�e���FW黁O�a� �X�3m���~���<�~����I�깑G&xT`�U�%�ɛq�^y�=*��;)��z�'ɩ��4���5觋ŧ�G��M�]�_u��m;_0�}r���T���m���y5��4�бzD��i��Hs�Q���b2���@7�Q�Nh�����+<aU���.�ՙA���ԃ ������k�7��	��P�Z�i�?��<�(%�j��2���i���/��[�+�v����P���F��+X2����-����i!P&����:u���>Y,Z�k� O=�d��(��A�^}3�����_d�w��g�����i�����b%���p�6[&��%����¸�7��|�CΧ,�2�@j'��SU�['�E���F��F��m�,�f���~sh~uc ���_���Ĺ:�v��V��zYR[ 9�p��U�Kt]V��`���S�L)x"�?�	�U�Ep�	c1�T���-�=�+1���}�dE�R��[r�]���&��nGN��`��������I^`�J+:�F��o�s�My-�J "��]�OH��$a�k�LF�EN�ό�Zm���>KG4�-1u�2�9��\&6�MZ7=��D�:�"�TSͦ�~��`�8*K����o fh H�'�mK���uN��.ֈ�w'm�Tӣr���mݘ�Ƶ!������`� n޲@]u��R��X��ғx!����Č��B�"cBW��������䒮ŮT*̚�VeD��\��cs�4~���Qiiل�ݩ�r�*�ٙ|�qO&f�d�b�m#��!�3�lt��ی #ju���t|+�*�ס���;J_):�%�j 3�buaN���Ăы!���Ҁ#�ܣQ-I������f�%z�]��&|�i?�L���~���9FEjB�]�ԲN\4��j�αp�ĭ��N�"���z(|S63� ��G�/\�2.��Ri�/�?J��.��m�J-�SH�����̗��M���z�%�VV����Q[{B������f�#4��>�6�<PC���?�~�����Us��$ܖRG&d��9�ri$�Sg���r�رGۃl��C`�RٵQh!�h�A���H,M5��^��+^ǂ�m)��r݈�6ޤ�����b$�� ��ē�O��G��;���w��h�F���H�!<$��% �E-��R��I��V���w%�참�SqYkc9"IA'��7����1���^)�2ԡ��߂Y��\f>Sq;�`�)[@��KP�ۃM�_��^m��@K�����m�s��nV��Hۦ�����Ӡ���P�󳨃 �m�i����YyR��䡆��C;ڈ�i�"���S��-�� ��%ə,��6�j+�ѨD�y~!�t�fm�J��k��Ų/,U�Mz܈Q����ý�
�`9s���Ӆ��0i^r��
jT9fM�A=#GU�����Lz���V��2	1�D�~b��D[��#�
�K���B<~\+j��j���&G���%���"�� 	��0%!����$!u����zfKA;&��Kex,��5��"�YX��P85�J�[��wԹ�����W��3x:)N�FT�2aE2b�������Dk�(�H^�;��&:�7g �LU�
J��$��}��$�c����)�NE|���$}��8�f�|l��gK��3G�ʏV�}�1���td�����Ͼe�z��
�ϛ44���h��y���>���o�ϕ����Eݦx�h���Bd]F�o�c�_�񍎬}�n�zT�H�,=�+_A���GV��:�< �(�*kπ����elȱ�lb��vP�x}�m��d�=��.�ZA�>���f�_��X���� �F9�b��byg��|��%���~��3Po뚸}y�u�0�u��I^%��)��3`fρ25��vz����e������=��pU(_3W����<ekM���J��Xse����=�n�o��vV�O��f�չ�▬�>7dqf�I5ZYĄ���b�Y$�>��#{�t����s����.b�=%W�a&�ʍpGy �d~�j���2�^�%h"}&K���c�5��r$8٩Un�X�&�ۤmdc�Z"�Urq"}L'9�~r*�oz�����;o�S	ov�O&���/�֔�*�z'S��������J>�a�5�}`�v�a�c��Q�������I��� ����˹=�r]�#�G�Ǧ8W�*��+�$�)�.S9ҧ�Zr�G�B浪���`��NQ��QT�Lo
;�5��/��D�_O>����5�<�iU<�,#����U�O�Sk}�;�_�bR-$147s3�f�hT�]�4�)��C��s[u�٥�h/w��� ,�0h	����Xu����T5�Dj��d� TU�+��L�{�M%z�eⶮ����	�\2<�G�A���5$u�*�g�H��$�.��Bl�_G&�"��a�3�G��y(ND��ڳ�J�QN�2�չ����s��,%���m�"�
q�JvJJ>k��c���#b���� R+�1RA����v2r���P	����9��[��G��!��0}�9v��@�@�t#��W7�{c��oo!ܮ�j;�s�a�oLQK7���Ŝ��3.�V�Jcض��O-g��kݺ����ɓ�Uc�+���ڟ��}�����w���	[��͹��u#���9pH)%��A��@�Z�f���!t���+P�x��2\�uSj0�LG{�}v��6�=t�T�[��4k/��g;!GK��M��;�㶀�0�9~��jGc�W̫d���$�\D>�N�ŨYՠ��5а ��os��N�V�x�ǩ��/�S�X�lT E
��]<֑h6'�YJ6�����C�g>5� �7�=I�uE����j��	:a�\&���M4BdK�.0�ϩG�����?��"4�Vv��ؖ"�9�����󁱣7�m@k��.��?U�yzh�����h�_�]��<7�,.�0�tf�ck�de�4j�Pu)��csA7ږ�.�����vTv{���ԕ��!Ԙ��	TE���|�^Z�]�ΐ�����`a��l������*�p�ȹC�]>��
��F�r�|��z�!�LS�^�j�]ml��$xb<�Lpǉ�(���4!Xe�!�|���p��`�o�"���d�,�P�%�ӵo�:��lT䫌��#a���z����x�G�@�N�+[J�I�#b��"C�ءL���F3H-2(˟
��B�8�;t�K��K/���8s��;�������ϔ�"U$̳u���X&�8(���z�|Mlt#��A���I[Y���v&��$<V������=�.�Ş;��M�R�<��j�6���!o���;Gg	d�nE��j�x�)�k0��E�5��2�h�'��q�l28����_P ;���Pz�l������������]�q����m��!4ƕ:v�Ldd�@k�~�B�v�ǽ��6e������R��������_lɡL����鷵��-�X3��p.�|s�f�ѡ��<0t�K�])?�5������AJWvn�ߣpxi1
�y=�����ʯ����6MS���Wf�T�����6��~�|1'q� Oa����E���}��]���Ȟ�_WE���Er�:	e�ō�5����|�f��Rdc#�%��]�lf(m��n�ĕ����7�|����>6R�+� k���*'m�`BX�� FV�i��<��%��z;�}��}�\�h��Ć�k����C�m�攳�@���VBB%9�f�B��>)Y�ǥP�cP��L�
ff p����9�X�����
�r�*�/���6B�@a�M���wu�50(\X�}�Y�SP�J�KLE���YS���jGɵ��$��T'P������-��M��g9�F�YvS��8�σ��oi�8K�GKWN�3g�l��Cp�N��Z2t��[Z��(k���ggb
FZ,v��g{�iP�3N�U� /������ʗx�����:YV�;�Rn��ߴ������Z�er����h���j�V1L�Ƈ�� �7