��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\���V�fnvx��ÍG_;�ȅe�~�>���9�>��Y;�0G�\�� ��|7rw8E$64��c�-Z[��EY�v�5u�͌�A�&���%��j]����K�aK$�F�<�[mA�������uQ#
��`@�E/�i���(#2T��E�f�����h03���>�E�\zj�}�Ҏ	̜K��&k7WD�"�hxM����eLK7�t[a$�kd�[�r�ή�<�+j���<��^���v`�k��W�z�ub
Fl{��iRǫ24ڋ�#p�)�%�G�NE��A���Y��A����1�@h��yG&�
��~���<"?/)Q-Ј�}e�v��Q�I�F�Q&��t��|_c���l�M���^�⃋B
��<p@�4��H���4Hg`X�oR��6��d�����Z�өN��i6�q�UD��^9i�+м;bw�ӝE�'hbs�ݧ��K�Xu��&��פ�obD��e�S�Z������7�{a����@�76��+�(��O���sNc:!����`\�%Yn�:eѢ�U�a4ɘ���L��}��s�3�K,�bE�>�x�K��y�����7�S}��{��zj�@p�0Pd�=|Q�� ���w.��<U�
+��Ygn�~t�;�/x�9׿�泝��QuO��>�)PyGC����U�7�n\����z��ܒj�3�iG?��pb���#�~�j眄��<$3����Q\� � ��������z�34���w cm*I�i�Ʃ�p5�sG�,l7�ޘ��C<D8u��IG\���K)���є���(�J�9���c=��2DK?�J��
:>ϓ���k�Gŋ��ZpM�!p�[:�d��Ha `J<\ƽ��w�Ң���ʘ�&��.PG�Y9�������0�7����K�R$$���5Y�U$�:Ȥp3T�4IZ�O�@�l�׌���V�Z�	0h��0����x5�Y
ո��
�+��U-�q�܉�x:~���,&>ex����"�Z�zU>��Oڊ?��������$��
�g7f\anf��Ë@r��Pq`aD�.A]�BPs�y$�h��?m�*��!O��+����h����HS�ܽ��dF�UJT-'�������Ljb�.��c	�8PaA�����닸l�� #�Ӹе��]���ɋq��v6�B� ����3q�2��W�G�+f���&#�HT̀zhV3����Y��as4�v'��'�1�ra�We^�
qB~�6��'��Rk�Gq��>f��ٴ�Gдm�����V;&���/�N���u*��i����z��3����=�2?ʔ�O��P�qE�L�9~���q�bU�f���b��(!;��˱�#�Gǧ@����<��#W�aX�p��՝�iT�����
���8yF]������x�D�G51IE��.B��;>-ד�,�	��������v�Ԃ�!	�>�l;J��A����
�Ç�l��T�yW>+ ~�� ����\�#!#.rkĿޤ�ց�p���	_:��5i8L�Zvrp�3��#�R��]���Y��Q�e(���-�ʻc��$*��_;��,,=��J�]&5�{kI���XYŧ�)ܕ �&@�j�oy7�w��	�����B���<�����A/R��s�}'㬛�xJL�;%�äl$�|�S
���n�`���	DX��;�P�!̈Ձ����rW��s�`�`ޅ��Df���O&y�-Ou�*la�]���`&ָS,l̖Ļ��[����g"]p}[�9 �2��߉��h�����ˤ#"0����3�Ϛ�HL�6�QԍFբТm�fL�������o8�i�^�JU|��'�]\O]]���c��bwh�颒C���+{�����+Ťq��?�t˨,��9W����^-��o��E��T&+���!������-f��;va>�p>@⽣X�X��E��e6��N�������d2�ZF+�s,�i�F�Fvs*��{����\E���<�<�\2�"q�O+a�2��UA��3 �:����G4 �;�t�)�l!_����Xٛ��l?��ꇤ�b�o��v�;ˋ��&����5�\����5pߺ����A���/���`�,b��U�[��+0�� �9R���i1e����� !��5e��ΔCx`
xS�P��8oLE�"��Vo���U:��J���o{�=�/J
�O�j�m�by'-؁�*ˋ��!k?�l��D#��T�5�7���[G>y�������!�A���1�L~��~8M��N �ץ�}	"���j�]>�޹w(�}��vUͷ1�I��ɔ!]s9y���ǆl���%ѠY�e7�pΝi׎5^�緷
b �ϴ�؟E�҈�}�Po��,��#�D,��7T���u0��ݨs6�0wʒe�v�"�O���A3���B�����؎Ae�	�B���H`VgX��/.D���a-(\�7�ͳ�L\�\H������xvOV��(�L�S����@Xh�;jg$�ս��n����y�~$��l�H=��i����
E�ia�)I�k��e�M�g����`!q*T�X�̔}0��䡵k2p6�P�5n�C�Jկx��fvX���(��->bݲۑ������<b�)��+{/�^�O�a�re�L�RN�7U�0�,�֋�;��-���}��s��k�r�zV�J�Q�Ʋ.�6!�]֡!��m�C��J�U�B2���^Ö�R$/��E<�c@jԆ\���+��Vh�����F	��=�f��������쀚^�_ (9��	?�f�p��v6�<#�G��9gY��}�F Єt۷�)�^;�yV�rЍ;bf��ɕ�U�LC��i<x#�c:�4��MϬ��q5:Ȋ@�7Ee��y&{�[	�&)z�#� ���޳�Е@j!�_-N �������mJ��*(�.�
*S�������5��ԦZb�}���|_��HF��O�V�3r�i��TX�o�l�CKY�w��CA���P�6��Kvz&�h��,�QH�K�Yf����� �rWRj@&h�/#��(�!���9[?� @>MU-kO�-��G)�B��<S��F�P���<�y�a�Sw�z]�s*k�|��� H"85+D�OBZX3�>�m�|X��<LT�8��{}��������i�
�Ƴ��9���������pƽ?������Ȝ�-"C1�mA�}D�G/���Tߍ}�{zo髢�#�Z8k�h2��.s�m�KXU�g�/�� �޷�m˴�������̵���0'ʞlY��]�@R\J���.YV�p��Ln�*�y������6Vk�p�`�r(�3�~��e$�P2�
l봢lyyc r�,0��m=Z���[�?K:k��$3s�l��X�V��b�9�lIz5��9�M�\��`@����t܋�a38�ߛ��ڭI;#�x��UY���_{����b��g���8!�T�O��O]�H��N���+�3���o���I��C��P��~젂��?c�b��B�}:k�^sJCǁ��%��EW6�L9�����J[ZvS9�Z`Oc�VV��`nګH��-�ZOӾ2�(���@�l���&P�һȟ��(�ar��	{��GF.GO�an��UV#�}_�H�w�Q��JCK���x� ���'w��N� ���7�J�����UHeDO-�g;����9Z���m۞õd��h5�*[&* �k���2�\�6(�`?��c�΁w/z�eb1iE�Yvm�7����9h:��d��܌=�
���ScB��0�����P���qi0���>0��z�㧀�ΏWք��\�Je�%&v\^~Ǘ��泺���zCd���CR��4B��V\>ƄQw]�/3ƍ.�����
aC�F) `����<'�Q>��j��FM#L;Rf��7>J%e:j�Ā���Q��%%Ҹ����2�3��K�����Y��LXq�����xr�~n*���ۭ����ѓ@�{�?����:<XJ�Y���ER����6��w�:���[����'=8�����=|ԴK�y����n���Q �ݹ� #���e���0"���2����g��%��_3�U�s]�����3~�'`?A)�>_��U��YsJ��ԅ]��j�9ʍ���6wuد��K�ms5hᣑP]e���s���k��3�]�YZ�յ�*B����sҊD�a��Eo\��"	8�.#���GRԵx/��\��pa�%W��ND���CB;�T��冡�L�1�C�G�&��wL�<Z���ŉ���:�W{�#�򦄥&H�K�KT���"��O0�"�'��4�saΓ�ɂ.= 1�����i�a�~u����k�%~$ݬ���_�y�['E6���/IMe��3j��ZB���o�\�g��Xf�5��"� �_Gt(�7�;�r ��b��i�p7i,�O�˼�=��>nF�� �Z��!�$�nW�� t�f�z�)����%�/��ĝJS��+��*��M
�f. �j����JZۺB���'7�on5�J��-?"� �҈Wc�����"�A����?0��\5�����ܽ/%�����Yx��mp�4���o����/?�D2H2g �ʸ8��owP�{(�M�����d5^Qž�B��%�`�' Eս��M��Ǩ��*[Ꟑ/�VR�4^���$�v	ևbZ�GÕ��&� ��S3�K��O5b²���Ma�f�U��
[�!�;(E�����^*3@q�1�8��D.��t��.���Lσ�69�1�Bu��z�Ȯ-j�cS7��]���3�)Nm��q�C�.-�����M\��K��N��=�	����8^,<8�'��ƽ��r�-�0����	!;��7� R�U��uKz�d(!�,�(1�*�~��HF�cr���B.q��B	;����D��ԑ��V���d�lX�����7`�k�����o\<�; }��� ="u��[�~�F�NRuRF���#P�\���^	���9���Q
%~�d��U�>?�L��nI�1�}~���i���@���
r+�S-�T!e��;l*�2N��B���jr�	�h������N�O�w��'�h����U)=�k�1�_7���Kq裡��
�!�� ��=m�-����y�������.�����:��5�� ��
��{4���om���(M����|e�
��
���٫�b��,� u2rw#ݬ5��a*�h&.�B���nٵ�����
,<�����j'��Z������S�v鰲�5�Ø�yG�.å�����d�'qWx���:���;����ŏؓ�g���`� �'���\3�};,� �( �ݹ�3�%4���"��O����U��{�6BoO+E�S��k�w%ā7J�b�8���j���x37�2����VU�)ў��p����U�d��#9:�˴-@c��ʼi�!�F����/����_�~���XX �K!�A��.[��W8��U��t��,��_�K��b�%y��{�������s��I�5,`$�����ߛ�F{:{`g�uv;������K��z�qi�E>qM���;���΄T������w'���$@V �PD鍢�?;�_�P�(���rsx��ˬ\��/�����`
�v??X���D
��%qs�=��1R��َÀ�?� �+��mu�?G�n/�`�G���I����Z3���}��\��uq�¬�2��D�n�����
���d� Y�v�tV|���[]p�J�дݘ"�Y��pQ�u��SF[���W���A�����@6Ч��y�S�E(t:�1��`E��h�E����>�b�<VF��A۵���5���j�i첣�&�'
�XPyXy%�佅�U8z�T����21�Q\��y�!7�WX˗������*�����Ϩbkx?@�&������Ը�./�5�m�a옘u��U<ݽr[��>arV`y2ڏ8�k����qct@��J �b��;����0O %��ڴ�8�T�V�4��c���oJ�~"/7�~#���(>Yz] {�t��5��=�'�U��}�ۈ'~�Gc�A%4��cY|l ��߭�c���q�_,z�����$��+{^:��	�Ѿ�hlJ�q�5���d���K d����5؛kC�����[�Z�5�C�Ȳ���Pb����8c�����	�9� ��S��D�5\��'��Yo����������l��L'e�|����0�S��[1>{��@�Q��0#���P��8��x����W����=8���gXo��v0U� ���8�VbY�T��@�*�2S-��P-�3n3�+�����j���!m�:g-s��g�z�r`L�/[C�A�f	��$�޿ҳ�z�kg�ʈ_�"-���*� �JƛoP�D������z)Y/���z���,`�^ntV�8y����?/U��;�W����s��6�3B�����-���ͫ���qT��Q�$l_�]����o�,]j�ӆ��81|*	W��Y����t�|nl�'q�W�F-]�{�������î�:�v�B��aʃ�냡P��n��)#+��䅕Q���'����>��bkz��v�%�|,�����l'��@X��
)�����.>���U�,͓eh`^I�E��g1٫��ĝ"t�ܮ5ސ!'���Ok�����&�q�s`R�9��(�q4�4��Ĩ�y)EW��6��5IVg;���-V�h%'��N�I����dmUm��C��F{
P�i���V|��^�(me�uP:K��U�q]saHQ�qq�Xי�~0���ڜ ���}^7
�.���9yQ�����2�1�v��̧H�����T�]��F�Q��M�_He=\D����Z���+��IRv;�Ǖ�z<7b�j%���?��Tx{h����a� 9�0��#\N���"=fsO�'���T�96,��!Ѧ�֧�L���}��V��RoW���H��-�K�`���r��y��EhT���?j���t0PK=��})�M��EH��L�����;B�|�T�C�4���HƆ�Fl͹��a�뿸�(<�L�=�����*?=��Y���0���:�1,���%q������
6�>��k���iD�6qeG����L-���C�������!�R��d��U
��rj-X��f�}����Rx|���bw�SN��\���#;,�V븶>����O�L�Ș�����8)��������7�꒻h�8���b�;��1��nZ3yh�s�*?����=g�,5��y����bw�ُ�[`Y��4*!�7��	�:�<<���8.A%�2���Ź�C�?�T ���̪o�C�ܩ�)� �C�IϻE�(���\�!��Y���V�Aa�]̗TQ �p~��h�r�sUd:���\��1���x�9A}�4'�=�(��$FB\���%���&i[���r���4��1�H�0N!�Z�WWl��Pb-�'1�
��y"�3�Ka؅��Z��1�|�0W��aH�_8�TH%4
S~��U1��`Q���כ[5q� f2�pf�[����ij����Py�xΘIŠ�B+n���ϧ\2b����IG�������0!���t�����踝�i���+�s�_��1�09������-ъ������/`=�Y��\C���9�͎����Y�i>-r�X�;���"s��A!�E�R��S�9.�4���H�%Ӛ���gR ����Fؾ��&8,��E��Q7Y,���O��-~����ܰ??B�3��ߙS���
�V���-�HW�m. �d!P�T���g����j��ս�e�	}D���R���?I�	����\�v÷�����>���^�G�0-�M�3%�"�  ���,�֫a��͐����\��/�:���0m��$�Ԣ�8��<^���h����٪~��)%���5@#$�o��^� V�
�{~9@^Qg�i/m`l�/&���x��h$��6ވ�R����X0]}E���T��S�P�(�����H�f�l���n�"��k��髦�j����7���ɟ�m�f�: B?r�
S���!#q�\hh��_2�?��+�)U�)P펱�~�I�	6'��Ф3r������;\V�O��}�r�gvv��iaYb0����劕�_z𝩉�;���þ�p�o�V9qs��]#y�����DV�K���9����sS�ͨ%��U"r��[�Dvp�7��W1�A�y�GHsqf��䱻=��I-�y����`�Ӡ��~�b�|.#�_jz�NS�C���\RՈg_��ڭ�|���a����o(o�I��$�44%ă��Ge�,T�,�:(���г����{��F  ;��������Vk�,���*b_EYjs������{��=ʷc�&�}��1�2p�i}�3h#��������4�߽Ӑg�,�ϓ��KR������Ԫ�R�fd3���f|h>�Yc�&9N2���ج�H*Rϋ���>�ye�z��siv;T�����Y�\0Ͱ���bf
x��k���g�Z�|yÀ�G�-�ޒ����{�J,b��x	>�\%��@B6-/X�bD�����.S*�5�ܽ�g� q)W[(;Iy�m����'�!䙤YQm�y:�ly���n�VՄ�R�q
o����s���6D�C<�d=U�� ֵe��'�Eз�%��;;�Fci�� ��-UA�w��ޖ.!>�X�)���BӐs�X��*�e�f�J|Q��U�Kh�yG�C7����*_lƮ��5��U3��Q�o2���Y;5*�/.� V�z�� ���&�C;`7h�B�gcOFK@����hK�H��?z}%�+�P���(�R۾���Yy�(P5��U+��j�dN��:AUNϞR��������y��02�J7�2�ɪ�+p ~�5UhC)H� ����f�H�y�����3Mu�N[��
�8�A�>Z"���dd��|��5��1��ˑe�f��c���p�o(�*��"*�-�JЏX-f�U�$��[j�(�F������¢���v�w��N#[��+��8�j��p�彈C����dD~ġ3x����p}��h�
]S= ִ��	N�.l���nU�S�T<H�&_	-�VǼy��L�rv����3����G��3��u�����0A � ��"0/�"ؗ��
G-�LV���
-<\�V+a��wI������ɵ*P�n�6��N�$r���� |��"�=���b� [��/��BLj�'\
 ���J����&.�?��M2=ӠE����P>:vE�� 5��hd�'e��K��~�[,�u�jD:+c�� Dْ�N�`OUBb,�ڍ�ȴ,=֯U�ĸ��,���Xעc���k�-WB��1$[ 0	?�YzG�Ճ}��6q~&}ްy	�f��}��<vX�Ke�G�7썾���?rbV���I��j�B����Iu��R'f�Q�/{��/�� ��w{��t�R���-lǭ+�W�U(���Ȃ)*����Q[���z>;~����vˠ.����s5��э�i/T�V|\X<�WQ<���C��0?2�Q>E����>l�4��p�VO?�J�����-d�{�Z�[��w�jm����ǎD������f��s� |���p��I����81��j����)!5s|B�L��(r��V.~���{�E�Eu"�S����+3.�O�"'���lޫ��g��6����؂���S�j�ѿ臰!΄e�*��zv<J{������6r���<.륵'����~�4���z*U�7n�,�M�B��	�>��9�� (��6�1E��K����N��LR����,Yޫz0��{�>hv��h �6�'��]=�|������T9�\�eA��)��LKHd�i0�:;�B�0u��A�=�h�M}��Ɣ5"����p�|���ȒM��B*Nޮ���en]�;�mD��Q2p��se��p�Nh��砂)�>P�7~��֦>,�C�N	9سB�Q�[$`�G�f2Ryb ���q����H�����5H3l�b�??r�ѯa^�}����$o<��m� t�N���`������h6^h		��?�%.2N��e�q���Ɂ���m�	x'2jO�a��h"�f"��y�Bn/�e��1���+�K�X��P�+2�c\޷ù��E�H�ը��!W|����z塈��ϙ=�ҢP�3��%�)P�M=M��I�e�C-������6�{�B?����¨���ه��%t���.�c��`
f����lL��#a�9S�N�yF+��0̼��e����Y���+�p.U�}E?jY��ʒhH�(��%�� ����D�GBxZ��;e"��R���������έ�s�^��yI�o��~�4�������tO��$�q0��Ȧ#y�,3YDY�Ov��j/Ӊ�����o�� �uS��4
���?МX-�d��BSW�I+aKȪ��d�ۗe�,���l���;*��\wq�̧O�ZT�]�K<oI�
���/G����CÝ9�����;��fI�����T|�փ<F�n�ө�Z�QT�g��0��Q�v������q�\�]�9�[�!�{ґ����%�ٝ�-X��d�T8��Bhe�桨lͩ�v��M�����WE�,I�������N�����Bŭ1�ظ���f䖑9���aX�T���#��G��OP���͜��	�$BL��� ���H����*�7�Z��AЯ�"g�i���03���^"��s^C�����TF�-��r�����j��j�t�2�y���/��ĭ��_��,~#�R���L��V�0�'~*m�Q�y5��%k;�+5�_u�k���,�7����	�<���e�Ь��#�(&Q�,������p#��~�ƃ�5:ԡ .���:�Vq���/�?檱����ӰA��S�+�����k�0cK�e�NH�)�@tW�xj>b<�ݟ�VJa5�|c�Ku��
D�ȇx:��Q����L� ��UOM�h��"�A����ľ���SR"9p�����(����<Ϋ�U,�����{&]4������RꌡOL|�u�?������"ή����	8�)�⚑ӍIE�:ޤ�iUDPh<d�%�PC~JH�I� �E_�(��Z �$��&�!L���m���,�6�����yA�2���~of?.=+!���?�*ا��2m;��>�\��F��B�z�C�`$����x��eة�^<���֜�}���$ �zLfAH�bg9d��g�:�|��%��)r1o�6�(��W�|m��C7��h�P(l��%���a���x%���o#�i��]����A x���G�yH�Y7�+)<��t�Ak� _��ɱ ?�9�>�K)�������ͧs���q8�7�R�����-/t}����<+�S	+z2����4�eP��?$+ڡ�g�X^�<4�$TT�퇻Յ�/�,�*U��Z�"�B\��0h��  �X%��T�fP8:��)��'��4�����p�qO!I���\�+,�0U�:d�� ,!>U���
?bQ���m52���l�BQѧ�"�t�@7��xΡ�$E�FYE�4^�J~����.
��6��Z
�{��_�ʥ,��g�!��وj�t�E���V%�lH(6��|D���f
�`q^T=҃����'�A�Қn�D�l���}��t+�Cm�����
ŭ�V���FY�/��sRϧ�D��J���:�ǡۡ ��v+õ��l�&\~)�∩V���K��>G�`6���ß/�oV�=��73~˃=G�������.�'o$��v lkD�8���ͪ`�l-��6�f�iF���*G���i�)��^�j�\م�6k�� �\z��<���L�H{�pV����N��_�}���èB>(��u�f�J��M�`���6J^�=p�� �JR�cc�s"�J����@,�_�h7���_�t��f��q1�73oO&�T���/|}~��q�̛�a-z�NF�>�v��nn�Y�ɝ�Y4�{qe��$�Ca��ɴ�s��Sŷ�?�7#$�>D�g�u=���WF7�(��#�����%����O�	ׂ=�ʫ?�]-��v��KVc�q��"x@x�"�����5�=TF眥��G��|�i� };��x�㮓0⤛�K��C�u����>��g��U�#3�nT���0[m!ˍ7[�^��z�q}'K��_�s���%���Ǝ��r1
p�K2����¶���֢��a���ᜱ�~�9#'G�Y >x6-�(���38朽CC nr1h�v�7�3!�%��r9�F���=/ո ���Qg#�+9�]�RT� �w���#��W���T�yB�t,�?1P��`��\�0/B�^�٫�C� ���1�f����#t�V�[�%״K9sV��hr��m����[3P�{���Ai��L��'�o��~p�Fol�2/օP�[X�(84��s<��$#[Nm!���a3��.l|��7ا��\��G�������o~T������]Rq;z�Ȳ�[[�Һ�G�������#�ӟ��5^�<o����rB���u�0�V��L���I�ȌP�C�����;#�u���TOG~��9N�lÏ��7�"\*���jj��t��{�Nia��7+��My������UG�re�&�<���ϋ�I�,n��Ͼ�~���!&���Jk.l"=���o��Ҍ��\�К�ҡ����2�+N���?�U0����{܅?=y',|����gf��b�.�K����=�c7Fg����,��L�Le�� �<y��X���^=��$���pH�t�׋e5`jc�m��o�i_-��d�5�b���0l�n���^͔�&���(}5ut���Q��I��RY�b�l�3l$h�����2^���X�Q�S�)���=Ɠqj�_�EWs�MEVa9R�Hd5����\�����<2M1�""k�����Gͷ��% �T�Zy�kI�[Y������X.��\���l�����\o=���O��u����� Ɉ��Q�uG����"l�2�h-��� @��pE��;��4,�;���K����UD�6����u�mq��^�G��W���u0��ت[����`n��IW����A���A �{C��Z˪�V��"ĉ�6�g�DV�R��0Pk�Q���B��뻩�vCFx�"�ߗMj�'t<r�'�z�yL�F��X�p�D�w�vΚ~�ʇ�L��j�o�@�/���G4�鯢˶���� �S��?2�����8�KIaޱ�e4���i���(�]��U���q ԱG���R=C0�P�q}��FI�j�">Y[�����*��
��18�=�.���^&Ep�㣀/-u�0h1�����-�`��>e<|������r+�|��T�qCs�!�y�y�q���0�Q�Oa�RC4�=�<���;RPD��۵Č5ұ7��)�����$�J#;��?�ͼ�b
+#��|��|?�4�z�kc�+�t�#9~��5F6U����QX��=�)�7�0z֣	?䟭�bɧ��R$��Ew���l�4~��^��n�æ�����6@�y�����j%w���[��=~��Cf��#QޙC���0Z6%Q��&��sx@cz	o$w>����ͥcTW�G�kR�}�
��l�7U�<�t	����X�7ּ���E6."�[ꪓ��JΉ��fsE�|-�:S��Q� ��F��c�:L�A�]5��X�W���N���J@7
�#�9!�<�b74,KK��ۼ��2���4�v��^7E,��˳jq�����;$_���F�8'�ƙ�j��PD��� ��<?�m���'�S�H%# 1��Q�JH�"�>'��\ ����r1%�O�M ���"&����.St�7��Xj�7��?<�ړ�E��	7��>�L�"��":�.��rR-�:+�/]��������!�}�y�]j�hl�1�/ ���/ɡ֚	�=���(u<�� lS��Y0�Tcջ��޲]��*/�%�5�ٹ�(D���?i����4��8�韎^	��-�1��
�jSm�etH��O�}:�/V��(߇�&�v˗Bl�^��w�v��E|W�! '>�a��u�d��{�l�׈Cŭ�.xʭ�|��=g<��,$ba��v��8�$;�B��])��KȄ�\�B��`�e\�՗��q�b����`�x��
�n6�S���锷�aS��.@�V����a��X�
4�*�K}iT�}Rqb�|����.����S���o����nI��>����s1,�:#ƶV�k�9��`��b<8h���٪'�.Մ)<�)�0-E�ƶ�u�?�j��'Kh������$�<�v��z����%�����Tq�>�4����sȰ���֤�ɇ�s �i"�G�B�#�z|);cY}�D�-.��j*�Q�ri�\�]jѨ!`F�	T�r,��ʙ쿌��'67C1^��E;�M
�Oǭڑ]�L��.ɼLRrU1h#��h��]t��<6�mP/��]̇4S��L��v�O}�C�B�<���;a�@���C%ݳQd�W�A߅��t7_.*Z����n��u���Lp���ٙ���/t
\
d;/�IG�ۼm1\��xjr��C�I��э�2S���Jg�_d�/�WX$7k���� ce.���2����^ź��؝?k0�Z�/6[)�'tr�ͷP�^���]D-/����T����OF|.fͤ�5�I��U-_��0�<�eCF�y�H�P��\r:���l���ۦ�5�A�ua¶�'���$��i��;��ܴ�^M���v`�/4U9_n�a��	���	�d�uP1*�.���(��]�2��}� �G��^��4tw>����đ��0���;9?��`�J&����:�l�2 �H=��˘�>��vi7�-�*A'����^�e�,�q�w�/J�+40��K�1g�
A��1�k����Ɵ�Ki����2�4��Jf8���s�!B��jH�Z;��j�'��.s̗Q�OT�lxP �5J�����q���$v���\�c���6q(uQ��D����wY�ı��ś�u���=m�y^ʲ�`/Z����h��Q�F����U�7�7���V1������D����e�&�����v gG1�JMm;V8�����7y��o¸�^*�J���)Һ�=j��?��F{&S�����"o�?�����gѮm�=Ǩ��1��w�Dݑ���6�.���z��X%Y$�n�x�C����Ks�1 �~.�M$�~���!��,����79�V���Ww��C� ͔��Rw=J��q��}cѸ�E�p�E{)5�
<�]�N���%HI����)�����F,�y���f������Q��!���(�#,B'�{�B�UF��\s��T�gf(Ǔ���^0@�ٱ�|����]Rz1�k�H����V0�1�nO�G����V�q� ��e��Zơ6f��*�Ȼq��-�ÃSz3;�aR��h�6�����CC�J>b�o�	��!e$�C��u�_��+JB�B�9jP�W�SX9�k27q�Uj@R�Qc�-���`�'�N��{���iun.��B����f������ܧe�k��1��UT�nzw��E]r�9N�*��.�tZ���c������+�MMKn��M����RϢ�1�<,�J��HS��0ǉA�p���f��U�q:�Ŵ��v$�b#,���Mz�{�J��j9W��#,�� ���ٍ�=%�&�(�_����b���H�.�?2�>��ŷ�G���a��5����vQ�Wd�N�w���I�hYÑq��yQh,gz{��Z+/�x�n�urr�&er�gH��E8��_���Y��U���΀�G(\��|R��ԁH���2
T�r1�N��P����mBf$����(Y9�d����7�gIn�3OJQM�9[��7���jz���%r���\&�P����h��㙈��,��{��/Zh�&j��~�Mx��
�'��Vst�Ln���$䷲����|������)�ɳ�7R+jځ�a���;^����AY���\ ���L6W"�6�\����xg�z�p-�B��a��92Ў����#k��s�&�K�oF��u" �R�:O"vDg�[?z��CK_Z�`��)[��/���ca5xmW
.S�$���/�==����v+�bVi�7��kDQ�o����[ �!R'NY�k�����ph
7+���噥o���6?C��M��7���w�ٌ�ឆ����|K��Ҩ�^A��^���,�!��LA�7�ޠ�|���:�v��T����43�;�	�h��p�;��6"bε��rR��̰P4���w`����]�G�f�����ۣ�j�!؜F���vs�a�>���V'8��W��.�K�
nփz��u�%r:��]�!��ݡF ��:L�^b`�Q�H'}���iG��}ftv̕uS�f�Փ.�~#�[�X�K=��%�Yl��s��%��e����«�#宦j#�AN��#��
���*ܵ4�/���z�b�6�N}��E�A�^8�jt`�^���h���ó|RE,Tl]N��O�(1�,�~� f�]�(K�v��`[���M����`�Q�����ѻ{	W*+)��c� �*��N\En��&�x���+G�
`!���t8���!7��ǫA9˷�M����vܫ�z���!�a��[vH8U��v{�8J��|�ڊ���<:�nR3��A��O~b��j\�#���7�[����oqZYN7R��6�D�]��p�r
���R������:s��K:E�ᦕ6�C�Oؠ����#5����a>�Ʈ���£e7Hz
0���-��O:����Nç����j��J�B�er"��ܩ�����P�\��ӂb�
�g},-L�dNT�P ��5�\��DA�k����EJ#�T#~�>@�|�h�U���hNI�<(F6�K�`��r{f�|��%�ȿ�No�~�)!w�s!��<�?/ߔfN��'�gM���Ҷo�X��_�a����aB*�����1��n7@aL��3���@���������P/j��A�_��c������|k:is+x+����=v%'�L���aȔ?��.;Fx���s!��`��s�
�[��kYq7o2��D)*B�V����y��"���t�2̓�[5Pܒ�l5�ro�������o��SJ��r[G�%����K{�O�����z%t��!���{�_k/M�� ������Bl'y%������0��-,�*�(e�2-X����X����Cb��0K<��՘���,E�ӷ?l�2��Ԇ0|���JTJ׾��US�<�U�[|��ʍM�jiI��xxv|�g(�r�J��#UN���q����r�#�7�-�Pc�V}�l�m�3WV��nZYU�@c���U+���N�1=�,�����qRW�+������G�#�˺un�#� /��V-߂�k8M-�΃צ���"�j�]z@'_`$�?U7�Z@\�9##�h��L�xF�:@W*E�]w�3
2^>�AHXg���u��cŶM�$�j��� �跭�+J����B	�f��^�J���RW���l'��P4Qp͇�8c��`���'�~���v����z���z���?R3�I�L#��v��Z��w�&~8�Hx1	�bd�+���%p�}&��0�>*N�_d���{�S��ܾ�
��u4=������*�}�{7q6�� ��^0B`&���ʙ2�I��%�Z��9��~������׶��Ȃ����יH`n��,E��7�d�<�rƔ{���Sn�m[0+]+��a���\�8�vq~����E!v�=Q�N�k5�e�QK�|:����y�m��1��i�R)#�B¸�@x;�t�9��`��e} /�.G�d�ֻ1�U�k��d��Uz�ο)��i�/Sp%a�[x�bă��⥈`�i֍:�xP�[�^M�1/�
�xq�>g��?��ҵ
bw<�+n��I\Ł0�����Tf����D�X���q� �[��%��Ēj���@��u��c?S��6a"����^��*���܄|xk�M�&TR%����WSl��
)l@��-�q���z����V?=����}�!�}��������g5�f:h�+�����B!��"�$Ϙ�k/�@��0��q�de����A��$ ��#_:kB��_��2��ߪB��{���-�E��;\&T$�T�}M-m{��r;�����v,8��a�-Ԗ8ʤ%a���2��)�(�VG��tD�69Td��V���k�0��Hm��f0�$e���o#J1�G�]����9y ���foz 
ʮɁ�
)vz�����^�MMf(e�����&+�;$��֢d\����O��w���W����O�\�-v�;�8fS��-�D��1UY3��J��B��!&^��z���%�ӍaL��>[� �^H�ȡgz24|Ƌ�b�_Ӑ���Ӻ���;��N�u,�Ԏ@�I�8��9�=�C�w����\/��q>��2�� Ƭ�b�/�>���r�~�
��g����4s'\7��z�����V�d~��n8뿉C�]`aa���׼!lj'�e��~s�>�[����ŅT�JP�{�co�<�ʋc=t_��� g8*����1�jdj��2��"�r�����A��`�yG�l&D [ އ�>�{�W�H�[V��\�I.�ҚCPGHd�:�F��2�����Lu_�eHf.�Z���k����a��iM�X)l�}�qz錦�0�2�Rv������r��L��
�; J
��X"^�%�E�0j�8Y�iI�O�l��\}d[���}�)�f�r��PKݸ>�rV=tOG_٬�r$�Jl��Q�����y�P9�qYڱeo�<u���#y�Y4!S�O��V꿦< �f�������
'���a�@��f����4upy����V��j}�P���Th���\��#�6Ć�P���2�N%�`\��c%~����$��V)½=}ON�]���"��,��H��}!���vTЙ���oB6��D�	�[��7�x������p�EcMg1���'�wjE:�Nq��m|5 x�������.�!�i����V�,����	
N���eys����V?T��3��4#�2�&Ϋ߆ 4{�%0��c��7�n&(բY�����C��⠜o�p��@`�b�ė4��H�H]��$0ְ�I|��gH�e�h_�/]ò,y+�]�k�鏟���0܌�O�U[U�#xF��m�6G���:��7���"a/V� ���I���h�I�*���nrY�)�*���*���Dݳ�ޫP�cKD.U���8�5�X�Ew赲$�j	~��"��V�]�r��L��[a�!0�6V	蹺��r�o�З��f�k�J��A�3�y�)s�zW��nIJ���� Rt#E���b�>����jDj�TMFF��A"Р�'�
�/~��(�4����U�xg�>����X�\d�����gsߛ�;'�k���ޮ[�驿=�*8�lFXQ:�]G
�pM˂�)�R� �?��\����	A
���R�
�����x_�
���j!�?�}���fb6[w��m�H��vz�.�J��0X9
	f�`vm�`� �e0NK�w��	Q,$�)(�	����↥������;��4f�F5����nG�H�"�o~��:��'���AD-��f�yD[*�%�u+��`Et�[?R�F�؁�I�)���o��iPSλ�v��Ǔ3-��笣��[�?E	bL��/��]�,;u���>/������B?�L�p��K���
���G���ze3�bY5�S7i�Gm��HY$>5�)�&�-��Z�OE����l*�"&���'Tp���Z_��>"|���:��yJa�}T��I[̋�Z�սT���!#��[���<�{�l�����-���5 K�v&g�]���Fs\�͐�C����A�t�(�W$�}�,l���,�1�� g;T���ŘE�j���IK�1�~=JHl��ä:�>���?�`�:Y����b?��~�m���!V§g{!�
'�Y�+���SN�Lh���N�,�%�y��n)�ۼ�p������ndn7��P%�������va��Y2�:�#��+��I�_�m#�ϛ�Ƃ3���85�'���`-�y�-(C�/�P���G�X_�K��~ו����{�Sm���F[t�d��3�b�8�h�q���ڀ���ӝюrӰ�?ʇ�-�����+'h�f��M-��Ѩ��_Q��E��sB���T�*��Sψ�)�/C�{�r>�,�0�J��=@���)8w+��j�W�
ޏRp�~X����� �b,W�cv��'�'Gk�W��Q�&xo��v��N�a�Tu�x�_E����M�N[�ǆ�V�çn6b�o5_pH��C�;���N�M��y�O��a�uX���|�{V�����q6j6�l�`�!����d��	x�t
�S�5��B���ӳ�N��P8�K��U��;pnfЬ�`�������
'ڹN�:u�װ�!��_21
����h���:J��I�������ݳV��a}���!��;;�M&���u�ә��pn�'*U���M�\(Ȍ%e�Lo"�ckƨ7���a�{{1Ĭ�D7��r�S�ܻ?r�� ����Z��
S�=Q� ��r��T�`�0?���m:��B9��`�V����w���9������Z
�+tR��,�*��>�ۋl�$3���x�������5�o�����hj�ؚ������M��?6�O��tʬ�D��T�p!���at�pk���M�v$4)��;i������B �0���E1T2�	�=.`�ڋʍ|Ѥ�ފ� �'g�ׂ�+;��:�9�*
օ�J|�pՉ��J�2ݙ�L���g(�̢�T�/�C,������0�)A;H|����9��E.C���:Rcԏ�d�(�Ƭ�rH�!٥FX%i!�q�;w�Ƭ����T}���`]���u����RsYA[�iCyN^ٍ�3�}{j'q����ߡ��2�2�]�ehP�	�S(Q'کx��QL�c��?a��ꮿHT�%?�_Gb��Ή7�}����:Rh=�I�!4&_ǖ0�I! ��冺s^�jE�p����R��+��s�	��"�b��f���z�*���G����A�y�:Mx�D���Ùp-��v?d���^C�_�8��������گUg���Z�):4Ds3��b�w�*��l�4�B�n��ȁ�#?{.�<B�5ʯA{f��â����~��	�֡�:,MEB-H%A�]B8�ڟ���1����c�ڒ��7.0��nq}�X�H�j_呮Ђ����}w� �h<s��䡼|�j���Ф��@n���j+��ܓ����l'7�Ö��(�Z�̀B��C�)!�β���(�G��b�E�돵��ς�yݫ�3@���h�7��Y�=��E�K�J�i3�7j��I��@!��
�`���%T�[�a� �,�w�`�On����}"EM��I̘�*���~ﳃ�{񞒖d)I'̌�����q��?�VnQ9�]l�e~k5?E�)RBEu+;������^�������N�$�a}.�R����}�]���%���k�tG���Vw?.��	p�\���Lcsw��։�pOS������/��}	O�}�u~m���"P:A�u�6Pɮ�_�-P .JS�	i�݈�e5�he3�,��4��̍��3r(ܞ�x0>�\�7{.g��F���]��<��t!~�ίD5���; j�9���b���[���9ڬ���m�� �z`O�5]5��$�W��i��gkՑ���+��}a+�ԕ�q'���h���O����8���i�w��3���@����s�}���M��IG"b,D�.�f"¹C����`+�%g�?��:c{hy��y���9y�&,tFO]�x䲐ӝ��0���jro��=��A��5���f��da��on�7H+���Z�����Xz��U�e���g�|��(�̏;MR}��6A ��ge�]�͑��C0V�
T+ �4	����+5#��|' �%$02�F����-��g��\�{R�L�q#��B�i�wN�[�w�F��f�"���ڴ}8���p�Z Y`�>���0�؃.����tA>�]vien]�΀F�7�U�}�(\{-��l�b��� 9�2k�����f�E�@�!t@�!��ٯ��M���D�L)]��-u�,0�V����C*�'aH�P0���.$9���I��+*�o����3���0�_F�`+��y�*
@ZV�R2Wt&O���bdY@���:d�Grn����YBu4I΄��c^i�L���Cо��j�����Z�7��v�0�8;�C:��n<'`���Y}/����x�pf=��{M,�`�����Jz�&�F���{��&���t|n.<&*��sF���7&�����6�����5��E�~de�ىo�9<Ɍ�g�(wB���Q��qN�=����o�g�.���Ud�}R1��I����6ux �u_���ΧD�3P���41QN5�Eb��I"���ȫ�������g��D���_yX�(�5�pᴷ��l�D_�R�E9-ߟ����d(�X�-;�� �n��T=���b�v"�\����Ӈ*�f@��a�S�-�\��k�����90d�;��Q�)�
���=��C�U{Seq���y�����c2yyi�)�rGJ��a"Fsm�C���5�)��o��[��;ׂI#�Q�ؒ!g����8�g]�Q'��'E�1J3z)�4"J���:���H�A���=-:Tz����r�.`(��W&4��1	?���@{�`%�I�A�n5������WQZ�s'�]r�j��?N���v?�S{n��(��;�>o�l���r���������֧�`7z�-;Ю�[�+:�<�������T��`�8��o�V	O����a���ak�$��/������m���	XA��"��aE���"m�����|�o�}
��`�$�}=�X0��œ�K�	c���rv����5�ק>��u�=�@v �j˅~�ع�sȇS�1�t�~*@8�����W#�f�*7,��Y�������?3���;"J]�̬�D�Z4>�`��@�2C\�a`O0�I�XV�I,+�׈#[��[\�H.c�<t�s��X��G���
V���c/T��C���.Z���~���6/cl�@���-����q�	��$ʹ�}�(/�`��Cu�����N �l��ߡ<9D��P�	S�0��r�Z�y{rl�E��리M��z��[lc��⾶�d?Rn4^]X�ePRO�=�V��+�<�ZT�f�M�@u���2~��E�0�:������J�/ԍ��pmD��A�7짜8��c�-9����P���q�0?����q���T��365N�����t $��M�rT	WP�mF��zy��g�����XN�hJqO�����T/�P=T���W�=R��-[�헛����{�6mF���^%�yy���,��`�52�k	���P��]�Z��b//�:��C^o���F�\���tg�fvWi�Ժ���U�����7_�uOg����d�ϠOc�r>0i:A2c
-��C�J����d�?�PY�3�Z��^������7U��)�?+�g��+�G>����6r��|	Ko;.�;͏#�ڼ$�7�!��l��*'��g�S�iE�N�:=�t�T��f�:aZ�&�P���������%b���θo�����U�5kd���}�7�ے��"�rTŮ���_	V��N4��4�!;�~���SX�� ��
\�`pl[����h���\%b����ZV�,��.�B~��⵼�s*)�'W♶����?�.:�m��v��ԙѯRuϲ?kۘ����=� HGՁ�詯X윹��V��~�*�>�s�9v��'�غGƴH����&�v�	�y�p��Y#D�Q����&A�b섊��	�����{��{L7�����:?���$H�+!N8�|wt�M�6�\m<﵊���F��9�Mjw�v�a�2e҉[��B`�|�>�y^� Q�Z�����$���Qxr����Q�G,���g��A붇5e��b�_b�م�X6�`�=:�9�	�3�Z��%�w,2�ׇ�fs9N�ŽTE�RH]Չ�yǮ�}S2D�*7t�� �i؋[���J�Y��V�3\�ތY�y�T��.��Hm��`t��Ӧw�A��80a����l���JȽ]<�7�""�!2�X���¬kU�|�����v�6�6��t��TwQ#/s,5Ե�JaбV<���}o��кm�w��:QО)x����|��s�R���bd��o�*�km�E�#&�f(�@�Ԍ���M�H�����Z�B�-�nL���5]o�Ҙ��Φ��*�_#+8'���e'�[}�M�1�Sd���S8�6���O�
�G�{:����Q������C5s�y�n���l7�5氅駴��y�����@u�k�3k�1вL��	���4�/��@ƁH��R�~�9�d���;`1-�4&��b��l�M 4HS�)�@Oɰ[��8 x� zQ�D���v�
�y˕RY�ޟp�Ϛ=������Ƴ���^�H�4�A�y!�>�PDF���?���h���?�|i6�Z�]nZ�f����=J��)x�Ɗ�&�P@Q�D?��N��u���Qs[7��6 �x���X�c��e:�]@!θ�]��g"�f��g���U)#����p8J���fҸS�hѷA�����zX_�k�[�2�y(A���"��@��
0G�,{����1-��SUϷ�����^p8��{���FV���@P�[3���w,^LT�]�U<�cs�;����6��]�l5���<���� g��R�x�h�cb�_AoS���ù���9 ���N�`�+�Dn�����_�QC�Yd������z���[��n�_(��z$��
a��~@Ծ�Є-ÄW��2����CǕ%�����ՙg��*�]Z[iUO�vZ�U˹�����SG���G����w��jg�����r�Y�[��qiW�g�-���Bh#`	2�x@=	�N�o�dBnb�/�f)PJ�h�~����U�*�A�\��$���o�=IĪ����R#w�o�O�v ,����Wi���_z{�B�d_|p6���#l���(�Y{mp0�)�ŊAU9�M���FN�n�M�#�k�)��� �iZ�bV�3�5� 8D+�iZ��Ǵ9�E� )�+ �*�;����F>��Y&q����2�wV��=��"�]K�O,�����(��qw�FF�(�F�ܽ���ټ��e���?Geى_��d�粻XkP�ќm�H��P7��oZ��u�\�[��s��Xm~Qa|N�V�{�ojDj�e��ɩ��b�i����ȝ�WZ�c�.^S�N�6$�Æ!�?��\}wU��fb�:�Suw�T�p����W:H��,G��I�maO0�# 1,�j
d-�� D���z�8��p����ق��> ����%��"&Q�����A-?f�WU��:զ<=�.�$��a�L۾����ëYu���Uu�A��4��r<o��M�`�!���e0��$̰���
���`Vد�,)E���-�-k���׈��
��T&bE��'Q�{��!���0� ]����[Y�	����;�#����o�:u��A�b��1M����/,�	R)�U��v�2w.O�j���ߐ���<
7Bm�)�6�{��R����4��r�_$l���K�U��Y^a������4�l�t���[�-�b,?�V�"��&��y��Vm��(Mw*��b ��Ybt%�@��}�i2��.a��CZ��Uo�9a �%�]w��sN/�"�xz���"t8;������:B��[����)�k�F@�ﲈ�x&5���=]!ݖ��	ٙ�D3��J�o��x���ًMB���yۖ:��[��+>H�9�h!��c6�Ռ�CfE���j��%1��_˰��X,�w��g��p������M6.�	��SMWw�ݒ�b���te�e���{�h 9��S~��3��"+�Ơ��c#g�k�ݬ�����^��D�) ��%��<�3Iy�U·GT5�y� o]6.<P�<�X���Ya�*~��D����||O<�B ��ތOTn�nV&�t��2ا�!J�c'�Ňs�O~s�ڧ���
5��%�6IӠ}Z�N�hY�6D�f�-}? E<$����'R����1is��w"Us��� �?�4)�&�-?*�9���5��ҳ���*�|��䔡m3�mc9�����is���5G��φK'"0�h�qUiT�u	"�l�U���!����"��v���aE�'�o�G�
2J�3�n<�9��Z��(�jz��rV`�p��9�t����Y�>1s�=>�@��~"9h��-{�p$@��Ë��P���;5ǖ����(��z?"�4��"�w�w����
2�y�#y�$�KF���)��'����u������JeN�
��{��W��gU',d�OZDA-׃������X@�s>�pT�Ћ�?�]Ы����x���n$��v]أ˷Lg����04_�-�ª�t�^�'}�����b����
��0m+�/\�(���ä�}���^_ !���`�g�*��{\�Ck>���r�4������X�mո��Pn�5O�{�T���a��"���A�E�����; �J�k?4t`�_�jx�����zDs��}�XE$>��ͯ�0r��o���@Etq*@�3�C}�(���8�/}Պ��੸�}������w:M�c�SfU8�� �����l2�{��C�� �5�p^�XV��T�y)'|���8r�����e�,�	�����*<��|Yٺa�Vd\}��Z)q��Ẏ<�諴���[ixf�8G��rǱ2:ے9��� Y]"�+cӴ����M&�^+��Tcƃ]�R�2�Nȧ��<��
�x^y��[y�ԍ���@�)��?@�����e��?���#Ml-����V<�<�rS��pϭ�+�S���n��0��9�:��cc©/ׯ@���+yxɬ��J(�X�F�<�f���% ��qT�K�q�ܚcZݳ�@?��M���jέ`�Z-6����߽���v͜D�Vڅ�Y���t��������.j����b:���L`��"��R�%$Ř3��F�^�INf�a$9qnN$��93:}�i<d
�� �V��5i0!V?�%���D�r'1�Qʖ�{��i�`�l�"oǇ��
�ء��E�t��¥`1�TK��D���zu�
�s;%�j{���T�-4��eq�W*�vP��#���T&�(���88�;A�m�J�X*�Gnw���<���j��υ�T\N��=��UB��� yg�>k(9��P۸A��(
v�W`�!��Ք�V�I3@gǄ�GF�u ��J|�_99*]�Y}�ɫ�E�s%�C����=�#�~�=�8�z���奪&�:�!�	�^M�;��f���D���b�^��Ak�-�sy.I3i򵂺�:���T�(<A�Jw���\������
Ѕ����M嫴���&�&a�u�]P�1�8V��-)e�ql�H�H��*�/^`('L����s��f��nD�qϭ����"?(����GW����%}]mC�HB�ޭ�A �m�W� �$���A""�X����Q�5[p2la��\�ɇ�G���7�,�O�Y)�1;	t������<��Ȣo� |2�Yk�=˻�=޺��<!�l���vh�iZV?� `c]�9�D�;WZtmGߚ%�oM5���3���:^S@5E�fz���`.E�p���w�u�k��ԇ��Ҹ�ф��4$H���t���� h�M�!=�b�g�Q�ӟ�_���-�Hȱ��j���ǡq�(z�SÁ"b�*f��Hy�~�m���Hl9�Հ���8~���,RHڜKA&�}��fY�ٯ�/���I'j(U��0�"���u04r������u��8�x�q���"����UHh����ƨ #�n*�Y���%���1[ġt?�Mq��s���EtW�.je���y�*7_l�"�a�ݩ��(�V���̍3��*:ҥ���-�0&H���-m��D|%f���S%�G1J.-JW@;A��ٙ�	�(�pg�O�7��-����-�]ˋ��DD�y���s��?`_鿄x�X�d�Nޮ�SO앹�4Qa=��<�;>�,��4��-[͆ZZ�b>���G�ϐ4 HNks�~쮠�v���O=ހO�N,�,���1L���9"���]����%��@D���{�A�U;���C_w������~6zm\Bj���gg��j�*~k86�$M�->p�{ �5R�
�0*2�s��)uh�� �a"�k����-nY�~��}ّ�!��S>D��٠�]+���\ōGtSfR��w�)[����s3^Fo�կj���U�����^�	��8�G m?��Թ���ߩ6y��Jv��VIrr��(�C"��DBr)�G(:��!�-���W��y���44�&?Y���)�n$��6�&����լD��>R�޹���{��U�kb�?_u���@��Oۨ5����0���\���q�E�G�fuU���\��h���yY������!��*~4:eH�#0�~;�*|4�N#=W�?��5�)�/�׽�[�}I��@�~yd�n�B�(�u��MR�	��S�W��%��%i���}_௧��mTj1Q�(�J�Դ� k�����WF�Fz����d�uy��a���F�L�>�S��=4�J)�h�Qʊx��c�Yo\]�����:ռ��!޶A͉�Ҁ<��+�'P
ݝ��u�y>�%!���_G#ܚךM�xhe�I6�y�h���=vS�h����ļ�0���4�^r=����
`]X����c1i�g6���d�1�"�:?� �4�.$�X�l��+�H>j(��xZf��/$\�:7�l�V�j�q���H��0�k��9-wO��ƈW>:��/%r�zg5J�2�BZDCO���N���N�41��{�*ˤMt֓��p_H#�����,_��@^~I�&�H�k7����]�N���JH_���.i����̴tp�� =�6?�N���k�*NN�#�gR'dbi�ȣ��7�J$+syd:���sE{iH^7"q.��ݳ�g�!E$��Ȉ� :���BgPo��(�<t(Aډ*�d�K�Md�j��=EJP�s�͚����l���$_�'��i��������'"��b̲�~�&�)���QP��-�(���6�� �E?YB��|��̜�k(ҙ�ۮ�]Dc_l�A%I�zO���r/YAh!��Ӫ!���"$�d�F��oJr*?j���9�{�e+��SX�UF���!D�/����P&��n�mp
(KYrS�"��igd��T��W�>+�xg��Nߨ?E>�k��v�]�*C��Z�^~�(,\�.���j�T�����?�e�N�F��4��?�u�=�+��C��J�6��K�'Dgo�\��D@ھ�VQ
1��\������@�0��\�d�T�N�NOը_{V2[�xC�2��I�����X��ǹ3���<��H2	�E�ac�s���E>mߖL��g	��8�*�g,�-R$����q+/0����"��W�qy�tt����IɾGhc��A��-Y�[�?�m�)lu�@ϣ�d7^�vW}(#gj�fOV/�� �MM�È�-�@�Ҽ���^(�!�[xK�|SD.���"Sg�
�QgiRӹ����7�Q&HK$��f�Ï��'�NJm2uiD"=�0U)�K���[N=C�X܁��T^J�}g�Kn�x��Շv����ׁ�-W�)�Я��,g�存�3�Oϓ�����(G�AQDQ�m7=I��9�V���lRrX<��9C�\��� �o�ꞖT��O|�����kԓ�	�5y�W�mi,FU���ZW���h��|h��F��>���Egp���J�dtc�����&��	�Z��F�K�Ti* �r`��39 �f�([P�.�Dl���z$��>�{t|4��a�Jvl���oR8 �� �c�����	�%xm
t���:�^���Y=:Q��)� ���<q��8eg�ܳ�	n?��?:%I�r�<&B��a2�K�k��Ӆ�3���bX#}˒�<����[S���Ўˏ�ww��6w��R��M��O��뫌����L��w�w�빚�:�6��O�3��V#m�ÒQH�܊e������~bj��L^nn��-�z��� ş��l����Sؿ�����6�aI[d��'���In��-�8�����_�p�Dl..�;�m߮@	�b�gٲKu���� I��)�l���d�R��C�2 RB/�mƪ"4���c}_�hu�Aexœ�|O�2�_U�!�߸��X�I]V�CoNY��XC��U~��B��fv�������i/|
�.�&BG#�j�v�\�iّYXۍ��ꁴ�0��:V��8����ޚ�ϥU��}���"V@U��j�f�����d]NZ�%,�1@��ݥ����x�9����_e��Jou���"Jܻ�b�g�c�~���F��5z��#-1����g@Y���@cMh�ncXR�(��I��c��[o}�܌>�N�&��Ȝ�ò���/Sr7dA�Wͅ�0˯Oվ�\��+�^���T�wh��d�ǉ��*4�R�m3� ��rQ9�O��=��/~��w���-��h�<;-!�^̈'T�tu7nԣ	������b ��k s�v&�-E��
�t�^�3��te��3u����y��G��`����s��z���������$d�c�@zY~+�:�x�9���iv�V��J��ۡw;�3�ro6�W�̍��.^B_�L�,�������@��^f�(�U���NXTZ�GzXR�6�~f����n� b;���ӌ3����'�/ �>HOG��R~g���"�"�V�a#y�H�Ԩ���W�~� ���9�x�HX��uǀe����.��:>!U��m*Nvٛ푼o�!�ZX�a���;x��CC�04���� �u;\)� 6�
X��Y`e�I��j.2б�HˢG��b,�뽦�#�юx	ܔ�7M|��P�L9>��C���- ��"�R����U����lh{Q�l�?
̇�(ka�v�#@���'$������]K=F˶}�R'L�숋3��*h���	[v�	�Ѕ��"��Є��o
��*��𥰚���g]o@�x1sq�L�'|LVūq���mlB!3�8�;Ӎ�����T��=���~�e�,�R
�0�Ҹ<v+���$�~��U���6ʎ`�)C��柾	���8�|������*҃� �B0}�q���*3��xe��[���a�����r�8��9��UM�c�����z�4*n的m���k��&LDV��g��
ez!\I�W_��5ih��y����g��p��vl�U5��Ν�1�"�ʭ<sq l�O��*)�\O�*����S�ӯ�K]hc�U�VnI};}�U~G��	k.�{|���,]Z1�	�	�U���1����{Q��jt�"�j%�`���6:CN��c(�vT3ҿ���M==)�I&�8�5�j��ݤ�{i`!�����w;���C����7�
f�м��;����<� P�d�8s+TP�/���c��;�HH|;���t�6\��=*��\q�)����6X�/�u��ͪA�_�T��7����N"i������u�㜃>�#~t+�j�m?/D������TtwE��f����I�?Z�� �W��������6������bp�Y@����܍��1�I�\����ƊT~�`�|��� ��N\�YxCHl�k���B�����p�P-/�����ѰVP���B"�݉s6�(�Ix��G��h�Vȵ8��Z#}�e�'"7U�}���m���jٰ!Z�֦X�\�m���O����%Ñ�{J��_�,,��K08�lǍ�5�2{���auRf��2���}Fb��Oi�$�94��_D~m?۟�]��s�{ü
���|�]'l��n%˜�,�iJ�'��u��mv�����-*��V^Z�L=�R�g�M��t�>�ޒf�,������j9[��|���������k����'q�"�*i��*@���&�4��1�b����'&ŵ�@��#AZ�<�]�qn���KZ���q��+���%wz��٤i�Wg��{;�1V�-}zR��՜���p n����� �͊�L	&BX�#\�y47HN�q{��[��l��l�8j�b��E#N��r��O��^�?������s�LL����C�A��Z�5����U�X�4�Q��Dњ7�&_ۅ�9b֢C!����W���Cz�<n�i�$	����Df�A��ZwN�������{�2,�i���)
����.W9���E�4֏-���7���iX|�i�q�><�B�J.B"]9X��g8���*�1����҉ڭ e�V���(ؑ���V�	�i��m�^P<cؒ���<�JI����,��b���WBژ6-�e��:��W�"5�O�z�� �� �̚`���W�|S^~��G��u������Z�_}B�?9Q�f ��$����������6���f�� i��M��Z�e��MA�=�!�5{&����&=�gP�{�� μ��&B=! �"���Z(�pGF����m��s�l#�Z5�������eN�y��v#bWu�U4�˜��p��Uv8Ц��d�M�a�2���q����>�	�*�� �5����2`4���4b	�Z�z�A>���:��u��/��m��k�d��xT��1d�f+F��!��3�|n�70T���I�˷u�� ���ֻn��|g2>c�V�  �X�37�W����@@?P�I�4���!eR%�%���1�ݮ��|�_��J ��F�[=�XVȰsQ�����Tֻ눅���O-#yM/G�ΚW���h)<�TI��,��(�+hH�Ц�h�D[�5Y�]���eR��ǲ�"��'c&���#��j��cB��T�j,=i#�4�z�H�q:���[�֘��u����!���Y���Dŷ��~[�[�����[���:�\�����&�馯�pG�7}�J豅��u����zc&� U�����8���̧�l�T+}�*V����"��k�-�����z�%���~���H�QY\�bi�S��g(��c�	SSϊ�:K�LVͺ���x#i�:w��h������-x�Ӈ��H'�O�,0^�6���x�&.$��0Q������)B�r��9�!�]���@f|�뜷�ӷ�����d��r�yX19�zncI~�*����_#�Q��"�KL�q�K��5����N<�>��k*�i� 톺0� ��n�gDK�N��;0�K���G�s{��ں��C`C8�?�%]��_վO��m�C�G9�^�C�v��M�)~B��8}�Ч�W��Y\�-1�\t�)�,�:��/�Y��k;���FG���ʕ?���Y�SkA>z���T������Y���4��?�����_/t����x������=J�� ��i�J2�]�N#�_�.k� 1���%�M�2l���W�q���KQ�X���p�ܱ`s7�B�tf�I����B ������n���������TlB #��zE(�z�lc7��4c�xd�1�w�Lt� �ʗ���3�DP9x�aGsCc��|tNX�ܢޣ!�se(��b5I7�hܴN��K����I�X'0R�Wζ[�Y��|uV ��<n�.V'�� b| Lj�|����4�l�7�Q�81`���/�f��da�K���vU����B;��e���D�ʗCݢX���3�}��dO4������hN��GU��5��_)p���[S���e�֟�k������y"1�Y|۞���03��j�<�_���]�\y�zcG��x9���aĐ�)������=���(Ӣ��3!L1�?t�(��b���؉GRb�> �Q�bв�� #1�m����u'��a�p�l�/�b��)�O͍��!�
���	�\e)I0t�~�
�Nъ��d~��ъ��&,J�V�L��q:MĆ9\kv?��2�}��;	��?u��������t|�ia8 s����a�^��Ht����|�,],��2�J%7åDHe!b:��6i$�}I'�JZ�w'�t�@�+&H�8������� m�˩㎫%��ǻ�$<���Ὥ25ġ�	L�1V/��5��a^BgZ�����K�M#��^���Tx�0���u;�W����(��8�����{�B��DB^(�(Ɇdk�f`K���g�>�sYL�3���lc[�Ȗ��nF�>'E�9�Ar��]H�U���=>h��j	U9Wk�ݼD�G��K�Mw�!��}�_:F�S�"����Vh6�8yuU�� �Y��T �����aF�;j������y<n�Q���hpaB�}U8������gަ&�� ���4�aN�5�lEy�7�9i�R��͢W�>�#��\�8��/q'�MMu7%�o��>(�;ᜐ9)�X�60h����)#Ec�����7�����FA��e��H���+^�7��D�j �7�K�b��Y��_>2�vjv�([O�L���f�Lבn�lK����.�vKҟ�6*~��j5]=$����3��qكJDz�L����M��t�Z�?G6�0�F��n�x�܄z���Ɵ�%�;en������h$�c�]tZ"����!MD&�J�!�E� ($������V�eR-7��(4�o̯7S&�)���^�K\4X���D��L��"�
������ <�0��<���k�{1�J����}�`fcI��m����Z�&�4S��Ԭ�Y����ם���K;��L[C��7@���3$�&��Z�q7�uh�t�D�ўMfn��ݖ�����W�h����=�b��aM�>x�)�]z=�������'b��K��P�9)i/�&�IN�h7�=bw�dI]�zE�SPjwp?�9M�찾
"J�T<(�"����!51��y[����O�!n�Sf��H}���{6��3���%��J&�	�O��*�q4<�i� aU ͕>p���_�����a���b���O�p��4"�ȡ r�7��W�(a�݋��]���l�mѷb�����<|bm�~��Ѐ΀�rohP��0��U6�u�W��2dϳ��֠�:�[�(�h#	K�zDPcu �jf�L鷽������-�	�!�r�奼�k��֜qwx��Ĕ�����+��<�8y`sA�_cUq��?��H�S����Т6���f��9"���ja��]ࠏ��Aa;�����o�j�+>Cv�Z��I/a���6�=�I���2�y0�ϱO��N	F�=U�T^s��+��<��=�Z�I�C����)��:�Zөg)���9mi�����JP}��N��̇���<����u�v�P��A��)��^����"��
J
)V�A4m�J"�+
,�+m�Ax��B8Г�]�1�G9�m�,Etk��$�yS��M"�Î����m[|Oiƹ�eҾ��%��J�rh��%�)r~�qj!²��nM�n�F�C���BV�6B�ﻷ���/�	�ݭ8� �Sp�.�أ�${^~���7.y!��U��b�5ܚ��-�#����C��q>�q�������̻�%�~]�'��2z�i��x�	 �=Wpԋ=p���	�̏�ʹ���sw���Px�@�s- �p:�����w�h��y@Ƌ��ճ�
��I�]�%u8�16tY1Oq`���A���<N�ӥت�����1�+�[e/F��?b�+��}�Ă����e�mS�v3���/#�'���{Ofp��_
��`z�����p���X:��V�礨�~�	�M�l��&�VhJ0�<Ћ�1�ӧ�q��(�E��F'E��b�s{񬖡]*�	O�W�R����������r�~^;��&�&w��c�7��f�:�gm��nexQ Ɓ/&1�P4ζ[OHFUqˋՍ�=�]Y�@~�JH���&�ِ�έ�-T�7�_Y��;/ʾ���ZJ\亠��(ڻ��i��� �Uf���Î�|z�M�[��1+���|����-zBa��(�q2� Q޺�ș��d�mg�����*?�Dv[���zՋaV;$��%{�.�֭MMn��ށL����4�s��k��ut���,�uG*©íąE�iFэ��l�ﳎ@e�:��Jɢ�������S;�@=o�f#��D�:��9���4ot���{���`�Wcg�\Z(��T�2qUB��!X�Oy�����6aҮ5HIh���x�E������u�X�;ď�-����8��GRB�\��iCN���b^�Y_���)�i7-���kK�C�^�<�6{��oR��G��c�z`G��'��pQ�)Y�+'��V�M�ױ1\B����6@o�^1���J+ �l�.��g�$\�#�>���Q�����M�`
���_c�L�d�e4<.� u4Ö~Qح��ҹI@������~|0�T*�WXj�v�������МoX�Jw��7�3UHe�����N�]��=���S���J�����z�JŖ_-O������>Y����JzQ��h���F�'�j)��g#d��}⫛�����u��mK�2!��Uhj�:�Y�p)���A�tʶd�k�~��¾	>m!� �G��TO:Q�����z0�T��BE�
	�ޚ��Q��kxx�����\�yp'�$!^�F���&#\�)<��E���2H��4P��Zy�*Qh~$�Fq=���'���#kx���n]ME�+ČR�̝gY�}I_��[9ʰ�o����
'<�as����+oB����屄�c�P�)�[8�N?�ĉ&�8RFE���k��)��e�y�Z� ���w�%L��M��&����n�8�B�AH� _����)6���6�9��"��A�H��&W�����v��8k�^0�o�g�=�X��E�N���Y�����n/b�	<��"Ӿ���@)ќ|;�R�vS��|��t�o�[:+'��0c6�� .a��!�Wh�IK��J��琙� h�G�+ȉAY�.����y��b�ͩ�e�z� ��6�~X�A+�G�vj���/�	8	�\&�J���׸��:
�a$�(�J�^bf|���G��x��oK�9p?��O�x;�O}��/�q���ZI�E9�@�L��)�9�r�j�� 1}��e���۟��{�#���b�l�;aХ_-ε�M
��*Nwi������X�B��A鑩r!�j��k��sH*�j#��}A�~��RP��?q�(-|�fHR*��=$g]&Z_���f�,����b���a!�7�"3�1E���_���5Z8��pF�"H�Q�)�(�P�A���~S���B����Q���.֖nȽ|�RK+1���tBJ��+zg��b�cQF(�4A찁t2Q����(��<�-�J�Q�q� �������]�_b�lRVO�B���'w�&���~���>���M�������$[��u�o�n#� �1�����n��$1�\�;� ����N&��^Jp���H��i��4��2��\�Bf���NVϔ��̱!�p`e'�����*Ř�T4�z�uVc#��
��Eg��Rf&�\��[s0#�L��s�'���m��V|qg� ��V-e0�$ڪ���9�H���b.m�!��e��laQ�%(/�WS����#���:/k ����j1WA{�dY��V`ՏTfiB��P>�S�5B3�Q���H��O2���u�R"=]�R�:3:�<�ʇ�{vՇ~���' p�{7B2ش��Mȷ@Z�3r�����k��(iS��pˑ����[�	J�f��tR[��������&���3�~kʃ�烺�d�!N�թZ|�{��c&0�����vG�	�4��q
;��ll�V�N�w{�ޮS�'��Y�m`&TqT�U��t���O�X�7hZ�>*�-n��a���GGS���w�*��!_k��;�&����FSeS��Q�����ܪ֗���*�����:�a��!׶F2r�m�EW��t&FO��ee��^*lL��܀��ؠF��U1�D���d�axf��x�����R�@&6 ^�ښڎ����y��zs����o��,+�]pêآ��^n���c3v�F_�%i��ɍ� 3��m3��igN���^^q迢sh	څ�9s=�+ݽn^�)�
f �:�%���e�U���K�=Ƌ�!� �O�����T�<��ݜzS����Nyԕ'�b�EzIa��2gb�Hk�V��5GT�� ��P��v];j�(��֭0�62�i_�&1���V5AXz}:țlx.�K8�"��H���t�T�- �B��z�s�	vex�Sf��6�J�Y찠~��`N�1��֪%�j(U�:�b�M�J�AS��Cձ��#Γ�zêoR��#$���;#�kUA�Ks �#z� ��v5
DR�N������yНS���;���0��UV�{UNq��?�u+�l������j|�>a�2��P�x��\e��=��]�i�ͩ7rl����sЎn?����[�:=���e>�w�G�֙X��P�Ͷ��Cam��sL�������}L�(�W�4%ޏ!�1W���&ՙ�M��y�F$��!���S��C�Wt���b �g9x!�h^�|��/��`ԪS�=p�i��8!� ��@�ΪF-�����32�>��jǻ�a8���wҨ�㥔�k�b��䣣X�*��~^F��+:xʞ�JI�Cd	���������������<�f4��J�W�x\Oc^�OK��t���O�%��7�ֺ�3���R�-�#� ᘴ��V\��5��_8��<5�r΃=y}�0MW�g}F�5�	��856���|m�*�����yU�+KNjĮ\�������VR��]OTt�!t_�|�|��z�ʧ�ZI�ƩH�j^�)�T�a���t�?��ju�E��1�n���u[wjl2��YUn"?�O5����A�1W$_�&��Q`S�}���%���!�_s�+I���ŏ�7�G[�Ri�ډ'�ZSڔ&��d���)�DC��=�2���J��|"U�����)0�=��3}��1.�>���2S�[�4�|���;��e'V�JU�ǐf�5>/���*1@���6�:m� pn���ь��j���"Ǹ��~��F驁�4y�h�]��*�f7�y�V�h �C��?M�����"㠃]HU�,ٝ.r4 h�.��;|��*�&�P[~���a�l���UH� nʛ�GE�����?���/	b��Y��&�`�~z�J�X%�@�L1�m!�v��b+��j�+*�7R�W��g�4-D������w_'����`�N��Y�x���t���K���g$]�j��N̝^_�Y!^n��ˮA���c1k�i���ޭ���,~�����6bdhK��K,n'�d勧�|24�|�g�J�R "��ޯ��-3��rZ�#�gtL+����W郗(}!�a�B��F���n�o�bd��FZtϗ�}���}���Ck�����S��x�7@�x�}�~�hҀM�}6@��'�%@�M��Ѿ�tTX�®n=��K���O��Rbوm�����)�>N��W���{���~��z���J����? L#Q�i��j��%s��J<��ǽ���%��TE�������#��X��|�U��쁯��0�d��7�4x4<��8)>�@��'wzƭ�bni�����?K(�#�H�ϲ�;�)H�o����-�{�D)_��*���zq��L�E��X��R��a%�1b��D,�я��ՐM_���eG��M[�.�����y�By2�%����Xp�8Nh��!_5�tE�-�"�'S��wv����"D����gۑ���L��Yt���slN���HUe�暎��ު���{��E2Эښ�9L���K�m/8Ԫ��H�2#̢���*�w�.�}�8�kf-�9Y�xq=����Ď�SU~ǾS<�a��O5��w���b.�A5K�
뙿��,�@+D���wPh�o�%�F������di�疔0�n$��^jI9�aOM߃eHzg�/xf�KիSU�_���`k�rWL��3��d�\�gB��#A��u�%w;���]MѸ��Dfc�󣜃� �$8����9}��Q�~CD�JJ�sm�Oa�F��8K�)���GIh��׷�,Վg�%t}�\xJg�]e�ԏ�A#�͊!>����@���yp��$ �����d��` �0�T�.x���2����h^Y��ASw���h����R�2Е��fg��^��}s6��_)���
��������Q���	V��E�@c~=-z2Zb{�Nz���p�϶<s�S�@��hީ�J�0�UCj�Mr��e�t�:N+W��^�R�e^Jn2���r�8�n��"�O�G?/4�9�VkY�R�w9|�W�W<�䆅qMM��|V����]�r�9c�^
��u�5���X���׌I5�i�@�+�37m�l$"��N)Pح,��19V
�����u������lv|Y�/>N_���.Y�������':� ���/���y�-��$�9t��s�2gޒ$�64sEw/]U8�O�*"ɍ�m�:"���kb���Z�x�I��D��k�ٸ��I�ZtdQ���r��
\*�;^3�<(P~�h�Z��ZE҅%rT�P���jj�1�M/ִ��
HۓPa��H�_f���wr�OB!j@�4éw�f���@ [^������V�
�<48�ܙ��SG.�{-U`���]�����#Fzciu2�NZ�o0���{(v�}K�e>C�e��d�O��p�4>�Ù����S�9,���5A�H:��P.i<���m��J�7�_�J�h���'�Br������}��XSjϮ+���Y<������d�����/�߁�92�jN��< º���yi��㚋g���rQD�J����,� J���3��{yM�R�W�\��H�>u��g5��A}֩	��Qe,h�W����qy��F��S �0MF���xKKp5^*��;!��
<v�ɍe[��YL[v�i�f�k]��q!'�%)X��c���Vo�f6�C����a���B,x�4,{�oń|��]/��i@�_i���9�z���l*�q�b	~�ՙ[͉���ri|?���a���b��%%��0�OBj�T��|a�>���4�J&a��]x��9uz�pQ�f���`�[��}\v�Ure ]D��n���� ��&HLϑb��a�u��5R�P�Z{rn��K�I�t�	X�t���,�J�{t�v,�l��Wrp7$�c�Ƃh���s.�Jp��a���Ẻ��0�<�@�Exc���W(/v�[��1tP0�Q�X_~kmR�T6_:[T�V(��-�Kl)��U���5��T��Hp�iu�g�;,Od�3
I�a�ՎI����1s2�vK��7Lg֦����O���APo��R�әꖮĦrc��ZE>�d��-�Ţ˚�K��q0���kUΉn�������hA%�̪�"f`���'���hW�A�I9���f���@��1�<��w�[�R^�]��毖�,{d1��3��aa ��Ev�<Ez9��p2�$�X7��4�XP�7�F��`�z1���f��'�\Za�>e�G�mv�C]�H$7a�R����z�����W:���!w�#ФN��;I�K2#U����|?�� ���A[�L�h����6qL���:���e�%����o{2��ya�{y]��G�,x�(�a �R�z�U����-�˯����Zz��c��`��ލ�����߄�Vp��5�!^�a�G�"�o��ƴz�Yqr�55��uG�j�x%�.Q��0\��̢;:r(FϪ�i�J8�@D�ti�QVL@�Xꇁ|u�v���-��X3� ]�#i�F>�ȁ
(�#a�ZT}������7]�hAݽ�t��>\L]�V�GN^<���*|�#�t,!j7���؄_����5�_|R����?��z��#}����Yas����ͽ�#	:�����)!-]n=�c���c�=ܯg�{����D�-d͡�pPug��Ǣ��x�Q�a���.�dhKG�_9_sC��x%s��+��/�s�o\Na�H���A�:����`�ojr��\I���.ʄ���,jt��� �{ڼ� r�H|2�">��:6
I#Λ�6�(��P��7�x%�RCW��[Yr�@I��q��'ꙴ3��`
��a��<�E�$�#���V	{c����+藀��K�r}�T쁵O(kF�W��ZU��4������;D�-zu��9]�M�q�ش�އ;������P�J=��k_�� ����� �՚AFX\��;�yL���<st����J`�h *8�y]J�P�/o�������i�O��4�b�z��&��#QgGi�_�%�#����~�Æ�W��@k6uV�ҋc��v���DU��7��䓘5Q3'W�t�� N�]QI7�ߨ�J��*-I��@r�X��{J����j�Z�i��j�� }r�����J{]�����_�/�GWF2+#wܢK������b������7H\�ǡ#�:l\p	u(ŵ��xӰw�[B�s���^|r�e�j8��_+���g�N��kG���/����j��Ǭ�;�r�`�p'q�p��I7�2��}r���L�̖��<�R���Ȑ�p��c˂S�+C����Ə�� ����^���7���L�|>����Դ/Ps��re4��|
NLb��� a�|���e]�}=WM��U�+��1Ѷ�|k8�����,�A��J0�si�H�5znt?�||���*!�9��W�i�Y|S�g\4�c�	�~�B=h�/��Uv�x�p�z� ��3#	l�0HM[�_��{92�	�S��B�|d�
�Z5��:�ݳ"��d�Y�������̸tp�ҖepSb�,a*p<K=�D���ae�Nj�B*>`ހq߀z7�� ^WQ��_]؁�|�	��T����0�b�b"�E��Q8󭀤T�X_�P8�N�ޗՉ>�S���.��m���jM|�]�uټ�oG�@&���W���.͜M�{��x�{�)�x�ӽĹВ2�t�@�m35v��4�ܘ*��z���1�^%�,^^�߁9���	�O�	EG��T�c�$�?���
���
#	��$kב�j����A�RA�Z6@���1X#��N@�z�ʳz��7ه��/���vjF,Q�|��q��Z�ѨP�n)o�/'/��7��&�~Gק�r�p,�>����FR� pm�Ry��I��J^�m�� ���i)�I����X�wmH핻| Mt�ԕy�����;OnO�h[��mp�� ��!�Xw2->�����	�����.��W=�4\�9�l'tC��R�.Au0��$�P��:@I�T�$�zTOMAu��}�M����]�M�KV��V1����8���v䁴�G�܅�{����0#>�=C@��j�E�)�X�z�"rÏr{6�y���P(�lc�_��I(VM��V3��*H�&Y��~Wj6�^����`i�Ԧ�@�ϓT�ϑ44�{�T\��N���V{�!^UR�8�}ɗ~<�"H�\0��`˄���2��U�%k�i�(u��q�yr�:ZR`�*���� ;5R�����'G��It@E�&Iy]S<>��cj�[O�`�\�����F�����6��RN��Ѝ�\�f>�En'���,����b�ä�qkK"G��v����  ����n�1Q��*��1-�y�X#�=��p��O��߲�>@�W��v7��2�]K
vOUE�6���/m���VҲ�;&�)f���Љ��Q-�� d�Gj��IB�d��ǧ �T@�Bd�f�����`�R�����(�!��}̃&��1<(�-�1DVD��q�?�q+W+\���l;�˰�C����<%�f��U� �i[؝��w�k:̅�7_j<�.�n��'�QQ��#��{�a��9P#<
�Ԛ��y�"ZLn���J0�L#�<[�r���Dl,�qQ[�(���h$�PT�&��_����H(�i4�-\�Vx�'�Lbg	��I�p�`_|� M�G�o��k�\mv��)���o�#[�#O��[hs�e+�/�6��R�Y}(N%�/���f�d>�I<�����1�e�p]� ��F�����&�e���v]: wۜa���ú^㼫!��۰ӝ�������-���y{�1��� A�ǅ��׵4��M ]�*�0vY�F�����t��9l�u�{���MоQ����0��Ж7��%g��/5P{�
_�Y�.* ��Hnu0!�J���?? x�y��F�N(�"�#��W��N_۾Af*�;[�9�I�����_�i��*���b�rG�UqL�7��Q
���t� ,1G�^h�a��O���q�ud�ݜ��51Pe�2���ҾXQD!"&�I�'}M`�g���?6��t����e�%�a�N2w�ш26l-��:�+���a*w�әM�/+uy���e�e����i=�S�-���,���W�ٟ(�}t�|��z��߀l#�eA�it�K[j��Ӧ�F�l2�9np���&�W>��t/$�Ǽ	Ym�QK�D��щ.g��!�U�"CDu)�K��gG�8�i�J�}kH�.�龎PͿMf�������K���a"͟����vWe�vG��ep�+�B~:���[8��E���o?�h��s�k��V�4:D�*���ٸ�2e�wҟfL�d���O��_�G
���<A�0��g!��I�� �[kv	0�$��;Q8�#Q4��" �7���<�e�"����i���ЋvmtH�;9������ g�4�տR��w�șa�Lx�b7���:MVv�_o���zHJC?+�ۿ�ݶ?�Y*��*����Ke%Ӑ��v�C���i�5��3J����nC������B���2ݫｐ������z9d�k����9Qo_�8�s%`��uA�:D��5��C��@�4A�u�7�HYS�0�-�a;0|EI-&���:�N��B[/l4��D�DV��zF��L�+�9H��
]�T�\KN	)���t�o>�z�S;���j*�G���h�­����)�3z�#�|C*��VI������G�/�w���ԯz��P�$Ý�dՐ�.�5�V'|-��G�?�ϫ�zE� ���ۇI��'=�GA�-s��ȎW�=i�a�槁,d��X���/Bڔ����`�85.�"c���zBmc �Ɇ��ƨu�a��[Q~�ap���~���`�i��A��YYr9��}Ӗ�fgd�nT��9�����%i&�n������qhd���P 8�����
�z�#���~��x����?;�$΁|�x�]t�>�<NF���h�z�I��$,g�l<��N�@d4�b��b�c1�o��ηz���hg�t2�r�"��ZY/�����-9g�i�3}u�� ��w��4SEQ��o{!�bǀ!�:T���)5wP�6�q#���c+Q�&�����wԵ6W��˶�en?�ᘣq�t;�y��/��5m]!c��!�E'Ha)y2����ϟ��!���`b�Og��/ND��̐f�춳sLHʣ��fel��PP��G<O�,ש(K1�+R�t*pP����a?Q�Q�r`��<W��J`k��@zFYj�}�Zy��X��ߜӕ��IR Gg&����V��!r��v斮R��X��!��&4g�q���
��A���$�O����~�΁��v�z|���m%��<� �x0�!1���%y��xp�0mb��:m��f����oN��=҇�-�=�P7��W��LE}�"bna��O?s&U�-���;m���f�>�7�7�5���Q}
�t�cu*��?i,_�j'�¯��R��|�c��j��j��C����S�QS�+���"����U0��?ZI��$�ڽ�j������홼'.�_���%cr*���6ћ�� �jχȴL�ڱ��Ѭ�!	� ����FӨ�����^ ��68�UW糯4�6 ���Y(-��۞�T�
b������&S��`/Sp�(<����*�'��B�ӑ��|5�7lE��f�<`�������M��uCXFw#䦺�T�R����gf5�(�P�e���t���N��l�'ݖ�[z��eZ^���}�f|ck"�$��oz7�>�fS�&�?��$�U�ThT09���>}k��"q�H�	)��vPw+O�r��2$�����[�d�Ҿ��,gaz���+��e�#Ċ0��c��|�p���FN}k�]�������I��w����p:�E��9�֠�+5*^���6�敷.z9"��;c�"�K:7X�Ś7*�I9C�>�w<�����إs���sgT����J�"���='�`Rk��dXTB|үJ���F���>�5�\V��w��>u�<9~;���v@��9T�Q�x�䃂s�]��+2�"Fxgvvϣn_T�Lq�/WV����X�ß�{f֑��H�r�Tr��I�YG��:U8��2��
Q�gGX�`���V^^�2P���U�EI��v=a�R����Y���(2�~�S,�W^ mڊSf�GY@�X�W�]��l��4��V.X�،��.���(FD�M@�y`�a�)��&����C��2
*���)��MdG{��E�=e�B6��w��3���/��T��� �V'/��|ҝn�đ�$!c�Q�Uǎ���m�q2itg���G���VHZ;�S�'a��!��ߨu%��$6}�{��	m.�	k6��������օƎ`���{����`���k���Ds&���?{����.�ݨ�13�^'����"o��%"�M����Q�4�}�<U���ړQjO�q �`_��;�E�M ����5"���|a�[��
�qIt�g8Z3X��N��>�I�<@�[9ڵZ�q!�X���<aq�{�-F�Ù�,�ǹh�L��:a�?���5�Qt�?eqOY$�p�ϩ�
M�Ժ��X:~�j��:r��גT�����_Z�_��GA������G��-Z��W�3X��y4�m�=,��=��4��e  hop�������"��4i�P���M�g�]�`N
}�Λ�F|���a�P�D���A���u)y�'Ee���?�$zM"���0F�K�c\?�ϗA�v��H&X��4��y�Њ�N�#M9�羷�����k��W��&Pv��`�q|���Hj�Q؝�LFA�洿Ki�� �d��6�8u�?����{x��6/q^�k�`�>`���\�����.�)'��E�*���T{�<�\���<V$1 ^��n=)�%���В=�D��GAcdC�� �N�E��?܎R�.-��
R�Ѵ^Nt� �0g"��Ey� �~>�����}�	��+��9G@�E�����A�^c4�κ-���X�(��e����\�T@dN
�*n��_ꭹy���k�b��_�V��Td�]�8��S:߷��B�a��@A�r��Sl�.>��:�J�8�Kd�6#��i8A=[���7� ����U�q���9�L�]��w���
fOJ�Ung��cB�Y!)2��ʀ��v<I����Ad��5u��	�ue���G'1��.�%����=Y���yTy}��p|�4[�̔G�>�6/�^4j%�E"�¯"z����L,DR��5I7V���;=D�n��R ��2l/Y�#�@4��3i^�h���G��W֨؆�{:����\M=ܳnA��q��Z��R���Xf�?���Rq�z��;�L��;���D�w�.1����d�|K�
N��j�j�}��yej�D���R`}�?"�m-X�h�d"�����т�9<������ݑ?,���߲*�a��{B6�F����}�*�Qt��-���ӠE�����"ǹ�/%J�M�}��pmj��w��\12T���3y���)�8����|��ӌ�[�q�	��N�m���L�f��T��|!�K�T5C�&��Ɛ�@�[��]���Z���G 6u�]G��>�Wb�:w����'���n47���_�s-� � ��z�����I�<|pԺa�̳5:�h�7�X�������l��4Έ�^��ɤu��ܛ�Δ���$��Y�ُG_�A��A3N��o���
��A�e~����Ǧ�k��<���0��O!��d
�d�B���B{_�����J�G|���[B?��XN�x q���Nf�ء��K��d����!UxP�Li��l�]C�n6*�\1w�oaL1�"����W�&�8r��/á.{5�YA0�k���k�����`T�p�wQ��24�/z�Z^��,��I���F�`>��a�&�WàV�/M��)�=/|q-���DD�޹4�������_n^4����X��O��ȔGY�w1�:��8wv�3�&Gٛ21�bH��\�Ա��������g��L�d��F�#�����0XKQn��\}�!�!F����:�(7�Uⴾ�3�y�v�܈�[�H����y�.ȴm`�:X0����_X��}�^ݞ�KD�����yV�����V��T�g���h.�'��/����1�P�+�A�܂g��l�*̛�đ�=���o��ٍ��j�����ٵ1\�]�,����#k�^!���i���TY�:�4ve����ҭVgS5��gs��Z�._�����\5��)LU�a1	; l�0�3�Q���4��ڟ��#.����@���?���h�|�Â�������-i�!��{n���2��U�B
q\E*͆[BG�3x�����H�y9N��%%1i6�̰N�������y\w�/���3���{�����}�E����蒈6<�MDØ���<{�
��	z7������+_���7q�2I�L�q�M�C��t6�Dy��Lmؗ��p> ������-�ĺp��J�����bO�omPհKt�$�>�D�^c!q�--*w�L���W3�0luqH�F�GI�=���W�W`�a�ݰ���6���W���[Nr����ـ�,6rC~z��G�-E�����A��zm*[�ؗURv���ƂO�' ��Mu �ڡ=��%���;�J��c[qWA��(7�ZĈ��mB�=��O.6�J�J7�E�ը�3e��d����G�$���\�i�k�w]8<�E?��7�^ xz-�I��O��3�E�O�A�[�i�� l�-LR�)f]���J����� ʢk�]�f�� �� ���>>Yek���#M}�>W�OL7�A{v:W��F]U�m��?��-������0^���^�2�
�
�^�\�|�]�xف\��H�7�B;����=��ib�S�}`߁�NDl�!�'N���@��TH���5��j�im���x3j������6��m�q6��i��-���Je�|COTO����oבf^�tn^J�O�!��,v��~���陈��ޒ��������B�t���jj��5m�5��:��]Y�=�ߎ~y��}F��[~@���:^��jb=�m	��h���j��3H�5������?.�T�c����0@X�ͬ�L��7�ph{���:�3�ܳ���U��r��șO��*dw- ��u;��Hr���{
m���Z���m�}߷�}^*GͶ���]�@Y�>@��y��[6y�pF�홼� |���n4U�=�`en�SM��V��������1�0���s�� ��T���陦	�_�]�C�Ͱ�Fe|�W�!����Ag}�GZ��]k�ﾯ"����ϊ��Y���{��R�c���w!�f8GѠ����Ӽ�=}�����4�7�D��S=��퉴FE��6#�|:׻�2�v /9n�,��|�_C�$���A�>�f�{�v`^��3LC�M�i�Mw1�>����j��m-�����
I�
O�6̉57��ܾ8��Ug�L�=Qv��Z�=�kq���*����n<�׀Na(��2ە�8����x)w�Mѝ�/D+N6u��N�
aaC�/��	�S�t������PTd��D���gR,�he�'��g�y�:�_|P�V�OV�f)���P�-'ĉ��b\�j�{��XZ�^,������L���a�Aȁ=�>_��[Pxb�։��Ыj=�}����	Y��L�2p�����b2� >���bT���p�,PP���v�G\B���1 �a60�5��{ZJod��4��>[m��2��"����I`���Z�B������8d
�p=���̙>��2� t�«;��yjWP�G}r���Q�o���ǯt�hD��i9(d�։�<8�ϗ�t�\��ߕf�iat�9����w-��)�rQX���˕�\��Pŀ�9|���H}.��؋*�����M��E�C;��,:�ˉd�&*�_��R�	)�b�NQB��@��SCo!�:���f��2\�#��TV�����Ʃ��x����x@�-���,�\K�.�g�>� s��fR:t��;��(�,��� H�`$+�{�MF��1��<y�B��K�u���=�s�Hl�:��,2"�.vz~�Lu�9\T���fy��×����V�پ"����OIw�T=Q8ЕS�(�5�IK�]	&f�o{꜕C�����*P����+/^�S��k�����(��1H�����U3�|�څ,�{H���3�p��"gn�T����M�塀��I��z���VR)�(�v�L�p�&Z�z�E��Z������85v�<ߩ^w�A6�Q3�Nk�Y~��'�)�.���٨`S=6����X�1�+�jr&���Y �;s�W� ���5g�����A����]�J�6�<B����W�4O��5s��{{�hV��5`W�1���M{�*V���4g�3)[��Hz� �%ͽX4/�|�2��tr�MI/��Ȯ)'�+�����XW A2w�@Pڤy����A�iEs�K�&g�:'³��B�qZ��;���+���L�ڮ���%����'u����{�}��&7c�t�4g����D�{���r�e��!s[�R:&摈U\�lސ��n�6*z��ө�(kp@�s��+�x����{�hYYݿS���r������R;������b֝��m>.^�������?���҆�����?L;�Rt�ʎ�`t��^�+ɸ�1/�f�a6Y<u?Zt4��b:n�i�ys�$�|i��d]�eA5Zu���N�J���#_������t�\O�	��U=���e*���s�0�Q�1_���Y�'�� di��XV�X��)�����~����	3�{CȺ>/����hw��w��rgb��2ѝ0[*�;ó|�� hI���M��Y�{r�n�Jx�1��E�G��:Q-n����En����T��ʼ�����-��ߢn�4�)C��Z��z����Ъ�~�Aǜ�dO�!��``z������Y�=�:i+/�*e�Vs�g���"�ԌD�ʫ�'��W��(�D�m�.�w��|.�`�q��.ܭ߸��nc���%�^������|��0p�,��Mre��cB��@ZQ��y��U�*��꺄Z#�mx_�%�p��b����h�f��I��)��5��q�;�5)S�\���ʨ8Ǹ�-�Z"c����f���$"��Lpᴈol����6�k��[|m��e��D�.�99�)J���͡�5-N�����7�.V9��b�h��{�Ip஬�#̀�}VG�+,E1YCm%(Y�è��Ҫ$b�z�+@ȣ+ㄧi{t�D?����2��BQ2��j���>���E���_��qt����o㦭�����o,O[����_W��5���f���n&Z#�J��k	�a&��(�/�?!�c	�����d�Z������d�%Mu����EN{_�=���v!_�,�4���Zs'��c�2������.������ �4�tF�&��C]�oOC:Ā�tV��GA��"�K�Цn�m��1��Ǽs�2А�&Ti(L�Bt#��Z�G\���H�r	�(�-o7����2)�,-��<_E	��"=�Gg�z>�C��T)��� �HYTl��������d���t�f�j�J�{�7��?n� ��`](�r_�)����}~a�;�4��ۨBL����+�I�3�eP֊BĀ�!���+9����q��KƁ}�]C�w�"$��� ��,��j�Qb�qu�t3��,�S�)��_όRQ<m���[��"��\�ouS�7h�e�X��@�	<�<5��0�{����%v���������λv�s�`p,�u�g��"� ��1��E�_#�
I>�8�+�3vk#U�Կ����1�	Ά�?	�]�fZ�H	��wlnǑ�YM�����1�Qo�EȀ���դ��+e%��ɤA�P  ��B�Y���q�?����v��7z�������}�/�3���5�r��o�����,�:y�W?�m��˩g�F��/x.�+<T���� ed�	�8mN�F�Ru=7���?ָ�@Jg�xJ�d�F�����,&�9ÄU�vXTk�_�<Y99"9m�����SEf���]0�l$Wݰxx�O���:�y�4��EƖZ����c79/�Q��p&��] �.�:�/!�ԟ�Ǜ�(�	Κ��jR_��%���+����jE:��ua?��	�$\�U� &&6��$�۔�����5R꿕��|R�(^�ϲ���ۭ��K��ˠ��)+��>I=��輻����`�o�(y�I�v�" M�5��X=8�Cnԧr��(�W(T���yQ���Hچ"��{nة��Ez���S7X�Gk����z�Sr��M�\���+�}��C���1�X�ׯy���˷�]�c���%�	���n+���'��^������0�`��!��,�p����k�ǡU[�9�kڳiqx$B>��~��Ԧ��2���@�=�����I�j�pa��N�V-�>�fFR�����g�`�����ű���3u?ନq�j?ڟ#A,�f,���%��z�1�B}e��w4��CE�a��t�S��<�A�>�������� *"��.�:���G��=�(��,Dg{N� Alq���sKuKT|�8BWp�ς�i�Xy����@l���e<��a,0h~Y��q)h0-+��rhǀW�8<�d�V2O�^h<MQ�V?���Ϝ�F#�[5أ���F"RG���I|To�q�u-Q�9�v˵�F���Ry
�<�xGt�HHT٦��q	f�C�R�V�Jw��H�hN,�ܓewB�ClA�Ɛ���j�R�Zd�Gؿ�g1���E��̝'m���&"#��tv倃�� W��^��y���ey_Q�P#Uj����y�!1�ls�(��y�B$H,���=I��`�W��S�S}�9�=<G9zo�.+
�v�o���T�y�U٩Vz2��'.6��N ����'�	U�%�P�AyC̰�w���3��G��r���v���,"�]o��B��ջy�=3��"s%RI�x�:���q<aC)}n��a�v��E8��bn�.F�B�p�pz:bj��Hq������s>�{�*���ܖ��z3�'���.�=�h�]��V�_�ڽj�L9J������EK:%��W�I��8�;H��n�а����NS-�b��5Ⳉ�+���k���f	yta{5�!R�u�K�+j��� #pp�oI��m���T���//ň��x� ����h:��YJe���g�[��ޥÖ�6�4t��=�Ƚ�X+�-�N�Eޅ��ǲ���;u�����{���Yy��+X��E�ƥ[���A����#R[(�տvE�)Zq��������{|a�s��#e�H��]I���+��5CW
������-�"� �z��E,xve�E�l��r|���l���>��W��`}�N��Of��)���Jļ���G��q� dC�l��o ٝ'��dU��:R��Q-�������fX>F��JnMb�*rl���9�m��hM������w��-�RFq6f�[���<���ͮ��B���-����=6�r��6�Ƴ�Q,�1IG����aD�A���	�b�u�����&9}��B��jМ�'�N��p'g��<wv�!�My-[�(5�e�(o�4���4ƪzK��j�2����+�j��'ByX6ҧ��7U�*M�$�bg6��(H��igL��~�[џ�x{Dq�'����xi*��QI��ў)�M��5�8R1�"Ҥ�.b`�lG��R��`h�0W��b5Ȫ�۪�Z��gH����D���ӱ[1#�a����&�5�g�9�O�M"����=�� �f���
�j�ǉ�����g����|�
�q-=oe�`:I~��!��&\�V �\A�Z�B���9�-?��'߿
�@d+�G��Mq����E�Ϩ�9��|��{��)��xlO����Ld��FE��j����ݐUT����MȚ�D��d�M�U�;k��o(h�;���Du+�Ʒ��6����J�5�Z�a���ķ5w�s��9F�3��B�~���T�2�4[:-���k��I�֤e��Yص�_|0�J��k�����$	3��2?\�m@����wC�bЩ Z�S��|$?�F6	�h����$Ե;xP�_�0êҌo<�������@{Y9��(����k���@,M���EU�^@���F�v��`,���18׵��W�NE$�� �!��\�\n��"�����rrD�@h���^�����S+T+�����M ������`�td�//�y�x�r�[p����@&=�e����i]D��m��<^���x!#Գ�`+^X+��I�L�C��嬊A(�B���b�~`R����7ٶ��nE�`S��g�CAgs��(Ֆ/�䩣̓��8�^�&hp���J䊟O��(�]���KAǨdoN���]�����"UT��:"��cNu��tZ ٵ������������ ��}b�ʝ|Т�n���D
:�DYcl����@o��Bň�K�\;��؍�]K�7~��i�.�s��Oe������������0EDAct�%T�M��Mu#Ƭ�$PW4DzΧ�""�4b��t\�+�'�S9�/X.�7B�Bߐ��}JW���q]�a#;��lڪ�eus��n�L�SA�1�)�7ᆖ��T��e{'�Ayʕ�p�Df7; sG��3��z|�Y�R"�>�B{���Z��e�+�����2:��D5�pZ��ˉ�,��=G�~�:У�>�%AO��IߐZ��6�*AXi:�i`E�L]�K��F������ῡ�iŏ�8yy��*F�t��#d|��_X�7e��:���e����_������ڟq,O
@k�kW�U���o��,
�yQ�y~wЧ��	�|�m
���")d�9���?n��L^��ZqR��8O�-Be��p2��ь��ޱ�R���S�ք���E�Aޮy�0����F^hq���T�c�bw��v����f_	�7�p]X�RV�L{�oO"RCf�O�/tu��Jn.G�,'}\��P���	�P��d	D_��-TI:�r���'Ɏ3�%�(h��C2�M���u�f��+~K�QI�{��z�q�Xm1
�O��w*�Sţ�n�Cj�̋�i���FfKkfH���M���c�~����7�,���@�s9�.�7�dn'�ΔA��z�#���#%�:��u�Z�r�E�e��qr��t�׮�qK��*���W�����q��,��*"_�7�Џd�D�>�/�麴NFĖ��T���n޾�l�w�Y���#2Ѳ�]��x�n�E�z��qdZ;�׉32�ˤ���O�_�9q�o"Ca��S�Pk�OW�ܐ�4���R)ݩ�fL���Z��x���,�r;�v���3-����W�7a��@E/��ߨ[F��u^a��U�duK�FP܌J�O���	�搰Q�T�fѓ���"+p�*������v�����8M�P��SN��d���x�����NGޚyp��uu��A��y9����ّ��.�;2ዲTU����l��"=~J���ŮQ���}�us��^��'����V��CϸҷNbRT���	�I���B�1����^��9��-lM�˘�|�����J3S�T������DG�;�܋]�O�O��u�K��gVd�lj��mP�Ӥz��C�ʝ����b����9��@����F�8�I8p�6�#��jF�=����\�6����!�)άǙ�1zz���Mjk�%>`4ge5S� 8�O�2�s���7�D���	�5tAvi��9t�d�5�nu��mw��G�O�P�m��A/�U�uW{��#j�4Fs^=�UƐ��<��-*[|X"%�E:�o�lEh�	����T���W�d��cP�)|I��������eV��lc��|���v?��.'�ms��C��4��T�}%�7cW!}�����giu�C�%��E6�+R�$|	�3%C���>A��M2|.(m����F�vI��^?⾣�`"�"����(�x�0a����؊�f���ZP��A���nֱ?��?�O��k���_��t*-gڿ�L��#���A�O��bR;@�,���Zl2�37�|�H������6��؟��ھRq��~i�:*��Ż'e4w�(vˋ��䘽��f�qm�#�#3�ψ5V�Z�u�7���07�Θ������a�}h�T��0�K�`0�MV%�Ӱ�� _��>�Ǹ_@ˉ
�w�y珎�^g�?*k��U��˝r��&�<�=��|�=��p:YH��f���.q�Z���p�oO.�A�yW}��s]���ԕ
y��_�ƒT	]�c�3L¬���}
�;@�eOh��]�@6,?��/2����n u�V�Qմ/݊s��z��'V �&�d�6����]�@Y �u�� ���CA��C�U�5���[�Zģ���_A��Q�W�o�ȋ�4��x�h�;rW�-P
b�3a	�IVu��OSq���'�ıfG���-Fǆ��+��C�fQ�~J�������u�xL��m�<V�D;R�ʞ��+M���r�e-���cTn��à<xg��4��z��,��3\�{���)����.d�����mw�! Y]�m�F]m����X�_�F�1Z�WC��&�NE{	�Q=sc��E{�k"����"ie(�2�"rEH�u$�3��'vBB)��Ov�]K���H���l��y����p��=JT�}�8P����>x
l�Y
�q�lV�W��i���c�����3ͻ�"�.>=P�1�"��ryiҬ���;g�;Ȯ��Nz�W@&F�@l(�#��R9�Zص�r�>�u4Ě�sN7`eUqFI�Χ(1m��R��?�IxQ�ny����v�I-�V�b����ݧ;ySM�ҙ���K7�T���*��'`���^�i`^��V;��r$�R����临J �DI �%�F����RV땝��G�\kO�mL�p�:)[pAj59a �
g�|�YC<��y�p������%`�t�(NꤐGh�vXw�K�\��8v��`�v+T��Fu���e�k�'7��}�Z��ZT��@�n��G�ͰR��8��.�c�i��1��Z�����d��� �c����A�e��K���Eں*�oHJ�&_�O�y$��jT3���m��R�(����mW�Wr��wt5�� � l��pY,��>�\v�7����e�Q1��j|Kn�b@{�INo���?�Y�ܮWFv)�Ұ;��\l�2�j�������R=���D3�k_��BAtXj[�֕	⃫�,O~fg3i�>w�����J����W|�vpW���C�''R7���B�r���U��e�>e���(�(vT������H��;��'5H������<&E�!�#��wX���E�E��5o�M�X��� ��V�é�U����U�s����N�bk��w����V2�Y2���{���>/<cx��e��-�����<�@��Ր�r�u�8c�WZc��O>��#��࿚<X����eA9jY���j.�#�8"�GbZ\+;�(ɛ�{��:�տv�F�󽁴	o$�!x�骭�"�/ ��j��A��/�p2R��I
��h�ӠM��	��䝈P`�����U<�WM����V�ԥ�P��10� )�59<�!5c���!�G=�P��ji�v��+�ft��u�dQ4���:{G����E0�lo�zk�R��/p]�P/��r�v!',� �S�:>ef���Ѐz���3�Nc���Ya���	8LPa/� Fw8vqv���5v��t��y<I�A��k�jhv�4�Z�t��g��R?��sH��Re����)��zTK����m.4�YEQ��jK��Ы2˖��yJpJ�T8$������ l�s�3� .V���ߖ��1̧g�A�������݇:RXN�f��Q���A�;���eNt����@ݥ:li@����r���ؗda��E�o��ժ���.	��z�"EhF�,w�b�}�q��r�O�:�H�u{�(x���'ꂝk"[�D�x�_�-�/���_��ZP�9�pr���b�D Ck�dd�*0���Gg��ʈ1OY����p+���wߚl+ӈ��fd,����Zu^�Ϟ����c�����^)֍�bn��.�,���	g�yg�FX��s�C��j�C�Mη� ��1��5��\60h ���![s�/��S�{��ڣ�&5m�Z�}�	��}*?���o,٧�R�����&�B����X#���@t!�<�Y&�Ͽ�Z�|℘���O|�`��s��<���p���(P�y������3W?T�p�Ӌ�5�U�=Q��r壭)�5!�� s �kI�HE�����oL~b������T�q�J��ձ'�>ii�db��9�v���*�X������)X���2�q	�`���ռ'�/�,w�WLȤ�o�g���׊���%U�8DY^��g�h\���hc]���tǥ]7�BN�E�y�v�+�'@/�q�ic`�bv��ҫkir_��a��Ru�	��^���.f8��l�)�N�)fl'7i���S��fY5�}�͜z�_��8����D8(Ϭ��{������m���㮪S���sG��r�ܸ����*�����aʹ��q�ނ T����q(�v�/m�YY�k�q{��o�ۗ���F¯D�,��-���^U�����9$��#2<�=9:3_���ʣ�\�)@�>�����P0�;WV�w�=�
N�?�_���-��75��z�c�+��$��0��^\�W3�E�����?���R�3o������)���B)af&5�礆aɒ��$�C>�a!����^'���yh������m����Rx��T�7�W#�bH�/V�ы�[:[�;�ޒ�E��a@K:	6��_P�Z�SG���d�m��ْф�r��rWW�&���+^�r��X:T��f9\��"�2�선�����SIŕ mq]wL�B�m�/`�l��} 	�軋�[$�X��Vx���Q�o����6�>�QR@���Ɵ9*/�I;��ǂh�¶���2c��݀��;U>:noZ$o?�
S-i����u�~vǫ{���x�mG��<�:�69܏�ϙp�K>�Hj�v"����g�e�}n�SXם�x����g�k��(�,�Kԫ��4�>Uٯ���}�W��Æ�2�"�Ū�����Q�j��l(�GśUXrZ$.@��*M0+Z�&����`�9{����֮'�F���c�Nt<׮�*�l�@��Kg}�a4� �,�S��vH��!{G@�/�h�4Úf6�:tC�!)�&b�M�|^��$D'ĵ�z�!��8���"HJ�f�"��>S���~x
��t5���$0�dO,�Ɣs4u��Z(m���(�b�9�_��ܽ450Ģ���`�p?qo5�cGE��,[(y�3�o����V]y�I 5	Z����NɮM�AP��ܽ�0V� �H�{]���j8�[�Ȣ�vŪ��"���[k��RԆ@2T��Am�Y�-�1�-����B���aߪ��I���d�c����r�;���,^�e3�2{�D�!�C�9.���b��Ed�i�sE��/ ����ۡ�]r�p��:��Ng����1��&�j� �$XEK3M�wL7e���u�\U�ZE�V�d�~X��dg�a_H���
!�$,�����-�x�	������̺��p���������������5�=j'&#�?&K�*u^ܡ-���[�͞�O�NV'N}<������CY[�L�+�X?�C�;�ܵ��R�m��r�{oY��?<)X�����_x�����l�7�����ӛ���vf �F?w�}i��9V�Jg��`3�ޚ��b���!l���%��c�%�О�����G�q���SX1��?zք�+���7�0�j9h�|.k;^?�D$��sF��rцl;��,m��.ѩTv�X�1m}� AQ�8��M�q��o�4�:�<�#&�bo��#���Tl��,>W�2Ӥ�z���|֞wwe���o)�{1���R��I#�E?(7l�ꛊv"`�UIWz��CD�q�cf?��\�b�9���)S�#�����em�V���Q�Q&J�E��P��nc�y�/��^�xVΫA4�˨E�����E�"}Ѩ�d)4�^��'���]0�7�Z���'����� t}��dc��p�C����V��!�z�`uX�m�H�(�ݝN�zg(�p6��=�  E���;^��1F�7�q���Ga|i ����-�����!�!��#��8�
��,�1ǻ�#9�Ro�^qv���!�_&z�_9������?���L�Cu�U�mO�®��~������ejb���(�F��h8;.�k�����4�� ZC�73����yh�WlF��(<MW�[�m�!<���,bR��L�X��3@�ژԹ�NJ��m���Qb���Hb8)^4UY-�~�P��,��t	��5�e%�ӽ�R�RQ��sk=�E�-��F�}�� �&��m��>�LR�+f�v�p�m
�Vt�/pШ��1A���#I��=��X7}߽<z�[�X��J���4J��`w��VьA�ߖ:+c6�i���Z#�c�۾��:<�"$X2����Z�z��p����,&MR��/<ۼ��BOr�)��(���,��b	�� +&�"��&�i,5�T���%�g�f�YD�R�gkɁ��.�.4���KG}XT�ޭ��غ۪/'��rF���5m*y馉�8)�)dY�L�#��t��[0��x:�1�M��;�2Rߏ�-�-�L�.���&�C��K��S;~\Ŭ��*?��{�H�Q��� *�Qk7�y�j��^/�����peg92:��%��KA*k��t���݃�J42kv��������N����ȑ0����sS�2�#j������&4�'D�|nj[��YU� �zNe�WݤtH��>C��B�f:���jD����9V�V%	`ʖl���H�h�����yec�-G��^�K���`�:�*�=`�N���g*!�.W�+�2	 �x�@,�P��Ł�8!}�%x~I���{�^���� jU%O����m�}PX=�_DWP�NX�]��c��:$�m�	t��EB����kƨ�����1R�H�R���*W���Vo����
�AOa7.�H����q�;f��v���U�_��vWD"K�����UI��\9]ž�m<��Sx��Z%������>�͵��Y�l-��Aʐ�`�P��Kn22B�ʓ]&S�������,�6�2�;�*WrZ1��I��17s��"ǘ�h�/9w]�������6�g{���_����5CS�>��x���ƌ�X��_��TP�26)/���U�'��� �뽡���ں�Hɘ����-�3�����h�&B,1b����9�n�
�VkWL��x�3>G��ۅ7w�g�
a�&z�A.���M�z�m���:9�U�ߥ��_���A9������57����э��zO�H���YL�z{�i3��[N�I��YE��V���I"��=YPo���U�䶈9P����n���u�}1$]|E)��m�hb}9j��;'43�	�C��s�ON���k����#t��-�#t���~�,B�+�V(�p�~����t;���W�A=Fq�_۝�+�&[b�>.0�@l����ہߙ��۵��S�s'9$���^_C,�o� ��q���!��3�\�.Dқ����;$�˹�g-K�zEn���� 1�D�����E~��#���]���en�۠}0�u��`؄;�I��-y����w�@a�����ʐ�f�	�;��+%'	�7X��^HK�{��@�U��M��$�6����C,��#l�d�Al+}k~�:�d���c&��^i$'.�W:atTs�ً��,]>���?̋^�gIE�R��`P3�X,��NL�mF�K���m~*{���g�i�a_�WE���a�\+�m��R�R�n{7����4!q��6tf=oz8lxX����{�h��g�9�C�U[G�*9<S��"Qd���Z������0C�ӿ삆��� m���T�z/��1�FƯ�n%�͐���cp��md^�z�B������ޏjj��Q��aD�m�J\#~��#��؁7&��Դe|h�a������`��W�d��(�J�����4�)��I���T�M���g��r����ׅ���Ip-E�qmi�h�L:�^ޛ�"�鬌�1<E�t� ��le;g�]ڏ��W!���P�4�G]c�������٘"�*�i�X��V�9�N��Vy��AJq�$š�::':G^PSk,,�!�w��eiS�o0�aƉb&��~��s��_bg�����^��b�f���X#-�`�'��A�����a���hh,�!@�p���R�I�jmƥ��$`\�;Os"e0�e%�Y�'��뎟bVpnx�I��4��ӕ8�9��%��3�̀�Y���e�+kr��B�)��|�����Q1���� K �|U���FDu���x��[��k=G,�)��2F<:s&'�>=K�Yq7���8��BXByoG&� �ԼVX���_Nf���l��%Ր�Z`W����͆ڂG]V�%<~7!�K�Q��}$�)�N�(���v��r��v��}�fj�~\��^���E�5��d9�Ǡ����
vx����E�p��W�$!���.WTZ�(���Z;>�E�x�.-�ip�~����┠.�zsd �c����/�*X��k�<#����#&�Q�Yi�}����8���;r�W��D��-��*7�)��ƾ�YZ�t5�h���T�3��lx���1�±p�aJ�3�Y˺-Ě�-`
pj��i�ݑ=�)�] ͛��L�c�F]Z�bXv�hs=�� fGW��5�gw�FQm���A^~f�����Ly�x;l+�,f>H�rI�U� �br����#�׬��xNHa���;7T�b���"�5������^�	Y�w�I��"���{�����-5�Z��^�"'��<W���6ԥ��q�I��P�Z�.Am�Kv�|�ɼ)Iqq;_�L�׆��Q�q�6�"Ya٢�?j����$�A>d F�K�v�;��9�����Ȼ����G� �ǚ����v�#Ǆ���v6t�P��-����}��gw��a�7�NI�LU@�7c��Ĥ�RCDq�$,��0��
4�������a��4�5���VZG��x�=�!��'	���m��/�����h��C{����QU>v��ۤ`��9Ѩ�(����C�G�z4��TI�
���U}�CQZ%��đt/~ӎyἚ��}F�y�g��)�\s�w��4D�t�u��#@�S�sS+"jR7�7��������M�<����G��7L�HU���l.�Lz�@��n�K���{ą"���V	������"��Ej|X��,6��OB�IXt���@���g��,�5�>��Mc�T�|�SUfP����(K$�����T�>��fI�SUzY��{̚nw�cf���>(�U��;T@e�K��(x����?�vC�,qBY�)��Կ��K��n0eïO	g�I��R\�AMo���e}�U\��D�d�ی�a�կ! ����<:=�}��+��E���'>NZ���3̠��j|*���ӎQ�+;��9����m���I�`$VY�ZWT�!ߌ�߳�������݃"i�ʮ06�#�z���=�p:/�$ʬky%c�,pғt ��<�o.!D�u�D��4�����I�:YY#b`��ӰS6V��Y2�חB�@"H�R��$j�2Ꞁ2m������,�1Ϳ	���,t�~jR@" p����D.�I{�G�|c7v����)��*=�X���4 ��]���V��G��A�5��~X���(�@٘Ƹs��of���CU����<g�Fo�m�:�,9\_e��4h��_�%c|#�LjW� <�gA5"�f��B�� ��Dv�@��2�~� .լwJ�٤�tA����_2sT�a��;��<ݕ���l��B#`.��!�"�vn�� �0��h%⫚+��e��@��L�4#8Y��t�Hԇ��Px���6�(c�����k>��IH��Z������@'7�Yz�X3�R���u�na^��`��ߩ���� r���|x���N�q��/]F�:(�s2�C�f�ϱ@	��u���ה�m���K�����g��w���*�Ih��.�� ،$ ����q2�Y8J�Է�fh��Z�-�>�Z֋��6�����7���ಉ?��p���*�{vcT�B�탑1f�|wȇ�cd}P�\���f����5)��O�Ǵ�"�䠥䫲[)����'N�*�{�v_[���Ym�.UK�DA����bOO%�/t�]J�MG��n	㽌�����T[��#�a��AV����/~3�U����-�aé6w3G�"�&h<c�S����}�vwD�h6��R��uH��jKٟ7��j��=/n�Y��Z��y�]i�^i:�z[�W�]=w�ndl!K_�hKT����z�!?���ه'LE�r�!.�FżXB�(ׁ�
P���Nˣ �d9�>��Ç�ZY� /��u��~�g�#��=;���lLW]�Y��	�D��'	��Qq�gia6�B�:��d��Q����EQ�E��$L��<�N���� �Ց��H�TS��n�&�#X�H-!q��]g ���#����c6k��r�Sc{R[0����"��/zG%��8��.�\_Ij����>q�nIҋ�Ň*'�{d>O�e�-M�C����䈒��(��OJ����P�f�2��� ?Eq�S��*�!�d��ﱓ%�a�T�W.{+��Ԥi脮�0��wm"d>؄"���G=�  h���ذ�F��9W����^�є���_�@�\���o��Bd�<��@�n"�%o�q�y�TG
�H��o�^�P�lTZ���U{���_��)�.PGv��5:��o"'����肃���:���V8D��bhVb�$�iW���si��d��Os[��js."H����U��3��������-l�:U}�ěFe!�����=�Y"@/
��)p^�i��)�����B�^'d-+&pV��SQ.*�֓����#�x�x=t?��>�	|�ĉ�
�>�5���������eَ�� ��T(�Ǽ{��tamS����>5g�2�����V���J�zG.����|mT��m�$����'!CZMQ��gФ����O�������XB���ȏF�1�����k>E^�݊Q: %P��g���VuD����S�� |������u�K 	��U�²i�A$��3�V��Ao��e���p^@����;�a�G��7E�O�<��M8.
��M��ʃ@����UÞ���gu�K��;�^)�GnF� P4j���]Z�=!
�}]��@M�X-�<ʡy3�����OA?�q�X=�k @��Hѡ�Fm�q$�&�~c��:�#f\h����C�u7ZI����)�������1
��i��T�����v��s�P����xgQ��̢�/�Ls��4���h.h���"�Xp|���I�w��{D����aVb�FZ�dM��������V��i'���@�Ε�Ga�(��e�[y�2�X��S��?�?
�3�&h�n��8Bnig%Vߗ�Ym�睦��R���T.��d4���KN�bW.�z�8T+�ٓʃ%p���c�:f*�$n\q^SF���C/vJ`��?�E�o�8�l���afJ�&�n��T�&�����a��@�#��v�bK�T�Ѭ��D]\?y��l��K��Y~���~���X'ǂ�1i(ӏ��D���L�s6��I�/��*�c%dq�̌Y�٨�����0�䳡�'<����l�;S/3��~�DCl`$�y�G�� Θj6Փ��
�j,;�5���W��	D\��x���N�6L��`���/�����?�~��f�`I]%�cH�v�m�*�$��!�:�xE�nzn���[v3L�l���,,@o�
��R��K�qƱ���9�����I%�W~�4E=��m{vq6��K�P�L�g�Ni�ņ���,��_��r�/�Yr�̔�gK�SM��4%���p����K�$�j4�X�F���zxk���/�o�7Y�^~��ť3���ܤq�|有X$���sdj��pSYY��:�=�(�"{.+�����}Q/�蹅�>7��=�P�	L���5�^LdV� mb���t�~~�����������3B�<@s��oC�o��D����""� ���47]1��z���^����z�.�$��6:%�N����X�B=7vMz�{�2G�(v�&F�����<�5kxH[<��":��(�Da�	�Ԇό. g�j�ǛLŨ�y4A�M�F�ɘ	�Ƭ���%��ش���Ϋn�8�oY��f�@D�Jn�Viݎ@��=�u��C"��m��2�����}�C�r���?~�V3����h�8��@p�{?*Y6��\�Q��aa�Y�[bro���X�L�U����5��r��d��[�O��d���f�[�cb��'$ڷ���K�0x��������Rڽ@P�AǪ�A�$ ��7+Y�CE����F�v$l9>E�>��^*��7�:��]=�K�tv亖���O���l�1�bU�N�fg���M���>}�>����E�gH��n�@Z��R�rAGu�C����tK���]��%��/$����a�1�D�������$���~�U0@�h��� 9Q�0�F�S��<۝��>�G�$s'9!�7���P��	�k��/�0+�������B�>�^tWΧ��¨��q&������tM��b�
��v��n��ulIA1�"���&A�ݩ�[P���y5c���E�>㣐k��wCr�7,�{�(b����3LH�~`�X�細h�1��.^�q���2�dE�5�bt��m>��~g�>����C��n�u���8(^�=��U~߈�D�EE�`��'~�Ѽ��m��¥�t�fM1[�$��-���1�}�K2�}�Ou�i�>��^|�ؕM���$wٮ8�<[g,h�ц�-�7�[OY6I;Eꗭ�͵�%��2G�x��W�&�s)GIm�3!�x��eFMO"C���
�Ľҋ���$z��U�V�lZR�Q�6/��Ҩ�z���]?�R*��d��c��ZF�衪��V�є�8s������P�^�{K�
1u7mT;t�%UХ�,Dl]z˳�t�+�*I��-�mk���:��@2���$�fА�:�r�|��ێ$?�	[��[�_[%I��98���F`�q4J��ą:�ke&%��ۊ�/ ��~��~:+,�[(�ΏG㜕�z�,(I\�p~1����%����#xxg��9妄Yp���6̚[o�ۙ�|;��S�qU)����2��q��;Ϝ5��+��sCV�˫�je� Af� ����g�^M9
hN���v���6����X����.�I��%E����|�]Vo�#�;,W#��1��m�.�+zx�O%�jR#��,m��G�� W>	�k�
ӟ�k�5$6�����@��8�