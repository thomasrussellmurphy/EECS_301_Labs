��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv �|�
����)���R0j��3I[���Q*������[�X��D"ԏ6d��{�0I���}@�J��1�^������W�Ex�i���)w�kN�n^����o1�B�1�����|��ȕ��,�3�[OU��F�- �[�� �o!������*�?>��i��3������#�P}k�1���ٻ��>\�t�Ʋ:&���/��C�o�%�q:��o��G��$Q�m��8�r��,����E��@�I�V�k���A�.�T��Tv�)�~�a��y�I��5�#�tK��=�Y:}��2�t�:H�Q��(�Z:����Γ��2mË�Ӎ�T{�/n��3Ң��o�2=�7�����w���`�����pcWSK��lfI7 �A�֠(���į�$n<�F���JT�������O�l���>�|��d�v�wo��_7
eSI{3Ch�M?6�1k�{Z��u����W��S��&A��(�ba��h���	��ߎ��(��V]�Vk�E��)��.�X���-!H=���9�F�V�9w�i�P?r����zȐ,e��+����)�qh��ܪ��4�[/J2t�WM�B
6�A��{��QU�Ŵ����~5M^%��w�$���2��9h��?��p���Vy3An�#�lK��z�e��xz�x�b&kM�2�����-�]��	V��v�,i�W�%�ƾ�&ϬcR���WK�X�|�B�;�e�3�$Tj^V�y�u��!�q3y��V�.�����vM��T@P���3sJͷmb�"-�Go�#7�]Q��~<��x2��9
�x6��G������Z)�����/�5�M���!�����u	u��@�Ą����&�Ă�	��7)��g�o�bu�k��m������S��i ]�_H!�ս�]�:V�gc��n�?�`�;��1�>/8g_����-K�>J�[<Ք��DIÁF�S66�Z�}�B?�O�%|��0�F��b�h��4���g�B�@~���[Q4��쥄T�x�רʹD�=�Q_fB��QE������,�^蓖�ƾ3Mb�H2�����Y�9�5���5l<0Nh�� Y��;���6ɮ���c�%�4��84+�:b���Rdg��}�oڙ�iy?hc��1���o�T�� ��Xma]0�b=yo˔6�y;#����b)��O.W[��b�"�h{������YJ��(����骓�d�����C��>���Yڌ���d�w�v㹝2�tr}q#�f�-��Vpy��Ǝ �I��/�U�QO}��z��YW�JD��N���
��p?ʔ��ސv�n���'�"��H����:����h�h������+[Y2�����,���g@*MsR7���l����i���}7Χq	0�v�W����0����
��E=��.��v F��V�R�T�7Qmp�R"�UPOr�)��3"�'�}�!�z��Q�q� o枷f��a�������̵J�����Ѹ3IGՒ�1����1��Qm��9~k+�3I�i^� M�f{醛��*_dw�-|�~��H���i�����8	�%�<o2�ܿ,��4�=!�
8�T�����+��^tRQ@������0�H���l�s^���M�r�Ve��27�wu8�[���>���[�$i�)Cs�9;�#�ρ[�����짙� b���l���Dsס!T�DM1�(�#��cy��7u�ٗ����4��'�7j�b���p�[���4q��s�����Bk<��-���T'S�i7KR��	�������ӃV�T��NF��j~�iא���ꑴ}��f��g���-�L%�7l�Jpۅ�s��\U�󇲣�� ����H�Y�U�߶X��6��*�' ,� �U$���i�C�t�xN�+/������O� ����}��=���Q|" <��	_d�E�INs#V��쎊XS�٧�U<���П��1,;t���Q99g�<6D��e�=�l�́��; H�wQ��EZ��G����T�oh�5W�.U�v����Fx���(#e��^0�@�f�u*{W�ֺ�i�2��������1<�v�G���<*���,�a�x�?->I$�����!@�Kqd�M�=pVr��b8�mS��X\>�Z�X�t?.fE����m�ʺh$���U6�ky3=i b5W�dp�]�H԰���k�I|e�t�e�B����uU�L:���]���/�����+��v۲�����5�:J��6�p�=��4��iV�+�Ve� ��{�����)���HC��D#c��O�洁T�\���hA�{7+|��s�@�VL�T|����UFH��5z	�舙��7u���\Hۏ8�Q�92���X�`t�k��n�X����&���	�o�l����U��P��ӵ�0s̀sa}����E�`�in�2W+*��笈�廫&�-��x�������z
<y���|��}��?�Q�`�ĥ�@��{/�M��ǈ{�E��iK��[Od���?<�f��{��u������oy +�F��"9Yd��(!��
���c�c6���q>yS��Q,|@T�~��p���-�X�g����:1ݢe�R���B�����RG���_�|Z�nIsj]������ݵ]+��jFG�R%ɮ��L;��PyHŠ�}���͓�mF��4UM7�gV7�*���qi�n3^�/M!�v"� ��a�I"=m�QJ��וa �w'��qѵ^V��T�lKG�g0������	������ҒRC��T����2OȕO��0Gti�v��-��R�=��V�aT^t�+��P���r�hiH���[�b+'�j��3q�s��p�
�__���6�<���ڦ�1资`�b��*|GA�q�c�d����͜������HfT^����SB����{b�ǫB�i�#މ�%��V4*~s�`�H`��:O��R?�[�|�]�$�?�-�2H�!����A�qq�K�U����>虭��q��΅�݄u���S
o�v�G��WKYC>�G���A��L:�v>,�4�����p!�G:�Aa8_��~�Hl�wN#���^��3�DW�[z��l���^Fɦfǯ
Q	�)�B|	F��Ւ6�&te�Ԋ&^26�1Nt��Ǭ"��6��/(�9m.�&�?�rJ�!f���b�˦��$�ʬ����Ƿ�B��"���+8HI�l���ѡ�뢲a���E��4R��w,�zRx,��˖c��F���꒥�]Q�\㰅����&]l�\�=Fn�\gϻS5��.2�_��Eͥ���"�Ya��=ema/'%9��oW������X��&��0�έ��5٬�D	���5R��5�D�x�6 Q�XO�� �<�~�I���0��;�E�PY,��C	�65�nQp��� ̠�ͬ��t7�	 d�&�_л���r���R��E��Y���ͺ�?���5`��{EC&obi��$��%Ձjk;�zp�X��_0�Mn9�C��X�������V��2�1P�ؕ�9�5�>�:���� �H�G"�w0�)���Ι���'�ɠ�@�;ki�c�/�S���1�s�ӡW�rkY�M0-����M���^/�#�IV�p��3���}�9\+4[)�)2�˚���6q�bcے HǨbFT�G���ij�i�ֆ��a�9�a�c]gj֮�~�G��O�z���ӫV��Ӧ��E�"18]���T�q3�^�X�ᎉ��+"0ʵB�W��N�/B�/��J���׭'5^���.�g��2gɵa��	������vl�P[q��J�)"}.a1�����i�)�Fy|j�e"X(n�������	��C�g69`�
#R�!4N�û�Kn��>@yLa�[��˓=����Bհp��h6��a\�����W�����cF`�HV�!�a��c7m�����P-~\� o�g5mS��1t#�1��*S7�0�6׉�����IN�=��_2�H�7�0e�]ə8${r��zbߍk�8�=T�A���-�2�}�TG�)H�}�>�Ͳ���:a�9��2�y0���oߑcC��r������n,R���_l;�m ��1�g6\�+�ԔGI:����R�YK�e�%�)y[��#��s�ĉB�l�#�����Y!e�p���c�m���j��"0d����2R�U{��5�G��o'�	Û�n��ZrZi*)I1�!�ԚUK�����w}nF@ dҋZJ` �_��k�QT�熖��gr��*p�D�uh���Ϣ2��>[��}'���xt�Q��w���L)Cw��Ѕ�׹zQ���2݌ń@���@�S�~���������a=���=��L�wG�$��7êR�1����^:���=���*�FW_#�|2���1`�q��b� �B����?��4�ƳQ@�YR(ŀr�LJI����Bk��EI�;m �50�Dt��h�������yP������X���X���E�<Cu�l\*��|?�a�^(�rO�@p{��E��Ts��p�����zR�H��v�k��6�K�����,l���4����֗�(/	f����>�
)ښҴ�9P�4����z(G/)�_����*�v�mܠ#��l�nn�"9VS���6W��/�b�w��<���4�t��Ep�3�f�nC� ��^(� ��%w��w9�J�z7
/󹘞�P�[h�;����r�qd�}��A�P1_��n��[�Ւ7p����)	�~��&��0nD���Ւ!����2�k���b���R�%2A�ķ=�)Av�dQ�Oy��@I�ρl	PW������P}��Ҽ�.�
|E씺^k��>Εů�"�`q�n�9�m�=!�0mO������ܱ ���r�1qc0Kj��
D��xz]���v�6�=4��#.�A1mP\���T8��{�<����ݝa��"�\nx�M�u'^����E���.lb�Ld�w�vEU��
� ��nC�`Ӊ���\�݌�Ʌ�6X�2$l@7�#�"���B�Ar�O�M��{K =�򑐪�x~T�n%�te��D�+5.�7���Ϻn���(\Xc=?�c��l��X���F�pP��9o�n��&z��3��fx�bו������g���S��ީ��3<IЬ����
[\ �n��X�ǝ_y��d�~��C=)!�<iK�����uo��^i7a溜w��w������+;��f0) ����ҡɉ!��]e�Q���'��@�iFX��� ��8n��,�@C^)�wr:2w�*����Ꙑ��Ц������y:�$ �^
]a3�x�*��y����<�t^�H�<��i�G{V>�/S_$(���#2��s9�Ӽ��f��>����1�|٫��. �"�{3���q�>0j���`�&í-h��g�<�d���k矧{�G|;��� ^Z_�k2fC����[UIA�S������BY�T����j���/>��Wt<��8���@�lVh���d99��㛬�#z��	H�e�r����7���Im
��T$��C%�ݖ	>1Vg��UEv|]?�s�����oc��5�鍥e�ƗC@F�����3xȎ87��av]�A��R��PJ�-�~ǚg��t��=R�{
R���s�r��#k�7���Z?P�=�� ��g�$]dح��ivp����+��Mv%��u�����`UǄ׺=R ���kX�����c�)On���߅���b�a��	����AbSE����@GE�p"��6������r\����<��.($U�$����7��='�<�%���/��q�v�ё�c�ٮW��xA�baS�5I�v�$�{���L�b�IQP��K�y����Ve�^�����xv����Z3U��+sf��MJ�e������g��Ҭ�n%&��Tb2�a��R=t$n�s9Nn֊���ws�XJ��g�\C��=�-]ךi�T��1�F�d4��w���-�ݶ�ܥd~a� k�˷h��<�鬂
���Є6�� ��XdX'����߭%����syq[{��&�Q|��-͚��d^�Lm�C�柢w6X<O��ƅ4C[ssoޮ�'�ؕ}���Z�V�n��=΃k�z������Om��C��]9�����ٖ8E�+y�1SQ��&�ć��XY}e�+�j24�`,/��  1g"Y��ڷ.��}\�X[ͩEה�1�_]�܆�h������\F,�~�ʜ"��eL�T��Xʗv�Nv�A�2#bƨH�@ȚTwMB�Q�匆��X���}�B�������B��_Õe����Jg�W�)#��!x�Y�k��?hZ���N�Ԋ��a'��3*�v6�1�$����^&�R
�*e�dF��W?BS���CR���m�gG�_��|��9��|"e�M���˨�
���!�k��0�1��)ۄ�I��(��PF�#xG5T-�nC�e��BTDD<W����z�rt�ضF��m
>~1%���sl?5�Z~������no���P�0��5l�D\ҁ���	�졵^!D^������B�tF��uX�R�����:^�<1[Č[�I������`hF>)����Iu�j?�xb�H!7�w��� �T]���M%��%����')2��!��'c"7��rF)�/=�����Z�<�.֝�}� ��_��E~	-me9xE{;�D�a_�N������%��\Rp�J�r�ߖ���tvgo_���s,������������)�J�9��}���Y�2���p��YN<z��C�$��� ��ͲTh7P�mG��JH����y��K*=�w�&�ΒA �Ʋ&2��*6���5�\�&��ܮEՎ-�R�I�P�m��"�7��sD�RC$�V�����A�f���k7*�y���*��0w��(e�{
N�Q�g�����7�h�&����+tƔ�h�:k�_��V*��l�'�s')�m��}��P9G���������̥�-�#�(Tw\NIP8	��q�����2(Y���Q¤�{t����	�(����c��ұk�P3j��5�[}��w٥f6d.K9���lM]���}>�D�3#(��0TP*�2/=>+;ۗZ̔�-��6Z`�D��L�Ua3^����OC�[����+-�o��Fs�����Ǯ�.�fN�OW(��|�>9�]"L�[\��2�)AJ�.�m.�"dH����`��X��`Fw⊷*='��L��C畇����4�������,d�g;�G�N��gnwb�7(E�Fx�_����\�B�l�h��%�%�6bR��P^S�uBw?�;*��Wm&�`>�_�X�TI��p�:
b�� ��%q�eB}C@�S��x䣆�B��S]Ycq|G�XCQ�E5�6C��"��Sm�CVR��,�y_u#�����-����:7��w/��\���n�I�1����m�}�h/��0ۈ��t�z��{[���7
T�6}�l,���k`�5\,[43�kRa�I��AzC#'V��;��,ܢV!i�VTOw`��Z�����\�z{]�4!���w��m�x�y7���5�E��fTd '�ʷ�� ��Q��ɞ����L||���%k�Q҆��܀�	s��t��M,���.���Y���p�"�1��33�fzH	5,E��+ie�9A�)�����&PS߱��-�e���3�ߛ�3�(]X��v�J�8�E<R<h�쎜X��yC�I��5�K�֓��W�7��h����K�br��L�����)��tn�Ikl����m#�u�c�[3��l�N�;|���RB�sM1DbKe*;�Q��$��8ܛX΃��2ġ��������<��	�՛��������}��q�׫a&��t�
�}߾��7oH���H�h@��/�]�v�Un"s��^�12�E(q"3:-���N^�{�M�� �i�V�9R�-�dLj`�#������V3u��DK�A�خ�A6�~j4pv�~{uSO=@����"mEC��!HD�b,�N2b>��'���Py�EAs�`P$݅¹"�ܡ�|�������|,�Ҽ+],:&*�f>metЇ�R`�1�כLJ_��
`|�j�Z�i���g2�s�j�:y�Oc�\�z�"��2$�������.�6Rk�B�}�\�!�Ϡ!7Z���{ܚ!|�¶�0������ժD�b	��?Q.B!�CHt/X=�0�����I��*�	K{�F)V�d.����٧�g��Ô�:s񞧣������ţ���R�U	��ϲef��YM�Ӟ����]�1u��$�s��ph����$G���n[��,C��$Ef�%�l(���'�g�`ax#5wL��� �_˔�k_"����xx��|Tt`K/����G�b��~�pi՝mp)��C�}���c�g{-�1��2�O�vs>�1qZHo�#Y���u���@�YU�G �
��d�|�3� oP�%X���"xbV�$�CUe�;5����$Cd��.#�=:_ڧIL7��L��!�$q��BH���˃@D��%e��/u��V�zG��AC�q���=�@O>1j:\g����Q�3�\�a\��� u��/f�9`e���3Q�G��H�T�+��s��e���}�� 8��S��j�{�q��B�c华�K
�7M�`�C �炍!�XY��9���?�7�ҖEƬ
��K%툳�s�E��]�_�&��w�:[���h80��eRXT"�-�<��G��7��g]�j��.�4:��Qv �=�O	�~y�����-���X��S��W������#�_�'�Ą6o�p�-1�`	��}#�fcE��×�C���|�r@m�c%���+!�K�ǹk@�^��R��W����@���Yܣ��%���N��#�PTf��.3��8}ZzE����M<����A#�b�ٞ@�2G��	��U�Slb�T�aX;��kL:̬2x)�r{�ttA�y(ߐ�N�a�&
�m?�)�(a)3�q���T�7.��J��%�6��4@�����]�r�O�L�ç��W/+���\��N�����K�0� b��$Q��K�}�ۢ	�T���5�1fj풤��\���xg&�vu=}	yji��M�7u@��?B�Jҥż7:|ـ��Ne�����H�쵽"�Z���>y�,���`5gu*����J��M��ׯ�A!GQ�����0�!���;�yz2,z-�$I��7�ISX�sj�ċ�3]ȶ�\����~A�M�f':+pޅ��9�;S?�wv ��7h�B˻!:>[����4�������|VfnH�9�;e�6k(
i�+b����4V1ۏ8$8}A�m���L@���_��My�O�5�'��U�~����Oצg��w�PuP�t�V;�<�Ђyդ.T2x)s��4���@��dܓ���lU����~��4AbE����G�����wǆ:g�5�p�!�#U`���lz�FP���T��P��?���p�y~���)�<g��sP�州Ao����f���J�18��vܺ�鞍�D���i�2�//�CTK�� �6Q�����=}O ��OI�|�A1[k?�s��7M>1�;{�ܦ�?��m�� ��"�zrQ�Bɉh�V���uX���0�2�#��4��e ���`
��������p0AlF��}!��D5=��8�w��Bd�	a�n&���0�u�k������L����O�dar�	 ��Y�^G�8��a�C�eiT>���WCeϔڹ�ld$p�,��:��3�I̬[j�
B �ص���H�����h�y��y<����RJ��[�0�G|��$x��S�9�i�]L�g�]<,�$m��U�xH?8G��*w�}}z��QT��e�mVX';2o�pg;� ғs+Ю���!�Z3ɕ�L$s��֢�/�Н�$�'	eŶ��XO�����K���-W�|G�5L>]�D[ԍ��Q�����7�bF���8�����h��r���<��ֳ��$�/Y�?t`��Ԍ3�Ȗ���ߣ���	�P��::�6���.`���]Q�"�?;�#>|:+��G@�B�w�
�S�s��,��[M.ƽ��-�DJPH��d_`'z�L~��2ZP@*(�	��]1�b�^�D��7���:g��Vj{�{`��w.R6�3|Ne��ۋ��-�=�`Q聞�/o�>���~��������V������4���G(L9��"�;�����]�j���+�m6���RpBF�;�Q��s"+��C�C@[�{�f~����V JgE��N*�:��a'փd���(��;}�랂�-����mo7 )��ѕuW�C �ZYl!mM4�@`��8H���K;9���P�&���7I�$бm���	�ꯙ���	_lӶ�G ��Z]xn
V�	Y7��'g�7nf�J��d��ܲ�}""<M��R_�� ׀�K�I������Y	Y!���GDh�ck�͐�S!A�;���{k	MT�P��
.�}f��8Fw��+f3�r	�L�4ŧ7��J�@YWٜ��~݈��?r��y�?�)��c���4�Έ������
��P-��_���F�u,��