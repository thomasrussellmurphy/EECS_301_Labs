��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,��.��̡�+P�FuX��d-��N��$%�I߽7>wN����u�]��j��ܹ�Ucל�|�=í[~��k�5�P�ؐ��T�5�����#�p"&�l�z�Fr&b6��,���Fԟ�Z�_�X�;���93	�����Ǘ�M�~���٘�2�c�D��������f� 3łߥ:ա�;kv��ތ(�}��r�{|�Z�LP�����!�Y{������I��܊7Է^f�L5�:�	�͎������W&��b��wD���Jݎ�IK��et��1���Lt�:��6�Ui�;F�o��!b��\#�Z��k!�Y�#Ao��U.H����Ƈ'U������0JN�]�[�萙��5��!M��	��1چV��J�-K��b@B!cٛ���qH�и_����d~��UImW{�a2�:E梂�L{�\���<=�Q<n�4�?�.XC0���E�9G����z)Ð��Ku<י���b1�����AtI߄;qϲ��ܦ4.���9u3۰:[lۄ�P�Ĉ�b �n����xkKǴ����Q�n��E��Z��`Z����H��JG�1<(Y&�D!�k���2=?�YkUcW���4��\D�ŀ�2,�y�[*��W�#��N.��u�SXo�Or�����!o�4e�8� ���:/Pu��T����@��Ro����wd%��	=��ˈ�ֻv�H����&g3�IӫVo� 儞׮<H�ƞ�D��2��v�H&0��!��]����`��Mc~I_���ΆA�	-�,23Ż�%u�(��f��i_Cjז3čK���ǔY�)))�q֦[o�$��'���/c�t�܂��9��.T �.v
�7Y���c>|}�۷9�|�ď̳e��5��_���>��VH)�"�-~[x+>�n�TGeQѹ�o���L�=�45IV�#pq��A��u�ƆI*��syxfY�{���by�S1z�`*����<����Q��@�j�C^}^���y�s(-1�>�|�پ�N���A��H�mh��D0�����~���y+{�[pX��K�����0�g���I�`�o���9�Bz������BS%����=$5g���E�:lC6c(���)EL�W����&g}`�@L�8*�I�o`��Pc�������K��O��<Ie��Ό���g�9c3���FGrT^��ל(m���S~j�F�k�Ot��!M2����<��S�Ot[���	�I�3g���]�k���]x�Ȯ��H�0bc��9\B�*�1M��	��I�'\\9�3���&Yuk����(pCx��+FZ�7D �R[b�z;2���	xa�䥙K{���i�S���\RL�~�$t�ð�H@+�>�_���� �Z*-���c#X��{�Q�ȓ*�,�𕯗qF���n��J�t�<VI�����6�.4dl�q�Q�$WY����}�E�$S�VʛI���!1h+����~�X��;�RI���EP�%��6b��0�k!��yS=j���M���8��f�.���{�6nk6b[��hoʺ�^��B��j�,|1 }�B��p Ȃg`��jܑ"�?��Ɯ�yw�r`��c��������g
3kq&���M����{�Gm8���uH.����J
�%ؘw�|y&�Q���냦���7�o�`,!D�y�z�ߟݰr2�j�K��ў!�#�GH�y$_>CEkJ�Yk'Ec\b��Дs��I?�]�~
��� �%��6���H�J������%����x'�^,�y&tP����mF�H�!Kx���[��A*-Bq�V��'���Ƕ��l4^����P%˖y6g��(���S�8���Xq_�k��~�_�(N~'��u|��_`|��KG;��d�n�K��g+�@Q�q�!V0�I���B�%�{^�H_���P�[Q���@,��X.o��0�����W/���6��Y�N�V������3^�>�������U�$N�5��5��1.3�i`m���}W:�RݖC���m!T�nj�ǶnB�L�}�6'�(���#�$��d�<-���Y>�y��<�&���k%��8�ZY���[�է��zխ��X�N�f2^<w�PFob�s��s1�޳��k{�oq����I;�be�)�{�x�c��o�vڪܮ�{f'��������n�%�N�Ȝ�n�{l���xk����w���\�bd����_�k�Ńܿla�R���ke��Yw���|�����)�"ȃ� W�h�w~t�iө�1�7�o�����E�� ��vݪ5 ��?��P��V�K��_�u5A�p���.���/�ao�p���rCl�QvФ=�����;'���5j�h�uޮ,���K&��t�����S��E���-*��>���S��K־�����O���QJP-��SmGyg)��lzB���x�T�ȋj^�?�N!E#���9����3U��W�y��-u<H��&{{Ǚ�x���H&2<+g���T%�E