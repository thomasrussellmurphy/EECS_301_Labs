��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv ^�n����w��M)x������8���#[� �M~���C+t��*t\il�(-�=�kej�'�2!�f.3��rw'nڧ)�*G���=hNa%�@��B �&jo�9Pdf�z�9W��@o�Q����
fY#؋��d��nk�l�%vZ��>v����:�"��#��{(�8YS�u~@	�L;��<��Ѻ�����@	��l�ں,�(vayfG�f���Sf��j?�<3�N��hz�ê�G�WQ= � I��\Ёw���G��,>x>7@қ�2�"e��jӕ�kO �����aW�Z�@}�A��KC�D���Np��e��|��H	����������;�p�Z�$��(q�(���Jp�[B|���R`g��I�gq�������[V�u�'�K*k{�����'fh
Dhps?m�����يx��F����{�w��A�.[@J8�"���P5eO��Aa��d�[��]����ljF3A��'�3:P�G)]j�O.�V��ǭ�ѫjz�^����i��I�"�*6M��=�L�d�P�.G��j	;�2����/sxi-/���%C5����z�	���y�p�e=(�Fh�2:5L�J���8f����=�?�N7;t�u�o=��� ��-�qj��NR5ݹm�OY�P��;����P���e��ԓ�w:E��c����yr���	<&T���:%xB�P8�^ �PH�-ֈ����=�w�D�q��bO|*=�-��I:�x����q�d�/�	������(�8Gk�hܵj�@��EQ��B�-�)��a��8�Ď�ž��YM�7ê��g*��u�F���`F4��B��uK����E��/�e�d�;�
���������Ej+bIT �o�<��.����*�S&�VP��k#��Kť~5B�h\E���7n�i�F3:yu���X.	���\��;���-HgJ9��mR�p	Oc�;Z����U��Z���tx[��D[.PW##Pw��_�r80mpf-݁w5Ť���T8{$B.%��}�1|����w�н`�:3�![)+�i%�`�sP_��a�C�֭D#�S�_[�O�\��1:W��@WbE��ʹ�'19�S�#�1�5�	��×靍ɧc��*�����sh$��m�k̖��oLZj��#���	z7��ba���� �ݫ�%��!E.d�`,Ӌ����/��.��4��/���b�P���@ZՌ^Y��|�<�#��D3�7�}x��aP��F�v�1�b$��\���fU���6H�4A��h-K�(� u��E[���H\���r'9��а4'�-sqy����O�	ǘ���Y�6i�W,�k�_E�ڂ1V:�⊵<�0�ņ����_^�S �3�)�� @5��6�J%N�:B��N�Q�֙�]�c)��֛b4��dnc���Rɶ�Q�:��4�`������l� 7_4�V#��ͩ�x��Ė@E���� �6��n��k��M������ˤd�qr�U;>���uɮ-[�B-0��u��7k/���=���m`����j�7�7Xc��/yQ�?���m~��F��n���C79�5%=�H!۱�����H��:�p��c��If}��;�U� �H�U9����/���ڤ���5��iG�Q$�lϯy_�qLX���Ǌ3�$�,/��T��)��\����\ȓĹ�	�t-���'�6���m�ԋ�c�ᤋ��֙���=�j�ƨ��όye���C$T�}�U�e5%r@�`�r�Dz�dwt�~Y^����P��]�S�R����x~�ujW�s}\G�sUa?�s�Y�Q�1� ����Uz~�E�(f�81�Z�<Jt/�,a:K����5Lb�>30o�t���>�_���T��6_�I��T��xkL@W����	�tK�R12�^�'X�p���8?ڃ�2��YHr2�]��:�pF��}z�V�NV��Z�ݐ5$��Ĥ���h����?cy�\�C$Ӆ���Ô]]�sp�V�n�V��q�C��jr5O��o��P��"1p����
�+�.��������:礯N���<��knyyeΰv�F1��]�!vT�����^m�/�����,�`�W�6��9$�:�o��:�,��MDS����2!��}fr�E�wW":�M8�Ytb�-����VE��qw����&rӑ��9�s�X�8�
* �:	�/[��8-���#{2kdw;��O�	�%�q��w~���(�ů�)%5��٢�M׽��d�\�n&�	�R�n#�ު)�=f�����G<^'FN4���)n��R����~7͜��II�cF��"���-�s=����&�Vf��x���'�#,�A��Ԑ,�{� �~��Q9�UP���$���ܲn[�|��!�g��]F��3��R��5](^�(&9��` ������&��
菪�;��UV���Q�)�Q.u�� ��e�P�-��l+��&#��{��/yB,��
����eA_W�v�����"�|�d�����+Q�!]�B$��=�o-���f&3���?�Nps���l��j/�?H����c,�U�I��1s�"@v�G��5&�B�g����.�Ͽ캎#����az�e��q���1���Nzl�${g}E/�ݲ6IG��C�ea_
��.�k$��?�%^,� za����7
�ok�a�Zfs�wI�E.;�y1��m�yQ��3u�XK��}��3��3J�@V��5�9���H�1���/�إ�e�<�ࡻ&��'�x�� qUH1V�[�QH<e�;d��Qx��`DJ�7*��t�R��c�#��#��r������
ʱBx+�L���������k:��byG�$�^�j���9*_��ph���^�[�8��}���A��;��~�F=WJϴ��n���21 �D�+��>7�o������(��>7hܚ���۴DR���Jc�x�P���A�t>p!~��1K��ֵ"��4��uv��k*px+FM�2����v����$�Y/i���r�duB򑧍���i�j�U��(�l��h�HA���~[���v�l^������.��x���t��dD��>I�m�c�x�7�ǋq�S}
<9n�{Y*���5`�6?��]t2b)B���y�P�mV�eڅ��!���X��P}�Sg&=���稉P�>r���� ���J+Š���"���FO�31���H&�g_u�p��T���!5�)j$�/�q��y�H:=��;�)�Nqf��<N�%�Qf�T���h=�.��ȳ
"�;y ����%�pCǯ�^Ǆe3�+�m ~���.���E9|�V�z+R�{�hf+��s�go�|5�.�LQ6 �54#�����"��Z�c�%նS<��Y40L�V���%:���~�JN��Μ����F��xh�.<݀�g��d=��@(�Z�ẟ&��hC-2�f�M}�S;�~6J5BCG�/�img���*JDly����S�y{�긇f�7�$�$&I���:�@�?P8��Զv ��S[�RW��g90I��k_�ƛ�ڞi����I�}�=�w�S�@�pϥg��Z5ah��L��gE:W�w�Gk��1�d�>$X�9�O��>�7�u
"�nQe�)nB K��U�Ɍn�&T��p��l���r�LU���Ai<�,����uG\<�J:�Z�I�v�a���"�s����~�}C'��1
���Ŕ�t:+������&VZ9kρ"�B	B?�E���D����¾�LY������0Ii�R�s3��Qw\pjZz0��8����7���^�f�R�~�pӆ;�A2���/w��ϖ�Q��#ձҎ��-�O�=>w�&�	���}��v�$\���]�b��t���l*]O�)���p�F/ÆLMu��]�<��f���%�n�ܶ�/dfx,�j�/�o�M�7fy�$sjd��:���S �}�>5���mVI�2mטD��i:�@k���o�-�K
3�=HV�&�,�l���DMbXK��D�*��r�1JM⬪u�I�<g=���w�O�[۪�S��G�E�P"�*	.>{6-%�MBK-��uN�_��2���NK�v�lk7�����n\u�MR�C�����{J/ڍȱ�B�P��ԋ-�my��ҕ�?�D$�%��j���*��0���x�{V�͜�j����5q��n&�̘i��MZ4|�<�]��E���D��V���Jz� �*�
�Y2�� T�X�Uփ�
Qd�i�I􃍓��hU�_Q�k�i�,\���N�:{w�H��fҬ�J�#�j;��FPy�0�����U�Lw�V
J� �:��Tb��jK�I,��Yi���1�����E �w��e������V��h.w.��Q�\|c9���R��s��j�TpV /�Ǽ������ܿ`��#�y�$V=K�k�����x���g����\}:����\X��;��۳��d��]1U���[y�ʜt�N�M�Ɲ6�Q������'N���Ӝn6��o���0ۢv�D�r���0OA�z4X��e)�{����U�����$�7w�`Ɵ�:����m�~����vu����o?9�uW)s�'z����
D`h ��}6U��L�����f���K`d�pi�t�|�����Z'<��۽a�$��d�*���E��Z>�����P{o�ق�F78��l�.���K3��M��ֱ`����9�;�,b\/��M�Z�!�Z���S�K&�3j6�#v���[�r����K�� �8����oƾ��ht)~��Lx��[�n��~��n��� �~�)�wk"� ۤͺu��@�ߍ:��fN&Y'3?݇_�U��R<C	ˠ��%>���9��-��V	I�:0�Vˀ*�wAA4n��EA��tQ�EHeY���N6�(�^�U�}�c8��� �R�����L8�WZR	s�J�n��+M���K�d�c�ŗ�H�ᡚL\p���(,׺8�R�,�@�KC_daE���=aB&�-��
t�e�2t����M��yq!n^,��k1U'	�f�zWa�[�,MkƀO�F#|� ��`�Gs�{zOJ��VMr`l�p��d�[z� )Dʂ��xZZ=��j�����*.Fi��Lg�S.ӥF�����838AG����Ñ9�aRx�t�<���,k$Lr�����s�2:^k4��i�i�����Ӛ4��>Z����5�����ŗ��S >�pi��QT{X�	og�� ��^m�K,=�q͖7�TD��.b2̐b>��^
� ���ho���m�PNn��sD��\/;���`K�K�����C��}J��!@�R8��8phx��u� �6Y]rH� ��;0qA�S�=Kڤ�nQ,������ofV�vc2��d2��.l)Sݫ��^��V쟨����@�\�$��o7�ء�g�0�a$>\M�Rw��j�J4f#�j��}ăY|��HVn):0H� �f�U6����_��պϺ�����th����?���Q	p�*��A*��^����i[g�$\����rzeh�
�qTǙ$��AE��6L�T��kHMF9g���o�#����	��Q���<�:�;F�{<b����@jy�C�ӣ�,|�1a�)�I�.¶.7����S�+:�̀m�����^��H�s�����a�T�8x��u��N�P6R�|����S���FS��Y��B %'�?��8C�[z���<��XG��32��2��-��xF[�,��C��<���P5�����|�`gh�z�jˊ$$� ��o����K[�Ȫ����C뇘ʜWݵ9���� ��7>\�R#����̂�ի+�i:�b�,"�L��7�J
�e�x>�vt11Z�%e�9=R�,B��u�[�o`u�k�m~T��-%�hh4�@�Ϭ̫��q%��8{��(�KT�����e�:B+�8f�����nrU���e���b-�"8
�n��n��-�t ��j?nG��<���tUx�
�O�ԡ�\��5q�ɒ��u���@��H�|�s-fr-�مRB�tc���q��;�EG�n�ٹ	6��U�4�M�N;8���/�R�F��S:x��E"p���d��R@������Q�����b�Ib�K� є�k��U���A��yP<��I��V��x�ݧ�����hd��vg�Z�{�c�=���B�\ �/��RE�Be:�B���8s��}�V�J���\�tE���e�:k������8�]]o��T��/��TD���o��QM�%l�78X�`�������AJ>�G���R�u��5YX�zzħ1�h����ڻ�˿k��x�X�"��
�?X�b�I�Pr �X,�p�n��,���W�NmK��ï����Y�lpU��-���5�d�|���*��V��u��$�-9��[�O�j�&7h2Yn�iq�l�޵<s�i���"Ӧ�kp��6�w��� sX�n4twY��8�^rj0���~��*5j��������>ڜ��� �2(���� �l�ڣS��������T�S��>����vovQ0��[�b�_��ՙ=YM�����0'@�Iu��"�r�v�7/�R���^�v@�}\AS� �b�н��J��C+�-P?j����l�|g��cZ�R�5|���X�&N��ˁe��ۈT7A�UӐ�Y�󘺳�&�H�*����J�f�O�����仳7k����rR!�iZ���9~��DQ�~�>'�w沓͍_rf�֟�FB���W�u��E`�4��Iv�?i�	~#rVΤ���h�&����*�T�`�� � : H��WOJ�Z�,9��j��R���VI����8�7���BFK[T�������:C���^��n��٣�3޲Tٴ#�ԥ��n��n�u�L�B�J�����L2�L�a2��	��K�y��`Zto�����E��޿/+�.6�|�c�@��j��0����� Dn�(Gy�-�!J��*�o�A9kI'w$��([Ή�,C��\Y��3Ũ�D�g����5��$���|4���_�/qh� g�c���p��؄E� [�[�;�窈K�$s��\�� ��k��D�J;po�� .c�m���a�A�x���R�o�O���E��)2��2��6Gd��+r+=^��[��#��Q ,F'�Ϫ*���x�K2�v��nO9d�:� H�D1��94�̵���a�w�+�(���Y��Α,3���f�̥a�}KfP��/��،�7������S�+�<x�<�v�#�:�5�T������
(ܤm����(�������@8M�^�j�xc����vK�XZ��.�p��8�-ƗR��$�
���|����G���<2O��M��� &8Mi kK�K�f/�z��S�˂EF鋝���Es���ހ7�DƢ����Z]a:Gx�����'�#��'�@�����v�O��X��z����SE>]����b���b`X8�0���`	!�qn^���a޴�����kD]k;.��_c6�H���~��T��k�M����80X)�/���(����,�� q���>"f��Wso]YB��)"e�Tpl�f(�*�O��d5ԯ� �nwn����4*&e��Ӷ��Hƥ)d��2R]\��C���~4� �q`�"se��G8�b7Ac2�3�����i�Țe^��5��o7���Uy�._��⨌t��������%����\6���,h��GDk�x�z���O@�V��&��,`�c
�w��"�_y$��i��F;B:$c�.[�t+0]�����p��gX�t��@����S\�{�E%�3n�bHEЁ	���B��τ,e	�����%��al�֐�r#�O�)��}�2}~>I�zUp@��#l%Q5�@��A�˹���,ĵ�d_]Č߂��|���O*��}v��G��z�+=���$5Ә�P����h_���$r�s�v3���%@PK����d�$�!��]Aq���-
�cV��tW3�.)2��;|��745�5b���Ң��:,K�*��"X_�:+���D��ZJ?V� m�T���U*r��:2P��p���
��v}f���ɏ����t+�-}��!�D��7L��K�&�J_��_��z�'en��$�Qk��ُAZ#yJ�!���5�U�wy}u��&8���	�f�F���О^�4��=`;-��ښ-YC�/��:)�t�����%ߎκDG6�# ���Ы_? oC�B�P�˿��a�Uc/�fc[�O C���q�* ��6�p���~#ޛ~h�<�Q{;�d{� PF�$�looa�_���?�Ȥ�s��3���N(/�:��'>�VL�i�&5�h�4z��*��v��H'1-�>�H{ �~�_�O��R�]������d�"�2�z}vRk[1���A���q�;��U�G5��+�ׇG棕a�i�#=��������� W�A�{�IB�l\h�wX �UGi����&7�\��m�!��iHN�{�)+p��:+�}���C�e���W�������U����n1�	�1�NL�|�m��JR��)�bĿ�p�����4�ݐ�:��3�??�IƊ�>��'Vm(�Q�A
�!26�&-����mdQ!�V{#�)��{[��p�T�i�[����Sׯb��Xںv�*��|Fp6�W�"��os�Jt��X�����ey# ��`�h��3��<b���C#3�I�vVô݃R��vT����T�� R���n�|�U�W���� _�/g�� �
t�ʾG���yy��b"����A��(��U�ܬ��P�������1r�ZҘ�w��<���i������K�����4�q���L+b�VF� @����!�͟�h,Q�Uc���*5�Sz���LB�m=��2���؅�A�+��B�
��ǎ8}�r�����[��8O����a��q��N)"���{m0
����7r�Eҹ<���E��t���n�Æ7Qt����.�D�I[�϶�l����<������˹p=�%�D� E�W[r���n�k����S>�8;���|�g�q�T������4��M���K������$�vqf����ƴ	7�7Fn8uզέ�RQv;^��$�5���P ѕ�xH�������I!sٳ%� 3����%�u��9�7�e��2�,�ތ�
P��5�9*�M�/��֨#?�>��� .�S��<Ak�&��ѩV;�J�h,Q��q�?�Rj`�O��/U��#o�Ta�+��V�ZQ#��e���������-̰~U�nu�T�"�͢?�<\����S������_��FϮ�F�#���8k�����<Qf���a1y(b6+[kv��f¿��2��v�.�hiS��š�^m������,4OO�p������_��#��h��>�j<(oIa@/��W��?T�8�E���y�=
rN�f����O�p_!{g1JĞ?���p|h|���~���PR��a�I�k�� �t1_a~?@�9���=,�z�&~��*�b�M#�-hd��:�/F,E���L�[X�IQ�L/��	�O��$K�����2�5v� i�$tx�ل#����4D|���qqŻ���V�H=�];:�E�Q�Q��8�8\%��Kw��]�{S��/8����$��^8Ö��T1�Z�,{�]%q�V߯���;�6�R��M�U�d��d�%~��5� no\Or�he�uw� i�e��+��A��~�0|�~c�#�Q_����y��X4�.>�2�P5�X� ���Ŵ�c�	m�yBM�?���*���I[i���,���͈X�O>�� ˽���-�mH� ��e�iɐRXE�U�xT��񀩳3���p;�}�N<�a��E[w�3��)��0�=����@cY�A����]�Q��7�KLm�(�[��YN�8u}f��o�kp��Aj��$��S�Y�<tHF&-���=�JY5��)�%P�L�¨�ikK@⋀ص
�mLpDӜ��T5�병��@��z�vL`>����/+�$A)�g��%��;��~L�KG�zL ��K{�I*	�ߐ��Q1����y�h��IvE��׬�u4 ˥��\�F1Mw�86�$O��HR��5p�y͸u��f����9��K���L���^%T���}�.vuY.��4ҋ�9����S����L/$Dי5�F������4����>��Y��_�h��t)��a��/�2*��@����`��=C*~c3YO�rAt�i�)�r�G�5�����z�Cu�|���1����oylը�߁�zGü�}��\�����(�����ۉ����"��9>}:�c�o��
��I�FZ)�=3�G��ۋ�3-�k�0a$�d:����z��뛤���O/�6�M��=Hܱ)���r���!-���w�ZE�n�p-7�������>�(�?��&R1JA
�S���U��d����r�A��kJ��۳5L;up>���<�u���<��������������w�#����4o^��K]�J{�(��ٰ�&r�|�R��X"��+��k�)k�׸}�s�u�W�;`4p��<�;�G5p��q��ס��@h�֏���Z,湀����`2���Z��O&�V�P<���u��5d�"���~bv�(��(w���U�D�i���#�7���+�/g�{�k�>�EH��*��{	�O:#�k�Rq�p�V�qN�� �_�+���l����$GN�ۤ�>{=���1���!�"�O,�[��hr����%��(��a�ۇt� �j�c!�^-m�x�U��Ln�[�u���^��x�Έ���7T&X�B�T.,��@���:>�����+1�*P���*���0�t���e��٣�K�h�1�m�
�8N��Ҕ7�)�nwx��0[X.̎�F[�av�`ȑH	-�hރ����>*,o����� ON,Z���pM�us�C)�_�D�%
׶�>���b�L�Z]�C��S�S8��c�,7s�)������]>���Q�DEh �I&G:k�P��\T|��}Nʹ�"\��Mk<���M���ɒK�$��ON����8i���Bh���w`M����]tp���.S���.���[8��!�X�k�"�!5�%AS��7T��I��������
,�ƴ���~�<���MJ)?тذx� ؊�=d̈� o���>��u8����0��7��t��>
z _�j�{YAKW��v��qX�K��@����|�`��̭C7��H���y��;4�m3�'�� ���0����m��}�l�����c2�C~��\D�K�8�i-'�5���6P��җڹRaJ&W#u$%)=���F�0G3�>��������f�~0���H�r��l��Ïʱ�}��� GD[�գ�k���D� �6��	�T���0Kϋ���Nɢ0qM�E§5; h"�0h��zpT�p�?��|r�R6s�v��S&8�G��<�[ '�.z���K���2�]���E�:5 �<W��ZZ�)4�J)��Z�l�$��UY���tDw�?o�f�ʸ�Q��.��Ӷ���uo\b�޶��д�0 �S�땣�M�����/�����C&^��d\WTs�Hj�տndq��@! 6�+���*�z��������}�d��z�~�hN�O�+n0k�7��M_G8L$n�Ҕ�j�_)E����!�DW'9�Y�	N�\���I��W��m���/m��j´&1]@�\o]�q7���Y�)mmwL�(�e���b�9U��H��`L��z�'S[��TĚGaǑ�������}��s��Q�l�a���Ը���뼭˜^wgnh�%kH�
���r�M�4�(�ym������7"H}�;_c�aP��^�	�d���d@}�O)�v��&G.'/���/nݱ-)9I�r���q�Aצ��^��Z����:��*檳��?T��ۣ4�1��)�X��j�D�;/(�|�X	�h�=�N��e0�>Nʀ��+8�^����4~����DMzl��<03�ݔ,�	?@Y( o5�Q�-e6�d�d��Xy�U��e�?��r�Qd�z���`MR�3���o�����-�հ�@�a�բem���r+�����8;�xJSa3�����:�I�H\�X\ ,��G��j`��ѥ����[4w>um[W�Qh�G�m����� ~i�D��v�*a��W��=�eW�K�ʔ���9_�ehp�,��3�?˰��Yc^q��A?��U�\��n	9:B����v~�nL~=�#�<^��aw�T ����ys8S�B��9�J��Q#t\�f �sŇ?�ȓ�r�̪J��{"�,2�7��҅ú7B<[̄�@1��MD7����/��hhǥ$;?&�NK��K��:��#� }��*V�%�S{[Rv��4���Gf���,��l�����Y��jc�Ll�)�UWܢN�i��ҍx��ϕ3b6GwШ�~���"�b��q�`�F�rc��u�p�5��������Q�M�fN88{���8���G��^�@�5 ����<����M�C�f�hDXX�\���pt7�ܘ-�l�W����#k�($�;��<5�Ј� -4�ػRq�3ȹ�?�	K�RϤ<ZFFO��tߚ
]Ki�HN��d�٠'t�uX:JD�GE}������K�Oў�T����� ��<����A�m����δP9���t~a5���~�X�"�Q��8359��ݎ
'��0w�;�,����_P�H?u���4��p�B|Ge2�]�՚�9�S��u�bp�p�dL%=��5�	D��í/������~0����Y�j�CU�̻˒��94��B2�c)@xc�%G�fNg�G��Y��-�WFt��V�}F��uB/��P�z��D|t3+�vG�,�5ř>���Knn��;�S=F��s����[Ė��ky�Pxp/����Q����s��q��~�{и[~��oz~�@��^�/
���c5�^qۥm�Y�R���,�UzR�壨�.���4{@p�J����y�b/�G���T�YF�����_�׆a0���UC��0��ô2ߌHNj��[p��;��EX����vÈ�G3 �Ȭq�v���4@�2��Kec(�K�!�:�=������]v�+L�23*[IZ��l��D��
��_qV�.J���4\��l5�������%�4\d�`@#쨎C(4n�Z��C�
L�	�,��˺\TM
(��֯B�V],˾�i&`�u��Vw�-!��c)�NnV�<(�w(:Ȟ���Voa�pj���PQ� U��]\�4܈h��+���/�|&I`\��5;�pM|�4w�5C���*U��	�E���]M:����W�1���P:+Ғ���'fJj��|����_����-ٺ�u��3 ~��E�{��_�Q%$�-9�F���j���;�^��5
�i��o���	]oX#��׫ߗ3G��>~8���֕�J���Fc���Ĭ��T;,'lw���.���
��4���sW���73�-�P�����g�닺�Udۻ�-m�Ut�����~UE�
 �T�J�]�w�u�w$j#=�5�� /�Ʈ}�d/�9lYG�Hn((i���x��>�dx}���5�|qC�{���3~�7�d�vS��{���0�L��i/��&bUm��,@m���:>by���d�1����>ʜ�g=̄� o��@X����Kq�x ݋p`�� i����/�P-��>�3�w&G�����S���A͡Q�+%�Ґ��w��[����E�!K��[P?���]��B㮇�����0�ĐS�<ڞ��z�ic�������t9"���v\��I���xO���x���KFL�f.k�"�ӡ��N0`jʞk��re�^����Ř����:���\���w�wrվbu��Sϳ55�[3%t�"�w��C�	��$g�Z,��U�CJc�-�N��#.L�א�k�pu�j�Mq�j�-��n����򘅑�̍m0�]��&7��=o<+���x�3w� /�7���W+���{�v�G-��������v���[�%_⡑��fp�+ǀH��l]M-��=�D�B�%<�ؓ4&����i6i�:�'UᏉڶ�"VX������Bt�P�۝��<2�w����	��F���fͮ��㽉��98"W�J����R�T|ix;?�4zu��K�����&�� i�;��������fufe��������q�� �H���ťy�L���e�����-�
�c�KNq3l�F�r!f=�Iv�'\������ɤ
lB���c���]�5��vvC�{��חg��^�&;:S[���%�j=.vw`,��.���Vɻ����B=��������l�&����l��|��v��\��&$�Wϟ~%��e��/�
��i�Թ�c��FΓ��2����'TM��7V��)�kHU~&3#BN�?j��rR�w�Z��j�@g[��(m� ��]#]��f��yճg�UT�����[��y��FkE>�T��q�Є湴ɉ׋�_t]'�Xi<'/:Ǟ"k�-
p��h?4#�=P���=E5�ڿ;�nr�?�h@
5���HE����#��뗅�!�S��E��(z,�Z&���'Rb9���hC��q���"1�K��	%K�y��a��R�A�^�}6��cؠT�R(A(+�@n
c.L)�A�g޵�w�u|�$�dV��0'��PR4z3/���gmv��u��E�5�OE�,�s��#��鈽:]Ґ �d0Pwӯ��A�릥5�"%1�^Rⓡ3'���
!� �i�6�D���?�uj˃�A�N4D�S��_-��r,��5=$%�,�XWl3���������N�  �"Y��vSU쮶�%� HL�~ۣ�h�k��^$a���px��ބ��r>�Y?�����l8�W�ʶ�����M�YT��g!@=�Y�a阧�i�KX$�ݚ��uIg��>(@�h�0?QƄ�;>%{��*䵽k�����k�"C6K{g�u��?�]�b�׆X/B!~ݕ<UB�sl�G"��ΰ�Z���[��T�K�Ѓ�J�����9���^;�~:�S�����:����б�:�����'aY�����,�@>��;sV��u��ݯp�s��8��`���W���Κ�a�"�<~)qQ���7)�A��x���,�����Q�B��b��;�9�[A\5�9%L?|鱯�[mp�}�L=ɺ��5T��V�ɪ��NUb��}�鹋����&˓���^8-$���+�0����m��n����%���%�Hªݑ���A��ba<Z�)szO �����R�z'Fj�+����-��9D�f���tyٯ4Y��c��w��~�ߕ�m����.L��Yt\w�h\;k5��<,��E�|z�d��,c�z��[���<��'�z;���?�>ݨG,�k9�*��Wn��hR��Z�$��q���0�qt�d���-��E���������6SQ(�#r5�6��Sd���hGI[."P,`���&������}9@3m �)�#kZ��&fȱ&_�t3n�W�m�������|�{y�Q�)2v��S`=���1��SM�?ܑ���h���}���4���V��>��o�������iPtТ�遯sg��2P91r�[2%���Gګe�Q���\UQ���6�Q�K"�.K
N�4v��o�����f�%N�����`ߵ�悥�p skV��H�����Jd.�P#�yb�ϰ�c ��%��D��)��h���X�ij���Ǆm��he�el1���e`(\V�>[bHބ+G���J�و	1��UZ<�@��a��//�&��E�T*��ku��v�f_��
��,�>��0㎍F�|"^�[��2�� K=0�K�5P ��L�E����>��R��K���Ɗ\��/a�^߃y�G?~|����$k����0�v�j� [H��U���Ԩ;21S�~QP
�7B���'Tn1zU���3�r��%P���⼱P���Z�J7�c����[��$C�E�����&����������"��n �D2�Be;�"�ŒMaR�_ǯ�J_��4�/5w|>lk9����N�(s`�s!���n��9�¿쨉����F�37ׇ1bɤEl�t>J�JKLb���	�F�9��avߕI���CNi
�ơ��:��! ً�W|�
pP(�.]8ţ�!1�qRjp��ޤe_!Ǩ�3<���b��x7M���"���u8��E{��8�}Ԅ�0]Ժ٬i���F��E)�,��
$��j�Bc�M֊K��YJL�B|��`��XI����3Z:��D�h=r3���*�X!���f�an����3��5�m>蝊u`�
�w�1��o���&.i>�h�u����s?W	o��^��U,��#�Y1�E5Ժ��y	&�:U��p�oC~Xٷ����Zh�Hgn=��ϓh��������A�\,ܲ#���G�E���P\�X��ך����l�ҧ=��e�,)�K��V@ܰKƧ�&�;�K�ǣ�9&i�R2��}��HK-�@�f,�hW�����{LH5X E�ay#��@L�Uu�����Xm�ou���ڌ�^�դ������,��bC1�u$ 5;rL�!Ü��/�}� �z�`o��,�% P�لI�D�t��Q�I0O~Ŧ�>��="�V�\�������u�G�E���|���ʹ�%[]�7.�;v��(�����k"��ρM��M��nrw�L�s�̍�,��6O��+�0!&��Λ����ʇ�5M_����9�E_����FY�.k�xA��|�7�8ā⛎��|����# O9N��a�2YQ� ����-�0���s�0��Q!���y= ��{��ɹ���!	��%���k^<���ob7�li�r?��-͖�=�,���gߓ��
5�᪟���4:RЛ�qmb���zr��I��v�
=�|T�<8M�UZp@^\HIHl2#l�"�\V��
EDU<�S
�
qJ���.����r���I%�V~��6��oP�+��;D�ˉ7�"���;�������\��e�KyC2�vh�i����]�e�fZyA���@�+�H)>&��}x�V�0��
+/M�ὪPkoN�&�����W�LVƠ���5+A�H�`�0�Q��³��d6&B��f�]BXC���2|�?b���Q��t��s=(&��o��&�0OXYq�O5f���K��ݧ���rm;���{u��7$-|xO&�߉���m�Ui��@�X� ~��� L�t�mz�2|4BR�q�'���E�ϣ�+'ݢ�} ��+'eU�����"��S��1�0��`�4�\��(n��z�b4yB_��6�E0�=�2E�KF�A�����A���E2���x2S������Be?�"0�>�m�#V��3�������B
���EC�I]��ܮ
y�<UG��<�:���J��8�%�$_>�a��$�)y#�A���\�Sҍ�l�L�����Z��RG>�b�T9@����	.E+��dA��j�O~Kl����-:��3*�H+_1^�W�I�PF ���<@���[�դ*����&Z{s�v�A��v��md�8uc2�ZR��J1�Ik�r���Ike|i��uġ.�%�=�obU�V;u��f܁G6IJ�Y�*(���}"|k�]@�EFw,I�_f���@`�:��[��6�;��Zf/~˲�������'�$��{���6 g�ջ�bl��1%PBI�q��nk�I �	�u����"]�ki�%����LG��6�Մ�\�5�d����V���`Nq�W����"���[f�{I�Z�@�uX��}�Ȃ.�|�kt}�T�������Y��9�C��Lv��dX�����i$v&h�yUjl-<��l#b�8VNISN�&ުw��%��-��(L	�pe��ħ�g-?WT�<�d��!�� eob�޿��&!�rd@�O�q�y��ށ�⪾D�$7��*ޕ�΁�#P��l�������{lAS�+�)$��hYL�Lc6R�K��-2QJ��1��)�qEÓ�m��P+
��7�/��h��J�~��*\ӛR�h�`k��h9!?ᙴ�6�״�1)�wY�v;7|��?4�
��,>:�G"����i�%Ey�7�*Ru���`�\�.��$�?�h�%��=
w|�[����,�,H$����#LթG>��bN���~�{/�ݨ����H�Y���d
���2��<P��\���X�Ύ7�*2�j����B���B���_D���U?��QOC�iPFXO�4X7>�B�1��M���tV/�����E�æ��5��=�j��-��|�{�jN���~'���떥���7�;�V�K��t����ݵ#c�F�3�Ϋ�No���BcDIU._�����ϰ$�FuE]�,��\��D��� 2��q�!6�C�t		�p��l��
/����L��	�Bs���,4��y2��yi�	|�ե�K�=&m�{�� �.\�^�u��v�ͪ�A}1O�G��n�f��3��~����1�C�AE�C6�"��[�"P�ũ�;�$��R��C0ȄR�d���_��|Hs���]�+��5�u=�����\��z4��+�*�N��mo���c�ګ�gN�ΰ���S��DW}$vХ�#��N�[�V�{��4G,�N�cj}��u�<�ʤN�]�\�2�枬�Į7�J�5�$�6-�֜����?�k{�`²��]	=w��N�vn<S69���T�����i���
��F�a�\��|���4z�\@�b�Cw+ת<M�I~@��	-M ����f�8��Ìw(a}�`�uѕ�
"�f��T��n�*�d	CEx_\7�C����ϊ[�'�3�iO���!���yܚ�#ZHsxDy_R�y��y}(��R)�=�����w��o��"�+�d�8,$���`B�����m�r���/nۘ=Z�=����
�m�x�N�I3�c%�
�$tZq����m'=t�D�ƀ1���B@�V �ŉ��xm&KQ���9��	x!q�5$�a�s��M[��`q���s:��v���y��� 9�����r?8J|B�	�v+���,�%=����K�?�����ȨX�5����Ǝe�7�D�ѝb=�1X���+��ߡ��W�w�Ө�~rxޜ�����ۡ<�~�`e�yv2��:�;R�iJ�t��?���
�~����Q�s���!�Aj�.;�b�S���� e�6Chq4f�M	4`�H Шb0P�`�W�"�{�9���]2��F`���4�j{�%gQˈ�(IW��n}�w�2p�_�X�&� mzAHM?t^x��m��ʋ�yH$l�������Q$!�=xYZJSWO.ŋ�<�&�.�y״���x�A�'���	V}4�}��'Q���JJ�J�S�p�7�C4׏x��J.q��~�!M���tom���?3�꿘�b+`)�^�K}@������Pk�J�&�!�[��\6��u�ۓ��[�/�U�s�2"!��z����L:Ti{Ks�)V)�O���bx ����\-���,��E�7Ö���Ӳj����R[m!/D�`�B7��n�+՝��UMF�fޮ�Eȫ�\4Q���ي���( �q�$���
9��������&���ň�Ze�!I����#�7J7� %לb;^xd'N�h�]$f�H����"�ݝ��r�� �V�2��կ����XX��w>+�)���6&��vZ`?���ej�wy�X�m4�+L��+
�1�ЋBqaB���}|Ov�]��C��
�m�(��	Ǥ�~H�T����9|	�'[B���ː
sBW�19�ai�b�s|��1QP1/��A�v��$3K������,�o!)��1�������1?6p�� 6�#��0 �S�z s�i���I0�V�3���h\dǧd�
���STȵց�vW:/g��̉�C���`oF�7�PSX�\*���.�G�4���JK�f�%�!�	�IW�ZI� ߲}��M�M	��Ê�RSd��8�Eʮ���ւ#Ǩݡ�d��	=+��.�0�E� ;���,�B�e^�_r�<oKf	��+�wX�~��w� Yiy���;�t8�4.��/8�S�V+��n,��Q��s�Xγ�R)"�3��tC%���{�(������1L`�>�Di��a�l$'�ɼcR��҈�6��Qz��0���x1��5�Q�7���N�қ��4�t�(�5!���I���Ju�+�E0��~;��[���kacd�	X�5[{�NUEGмmT��r$�e��c���r�$1+�e@MCZϒ��X�ڏ���y�^��;�k���)��l'�H��?#��p��(�&o�1�x���z=��,��|�]�G�)ی%N�#l�+�3d��/��1t×�T� ���X
~J76x�؟]R�ı�t8�JTE�q�����EǙ�ӈ��V"��ś�M��FLrF=�URH�{U��g�:0��޸���{���oQ;�ZJ �	K��9�I��-������T6����q����{&~���b�Y���V�C�SP�
�G͚˦�&��ث�v�i�1G�1{�������/÷�k��R�h��!��M�R�d܄v���H�z��z�s��}��S��,�*��ˑXÅ1���h�/T�����YR�\¥�K�D���%��I>QD�
�>1�'���/݊���?�����}�׸���}����wtw�A^1ʵ�1cm�%5]�.}�e�Mu�u0 ��W+	,������-�j[�2�P�.�K����y�-d�ű6|��U$�(yT�H���%&�T9Ӧ��˸�]G�_��z�o����_OL�ـ�a�T����cF]����&I���_M2���l�y�=�������&V��6���u"I�_X��/��#2j�5$I�z�p���к��*�D7�Kϩ�b2#	�c��c�ě�:u1%
���{�s�.K�o�¤�uS�u��20bE�'����WF���A~����f�oi��/Ո��E��
��=�r?�6�Y�^��|D�ݙ��:�.����7��#���h����-�q����Ȅ	(��">�Q�eg G�\{ʄj?~�"��aq�W6 il�F�����d�;��sO/��P#Ά����3r�,4�����U��|���!fɤ����?�ۮ�K�xܸ+��/FA�]y�֘��/}1g���[��;�?Lh�,F�4z�AP�L�8>�H�6E���	T�2��E�|���};,�	yy����r�M�&N;�&i���0>q���Sלm��ڰ�&�t�\�̏i��)��a��p�B�ፑ�b�ˆ\��H ���"s�(�Y�'���� e՗m+����_�N*��-� p�<r&�p?*_�q?�
G~a���?ׄ�i@��n�vL�_0���V�#�B>��k�^�i��5!�^�(���Y�?�t��k�_�5�,P�S��e�dq�x�`���H{��1�zh��D�,�� �������(Ք8��+��e�&'��"
>�=�T��k#q�+?%~�5��>����A�K�vhY����G��G$�|RN�W�5c$���Bi'�JeApm���r{Bv��r��}��د��'p2 ��Jl�c=Ob\&�"ݿ�S��j�`G�u����'|�A�h���]�=�:�����+�v��%[�]{�q�A5-�ߤ�5�SQ�H:Z��_�o�?���-��.��=���3S���!�����:�,w�Uz&�Ko�>���AU���	g��|��1�>��9E�Py�<� �/��"�	E?�m�	y��Z��pqSDP��[��y��4����H��I5ro��5w��(�O��l'���x i�V��Cw����[G_�$��4�P訕G��H�q�C)�Աӡ� ���YR�6���� ��N�5�8:�p��-�U��1�� �������Z}����V-4�~�v�חûfK���u��
�a����u5�`��{���46�M�����@YE]Z�\�c��;�u�2ulYp0����9�q�W��#��f~�l_�c"�C�N�LUdZ�%G�e���Zw�x5��&���:4ݣ���M�%��lQ���N�2����x[HK��U�7�@�If�Ɍn+G�i������W��Y���65��~X���W��:d�wۤ%�=x��4�y�m_����ƙ��~���^��E��������,_�(;���e��H��[�m���*۷��;z�_�qR�J���~{o�@˰��lg?2��&͓�#�z"2d�6�6�I�N�)��;�m�&l��$�*.��by�Y��Y�