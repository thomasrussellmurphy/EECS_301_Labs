��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�i��a
Α1S%� �uj?�L�3��TLei-3^5]E�$��f�A��m�t����&W����*X����i\��n�$����g������ix���V5�XqơƆBL�!��Z	f	D����F����}��'��[$�]��Ֆ�,���B���;^膭;r��te�̔ �<�p��姣v�T���7�D1�R#�ǋc�g)Xx>H@Tz�c��oa��:���~g����ž��4� ١F	OgzF�la>d�.)ϑ1=�I�S�\6*D���f{Ѭ_�G�����6�T[�@;	M�Rg*�0����Pa�ܧ�7	�yl��fel`�h����ʁ'e�����Q���M�;t�	$�L^�x��� ��ȑ{Ab��%r��i��T����&v4�ʸ���0��Y���{ �m�_&�Lh�(,����ę������o|�d��QT�8[� ��䐡��k�\��1���͹�������<?�"����2wX_���;�#�6۔�s��=ǩ���`Pp���&c���&�A�\}�)��=�cY[*ؐ���F��Z����Y��[T��;��"�GѳZ�04S��,�#�FOշf���ˤ�5O�ֺc��,70�q��q�w��#@k�W��{��;Y��}�
du@WЄ�<9�M=d�4���ǞM�YΊ� ą�y���{��c	7���aR���I<M)�[=��/��f�ťl;㱡R����f�Oɠ�w���:{�[x�S0���X��⪝Po?EK�GoNe��?׶� ���x@/�ǟ�$�xi0���Dkq5�L�$o���Y�c ������z�.�U���i�[�?<����΃;!�{�Kw���@�E#��uh�hhq#�ƥ�ܤ�+R՟�tהB~Y��Yo8G��?;�GQk�=���%l+5ldI���h����E����q����$�c��",z�D�ŧ/�5��[Xq�\��B��/�j�K��I_I�5r�
q��R�Z3���Ǝ$������p5ĕ����AM��=�i�^A`V��q��[ �e�L���xs8�5���_���9mރ��)���p���AM�ԖW�p���B�'��0T����|PI<{��aۮ��1b�G���V��%{tia���ب���g{��aL7t��A]:����۩�'���f�@�q:��Ò�oZi��cT�m��gK�� �@ME?k�2�L��ھC ���G4�$P::�#]&H}z#�Q�o:�����It!LL*���21����l�vo���b�-]�
;F��dX�U�$4d��.Uy�l3�?
8��a�k�bq_u)��h������)Y�zE0�Z���!�^h�����8�s+��2 0L���yH�ꪨ���|5p�4IC3|y
�-�̤e������%m�� ���G�/�pO�l]�����	���D>ώ�6��Z���¡�i���b��y���x���U�H���EETf�I̥�����G���@l�ܹj2����<|�h``��t�9��� Ƃ���@j:��`n����Q��=���V�Mha�nd���_ud����O��@��n�Ex[���W��|����
V����/����muk'�8id�hϠ��8��XN;[�����(I[gmX�"0$l���;��?�������yr����@���|�����	���~�E���۶A�	�m���O��z_�Դ"g+>��@:�+Fa{F<�X�{b*�Ŷj夆�P��I��>Klu;�i_�mJNw�B�̈́�N��6�w���H�j��ݥ[���1,>�7W77S�i@��9�o�A$utA���Ħ_U�,���Ϩ�ɻWs�,���k���ٞ��s���j�aP�=���n]^�[�h�*��8�ȑ��������"Ԉ�`�uĩ�'��{��y��R�."� %��.�E݁4�8�{J���ٲ�
���d�#c��	,�ֻ��Ex�L��*�s��>�DP�E���NcdCR�'$w����Cw�c�YѮi�;4�ʗ�g�P��R�G�x�h��e�1ӣ��@���I����.��C��h
�h��6IV:YL��(���3QW��9
h�U��|�=p���k�+���rxČfZj �kܮ�?�l�-.�@���0T�&���K����%߳�|�B�n&&��Gܜi_[q1nD,������!����DI H>u|��t���R�e�~P�>�r�Slpt#��s�Q�t��˲<�K���ʨ�<��a��tX�����I����C�+��������R&�*�����V�o]����3i(e��>p?Se�!9rg{V"�,D�P�Ӹ�J���E��VY��a�.�Vm ������]-j;��@�=;�3�]H����7T�VZ}�U��*����5��6r���"�UW��� L�]!OL�Mg1!:��}O���r
��R�f<B�����V��|�mx(��q"����W�n���,��!�UF*`|j������+R�>1�/�L�4�@R6���>�?��Rz��z**!ѧte$�r���(L����)�=+m4
�+��y��X�Z��CSh�kg40����OW];O�p����Hb`|fpcS��D�琫O7�R񏶠��7*7�}]cW5�޹tpG�K\	Q����kWcZ�m�(K҅�oh�B�����_/^�q����1�����yx(\
{i��� ����v��C��ߟ�ⓞJ5g� �%zBN�mߋ������2\�KU�e�s�P���K�i2Ky����po4���� �x����n��ЯY�A�SYJ����9��5�����T+PǢ:i�\)p&M��#�k�[0! y�#xe�̯��T#k;��ИN�$�fIt�o۹<����������Y�U���%dw��f��u�JR���֢��'�]���<H �;�56�����������,5L�(�����1����.��G��V�w%s0�ͻ�Yv����ze(��Ԋ��(A�ũ�E�j�4���|Xw�m��?n	���Y4��0�y�2�p�#$R+�Bg�?���1��-�w����j2jon�X�=4�c�����	��wS�h�j��4/~�ݖ)�� ���W��ɨ0����?�@�]%4��&`K��;��?4-&���t�~��P��Z�<�2y���R��v��0H�!�j募��{`B�ݷ�g@J#��C�����##ZN`���O?�
R��_W�2S��O�I��ٖ͆�dC��$��Q���|*�Sp����fI�m�8'�Q�w���Ԙ�*��M������J�R�}_zn�9)4AK�5��׆��1C��[� #r`O�܁�@Y��1m�r$���a?�N��P��|����x�A�� �� #I�k��	��X-t�����`�\�Ɂ��#W,�Lxq"��'i=��ϸBd��-��H&����`�����j��[AE��BH��)�,*�,v�L������]�?S�;#܈�g#LU���?�ɈSI�G�3�5Z<��S��O@P[�DAr{��$]+M����η۳�ѽ(d���lǢ��9�l�;�U�|�� x��wN{�uY�a����늂�"D��!&c�pX�'���{�gTK�^��8�����`�/���_�0�s����7�")��M|Y?�^�Ts�a)�S�7"�DA`��������_�>'8=�V�X�Q�1"�Vy�>���vRܭT 3����Za��|OI�91��A���n���'�@�d5�������^��&�"��ճ��U�f,G��Fl��3<�Niӓ8䜱�+�;�����O;��6̄���b�H`�i��Q�����Ǎ��H���Q���v((K�ʊ.����|��?P:����yh73r�fO��"�x�>�#fs���B@T�K�,(KV2XJl8*�Dn�l��9(:� ���n��d���0P��ل�8'�`�씂�Kt�D3I[K�;0�~a�;6ab쵂���ٙqb� qqr�Qу��7wt�xT/j޽���(�R��bbu��1E���@uka�r��z6���1&��wpT7H��~tx���q���>* ��X���?\��#�4r�ddW��-��_�0Մ\�n��j��J�5/|��X�_s,MNnT+�ܯV����-`|8ݽ<q���W�f�W.��X��aR��jh������g��.�6�`@#���"	+?L�}�t紹ZR9�5*/��� w-�k��z�mr���s���/y	L��Z	�(�&�D����ul��՝�>�-�ܭICN�w��}����Z���)���>��BGd�( ���e7�����p�a�-R� *V<	��':{ѕg`�J�B����<�Dy�Gգ�bYR"[����s����Vq<l��L�̼l�v�S�+�}���zt-���z����J)��,�z���>m��j��A�k��4�`�vMd[i���Ҿz�|̚��n�(=k�úe�.=V��0X4��:,�2� u�Y�yX�kLX̹sG��'~��rs2o���a��3���i���[7�e�7��
��?�8ۮD��h� $����I*�~k�DMs��c�x���kQ���~�|Te�=��LrFG'(�!G[�{x���E�X�-����d�jw�J3A�b�m�q��<#m���1&�dz�\�TI��i�	^RE�u�u�5a��;���SkUͱ���U|{jN��>5�&�TҲ��[ZV�*oe��_��q��d����T!p����l�r�G;�Ha��	v��&̜��q,/�¥���?VJ���mrjC�!ɻ�2tx���V-"���CS\�6ȝ�p`�;Y�X5��6��{�D}�#'��lB�ق��7_���oCBS��f�b/��S�ǧyALWJ|-�*zo$�v�(̮xb�<��]_���c�E��U/�';��Ik� H�'7����d
����/�:��&��Q��\�����nMf8�V��.eű�M�W�zm��GM�y�m�I���c��/�̤��Рe��!73Q �;�����%��p����R(�
rŭ��T8������Y0���a�����ږz�G�1������Nu��d��i�1Lbd�k�+r'���egh^���쩿�:�t����;���E�:��0{*��������>)�f)n~Tw����{�E��������`n�$!O�e���hF��Z,�C�����g$2���|b9둅AH���w]���<q�+H.x)QMyɱ ���sd#����	�5/�V��f�j`��nߗ�Y�����P,n�z��pB�Y+Qր�5�8�V�Τ��z��;}�Y4Q�E�u��t���:��R3�{�yʎK����3^�����0���4S5�<�Df@�E������m(8tI�՞����.�q�%�D?f3��'� B���\P.52�Im����7�7S(M2���[�C�ǺWѤ�_%Uĥ��ҥ�^��W�y㩛��B-.���z�!�
��ح&�	�"��?��0�r��q�/2n.�oi�̉u�[{�R9�3�mI`�;����q�ͳ ��'U�t���E�l&���Q�?,����"R�8��&�p�<���|�[��$W��	m�À�r*/Z7�I��Ķ>�2�Q��25����pI`qX�la^�bټm�`�a ���#fmta�L��ĔXI�k��	��,�4S)DG�'bN�ޓ��y`��Ùh�A���<����?�^�K_�6�$4��\+:�{h+cu�ƕ�j���<�y&�
L܊��ww	��~f����x��viٟ_˫\A�W����3��Qo��=����4��mw�>����~�o�f��:��Ej�+n�F�#��l�JK~���i�uj��ꢱ�X���+���4��M���8��-q�f�	;�ѕ]�<S�z&���\;sp	�/�JO�WF�j�_п޺y�q����;i4�DS[Շ�	�}~���e��5ʡ��JO�� 4��4�y~(`���Qǧ��j��N��c����߃8Y�
��ʍ���>���.bXOw(�d��j�����e�xΜ\'.A3���┑I���qvaܦf~��/^#L��7QܙE�I�Zz��:v��S�jq�4DXi�b�hYU�M�:Y���]M�2=�'����Vxaś�X�"-����{��. ���_����5� N{�c���[�~ǈ����@l�,�}
�:�Sp��]�N��.jІ�џ���J#O=a���_�h���S�X�0��ON2�`N�� s�)ӓ30t���T�U���*T}��B��gN$� h��x:��;�pج�R�	��,Ǖ����<�}MG}��?�L�g���Z�I+����٧�Ra$sC[���x�偩#d~��JU7�v0�I���n�g����;!tp�$�fJ2��`7�n]ʿ������[�I�	��~�&SA1$�D�Ꝩ�a�`�`+��]�yRo�J�9Sx'va���t�������7	��[�J;`۳Ms�O=�C�����������w�P��$�D�����9�Y�5��覤Oy,![� ��V��F��V�YGK0pzI�xM_���1'�1^+$��P��|�,�X���f��6��x����`v�~�&��/��Lϩ�hZ9��������9�۬T�muo�Ԟ��X� ���yi�&�x��f�4�#�4$N_c�2��R�E�\�a^M�x�B���PDa--K3�����s>�Ϡ�6�7?�Eg��|�'��J�9!#Ta��y�^Ga/�Oo��iE��?[6��@[;p�F@@�z���"i]M�Ð,T��1�H�`ݸ;�bSɈ���UM��Y���Z�j�oU{$vbjFu4���=1��������?��s%EԄ�r�������i�����`ff�|���:1%J�����k|�� ��h�/��W?~f�	E{J��\��j���3�&+(S$�:��	߮��!f�+h�&� w�B�i8�$�H�C��z )*���ݸw{����E�c��=�����m%	{���q�/�t��;�*�Ү���)@l��4�M�I+�5�/��fz;WІ�ɐ �P���D�}���Y!H@B����k�p���I��-Cj����nK���A����_�-R�r�@z�C�h��OD!��Fyg�[Z77���(�"9��� �(�j�H{�"A	�W�ՏQp�TT�q@Қ|���&��O>; �>�U��&!
�e5+�ST\3�ܥO�游��F��R�x`�~��z�2��N��)��#�����������G��B���(���ӝ/�H����<d�����&=@��w��u��~��6���Q?�+�_�)|^��0󷹗�צ+jUd&�D�Y ��6��\�|#	⯸��R��I�^0wu���a�S$�IN6S}�}�+mw���]_ ��L�+#��?�`pH%+�QgV? �`4]�ٙ����.q��7$a�M��=���pSE�Q�xs��K�����Q���˗xѥ�����BP��,��v��v�N���@����A�طE2��C68�4k�e�/�Z��B�����n����M�����ܔ�b��4�Wk�J��ifl�}���ᩂ��Me��.��!��R��O0Vh8���anf׭�d&��D�RY�.�V������;�^e�S�4e�g���9����k?���K~;?�H��}��Pyh�G��\-#'�����Ҭ���K(=�q��'��A��Z����ts��T��B�o�|�5�/S�ڈ�y=�&������X��b�B7 �V��X6�oy���c`�j�r3�q����=�2���IǼW���ɠSV_\]q��P懵�o�ɩ�Z���7�:@b1���n>�Y֞���K���_������x�>B@�N~J�{�ٌW@@�6�Y�(�iǓ��������2tb�1���pb(���R�.k��lc�B`��,o���e"=Z��?U�%��)�����En�o��o�:٣�����
���Q��jn׿-<��T�oJ\6�U�`�K����K-�X�&���`���ĚN%�R��vv�p���_&p�o�Me*�|/�/YFL��ř:����_2��s)q|^}&�,��
���G#^<d��t#�0��_T�c�~%�@�eB�4�h�p1�7D���E�rW��HS��zDT�8Ø)��iA�CZ�-��n���D<oC��m�� danI_V��U�;��C�h���F��ȹ+q�lKf�߸5���Љ�T�E��l��s�Eތ���D���?�-�E���.ZN�Dcg��:�:�I���Q��ͨ�ZyM��I�!�ț�2X�P���y�1S�T��yD5�!��E_��>�7���-Ȏ	2R�\PĄ8�.H���{��ɱ�н�[!�4!��/Vb�p�K$Ұ�����~d2`Ώ����T`˂*J6����7AY��~3"�q���ZP	�,�ֽ�})��r,#P���d��%vd���c��E{�nކ�-���h=i��rþpm)��͓�X[�48�+������%�bo�^)�d��m��{���X+���B���X�w��$��~	O藧��
M�al�Vu-$�%Ku�V2N���,vlЌCY�ܲ�n78z�&�qp�}���ev9q��_J��6��G���=���N�l���6�_�]D�1^a2��X�W2�|�u_í-塻#�G3G��������a��ۿt\��C�s)�Ob�׬�'L�h}c�� dT����-�!��-��SG���1��k���}���}��rǍ?�	R��j�� Gp*�<cS�r���ٝDE�J��T��	/˘6��pF��&��R��U��n9O�Y��~]3��|��/3bm̐��M\��}ļ��Q
I*���[O ���6y�
�Z�\.��B�y�u���{�>��$|
�H���r0�6
b��J���@z{��oe����X�AX6��;]?��xQ�P�,��-(��N����1�����&�D1�;��z ��[g۴��	��E���n�-��J�C������Jg��v��X�=������E�^/�\���}�nBGeL9}ݞ"������~��Ч��ksn��/���ЁՋjE��*\�y�(|��n��o��Nz�G>����b��N����jqF�~cȊ��,��� -�D%�������H��?E�)+̠���2/�@�HFi�i�u�m��m�����(��mg�Q����8��5dO�i"2ٶ�{(�%�w^h�
���u�i)(_�Q5�oCG�ƙ�>���*ie�^�_#��ދ�~�C�p�p�U�Q��^��Ĩ����*^ �J�b�p�=��W�<�~�Z ���\ݞ��)�U�b��Nˁ��,J+�h k{8�GI��*C]�"΀5��A��x�>S���W�٥Ñ�m=���t�>nR�����5�x\kBT(MSr������*G�+��u)vfJѢ�*ke,���c�������~��ycKq����G"�8,���&����{'t#���/~7���]$�ʵv���e�<"kBώ�p���M���#*j���V?[	���d���w�\��2�"}��_i�cH��B�v)�מ��:A�/u�UqPC#4z�uZz��oX�DfS��Ø"F%��A{sO<�����KzPK�V��J)�1_<�:V�i����z�-�B�<Ok�a���c>�&"C�p���s5� �^>�oVh�����,�5�=Z��M�-8����#m��h��])5y��p�̜�ʐ�E.n�2\��R�4oHp^�ײ�q/���I6�̷�y���~��.�B�N��q'�Y`U�bt�2�@��8����
�/�J!��p5eoz���އ�V��®��,�['��B��|�>� �.>�e�_�eWZ���OR��� O�fA������рqya�&�,�m̚�K,�2�%��a�$�;׵�~M�� o�E<�c�p�&��9(͍M���\q�;T.o�t�{[\S$����W��x�)��ݑ��I��nǖ|�_�����k�ә��`�Z,ݘ�T�<{�l�ϝ��qښƟ# �z�{b�x��99�㲃�c����Z�-��&v�jnv~M��E�!;��k��ޙb����b(| ����靑w�m�2�x�E��g��/�Dx�J1:Y�v9����"����~����9� `���(�	^����(:�Wd�G+{i����`�+e�?�i}��q��MV�����s��a~�b��Y�&,}�Nc=�� Sz��=�1��wIF��1��[GV���?ԛ~y�G݉��;��6%�{*��Z����I��~���C� ��n��o�A�o� ���������E]�~d���o���[ao𣙬����ۍ�n�P|�X'l�d����ԥٹ��w�Z0 �Z�<W֬c���i���}�=!!�2L�ߑBOY��sP�>vln�>�àyy�O� # �/�~e�߅����S5[��8M&�8Ă]����WA�1���D�|�Y�f��U��,-�L)u�'S	eEƗ��k��^8�Mw�iՅ���4�2e(���7`�U���/�D���e���=by�����<����b���|`�X
�W>��iL=>JEҘq����#W�D�������r	~[1C����@WGm�z��n�%#������T~[��ea�N�m H��L��]h���f���RXq�Jh��PW�r�i�)�-�l ;M�3��֦)����P�=�q�䎆������"em�&�����0�_0*2b��_`z�1� y���vU��������N�olU��S32���"j
0C�mB����~�~>D/G\�iϟ�<e��#����r���m뒫�+�� �>�W�p808C������>6������Ηb%sn��� ���dC}Z��)�Ր�_vIޠ�d�|�W�:SI�;�(?��sΨ$=uW��p78[l��hF�J��;X�`ɯ|%U���,貾��fLD>t�Yp/���Y����1��HX��0,���馬�G�X�����>FY��J�#�}���nL	���ay3����A#����(�6�늀��QY��pʕ���"T9B�JX��:��J%9�R��,������v��*���6u�@"Ƽ�j�)v��~��^��uUm�kp��I���_X0hմ�����U@��#xu!ا��H�o���h���on/K����O�)�D���>�I4WB���Η�y�w�Ӳ�v~�J7!1��3(yQ���Y=��<��y�.Z�&?�"ផR�]K����
	�D��kh��TH#�<�1UA39�ͪ�!B�WГe�gq������5��&�~�q�0eLp���H�l�*�T+>��u~\擶dN�|��)Lx�2����>"�כ���޺��]
��s��%}]�\��K�^j�'�Kr"R(ML���wf�,�D��G�k��=N�؋��C�i\��P����Xi9��m�Zp�֙�3��_��m��I��Ui���l�_�׺�\�+�1��6�f8%d��	J��0�b�4@��զ�lk�e7�Έ�c|k�H��f���X�`y*��@G���hcJ�!>�2�+�|Q��� ��:�@�Gّ�$�KG��?����ʨ��w��ǣ�YA�|˵~��(N�6����	D���)�j�(��+)+���j�{/j���g�6��A3��A�*%�9`P�%�,0�
��R��D�\����@��@S?L�O�s���{0����ҋ�"|iEK~�者��'[����-jR��%��%ޫJԉ��Ԥ2�oK�ǲ���#/1J���_��Lΐ�/�m*�����&r��i�"�r|_5��8I�I6uX�tIY�0�~8
���� k��2��Quz�A4bE	�������i����*(�A��u9�F��+��a��A�����Z����6�k"��u�+���4P�����Q̸���!I���<���S%�(6)�����G�;L�JSD̾��\�)+�47�!Ǘ���Du�(pč� ���G�"�Ȓ6/����Q�F��$X��f��|m_�4�0��&�r��K����z��a�)qR!�h%|ըŐ�_$��M�2{��Ѕ �������0����2����gw�L���{�d) f��^,D�'�Wy��,TKaL?�������%��.!�dVobü�þ~�)|"�&��&�����o��6~�[F���>�������	�#�nc�	g)�3%Iu�R�0z����P�4N�D	]9u}�w���U����b�7륆nO�3��θ#��7��
���A˔�� Ъ������&��xM;s�����H�%��ίH��{.��i�<��n%-�E.�&{C�&n�ZXa+oB���L_�2���pZ��R��~��$Iw�����57Q�%�!�E�$��i>M`=nޝ��e��s�H�&Ț��L=]vK�9���#-|n��l;�x����}��K���psܭ�Ŧ�l\Dj��fE�������u7���q��7�25}�֓�A��n��`��R�p4�ե�b5uJd������k�_��]�98�H%�,����Y�a�s�z���Z�	q�F�˴�Q0	Av�_���\k�:0s��n
�E�")���O��)���{G�
�u�3��2�?�g?������n�@���25n9����k|�!��@���j�T#����d�\��I>�MC>�����G�$&�"wSRD�������ED1�*헗� ~~U�@��Fɧ���],���&���-a�TK���\��N��?�?�T��[�1�B@��|�h������;\7���S*7�/��������L�W�����y��|N�����m2��XAe)��������5#�@g����g/��R1	D���[Qv Fo8�K�*�9dҷ��.��ޘ~�0ΑpKZ1��=k���ՄqWv[�qJ��ہ���B���:A]��\��zǑџ��������*��(�H��Z�XN��\*Ƒ-�M��FQ��:!�;�ǌL�ǚ�F�Ī���1����Q1W��S�����I�7��<�bj�K]�*��E�qxU�ދrj�m�r�^"h������-.�0L���OT��)��&{��Z�����A�����s�r�� (����W�2Ι@g9���
Ck��ļ�.�j#�B�R�#�B½]�؎n��̈Y���UH#��k����0 6�=d\X�u0�C7��P�Z˒��h/x!19m;�;�Q��nm�
:�>}m��q���gr$�����VLn[�e8��;c0�|�N�:vP���p-W�P�Gx�͚
�d�I�쑶�q�b,��|�1�6����v�h�Z皰�(}����e����T�XсKA���oYv�Py �>]e��-i�'k���r�񚕷�@�kj
|�nԱ�V��n�U�Fb_X�]�;yb����K�b8c]���
��鵁�����D	���C�D�k4�rd1)341�,��n�����n�>���W��}�Ia�����%L�s���"tq��6���<f8�LB]!�[�>7��ɢY�$��I���qg/�t+m�>mr�D=@�Ȍg[C��<(�w����*��bL�!��ԹY�}
����C�N�*GE=a�_�����f�����]�q��A8�g�	��֭}�,�
m�[J1Bl`a5�i���� T6�[nJ�a��NDÞ}lDn�=�%�!>�C�j�n�5b��	ϧ#z�暯��B�ak��A\_��5�ý���_�Iϕe�;ѱqu8#,F��迾L�*�ϸ�j��ih���Sb��@4	��	>-�����4�ŉ!�;x���j�g��#��� �R���Q�]�`$
�5�f�Nf	�^jb��Ԃ��P0�\-�kwn����j��j�lLl��Eb��V�Z��U<��9HZ�ɤ��X
u��{W$fc�!�X6}����d�H�	H<� -��sO
� �/�N�����r@���.=�.��hUyG�A��"��W��R�!���abL,FzBN�W��"7�8=#�T�T8n����:�Jj�n�Y��J5�FRI�"�h"�ꫛ�M6�d��U���q�Ȅ�$Ā6"v�0�����Fhz[pYb��M�G=���nǑa'BT7f5�ۼ��4X(''�ȯ0uµ�-x#�iR��И��Vjǆ�;t�MZ�L8Q�ME[��)b�	9��8�n��E{K1)2�S��\1��j���WJ����=�
����8��T��rL�5� �9�N|���sh��d�*�z�	S_^���\��Ok�\g$=`�� �4��L�K��6��'z%a�5�9�>���ExM���hC2�����xpj����m�dop��l�{�.�_��m�]K;�S�}�U[�4n��3xL�-��A�JL��R��6o������y�ބ�D�e"��k�I��CORQ�[g�*م ��̸�����u�r��;�7�7��"�'�l��?e�(�����O[�岏z���c:u�Njfi�
�wܸ��=�JEV_�%�!���	{���>�O����m���+QsL�d��5��Pi>�:���L��OvVQu���a�a|��d�Z`ig���=dOn���.t�����@1[�����V�9d�ts~;��9+�����
^G"���k����j�#�!���ٯx�/��Ƈ����p���/��Y��b� ��7�T(�sr=�"�u$���X���	��7��ϵR��>�e�U���$�n���8���f��vP=ͭ��u�&������,���D���oН[����-����J��{L~d��\�(�@�mO���X�	�6&���q؟���'P�ެz"�#pob�Ԣ���9���n���M[��C����������]�#x.����@�� ¸1�"��+E	���u��b����`m>�b��
t�yo�c�F�A��ņ��g8M��ϥ|��F&�T�9�a٬��x�?�Q;,�Ӻ�e���}\O��Vu�1���$�����Rk3��H96���ldK����{=`{@l��������ȼC������v��k���؞3�d
?6���`^��
P�-�M4��1��� �����)wW�0�̥��W��9Se�3�)yK�3��Ӂ�UY%�#qF��~6$�ޜ�Y�	��O�� JjJ�-����\�+�s��ipz�QLć�(��U�Ճ���>q�R�4�&��+����*D�Q���6����(M��VV�P�����f-9�Ze�fL!�2*.�'{f�;�E���U�Da���߂��L$1�H"�`���M�n;�G.MWm������)6�.��,��X9�8�43	�t�&����FVfE'Ϥk=Ӫ���^�����<g�#�ֿ1��%��d���l�`�+�͛�v�$,��ip{�j��po z���.��Z�� i�*�$/6�\��5��k�{�Sf��4�%�8��B��վ�[6-ԋ��m�N���_�b�6���a�P�~��yi�5JL�k�I�k�*P��l�ڙ۶��0��W�/O��,���U><�il��7Z�̓���Y��i�P��i$� �U���X�AP2h��j�`���	W����O_�o����Ö�-���K֯�aGv�]���o9���R������t�.֝_��,#�򃴈I�SK�|��w��r�q�B7�]Z��L�_�#�/��`�_���rAӾ�V����͹�j�g�v��*���:"	����iG]ӯʮ��Ō�F��bo��h�2y4�h�W�d����!�J1YD��^�Z�db���+9���9��4�P��ɒOl� ށ54�G��Ƨ�#X��c���?�e�"����-��p2��UD�o{�ct�Y5��3��tY^�̙�>�?������N��+�|=�����H�ZWrhFxT�|��fe�Ԑ��X/�N�XY�pF���!��3p�� �^a�uZ%�ڧ��wh��~y)`,�����lg�?�#�Ĥ���O3�8o�h4��p}����8�M�!� �S[�r��Bf
�Hv]�J��aЉ+!-�{p�g ޮ�E0��Z��z��.x�ױC��u.|�g�5�Lȴz�

+i�Z��������7�����Y�}n�<�}4ު��N��<�r�E�]��%�|{��u��B>��2gj>�s f�)�.���dO��lu�����g'sP�史�UX�rxEؗT��z��['�@_H��-�G���֑����]&j�>�k~tw�F���g��tjí�$B��,O���P49���+����;Cw:�)��r�J4{�}�.Oo�R?<�?�a��I����R�U����T�H�cPn�ӑQx0����K�/L���AєlѴ�뜟����l��'I��W�����"�L,v�*�7����֖г��s&&X�!f�;�%���R�+1o��N��1��5.[U�[��kg)�oH�e�_3h�}�џ�6����yX�S-��x�~ܥ��E,e+����!&�z�gI��5L3/U��I��(�̣�N֍�K�S�
wc�8S�5���W�hNv�Z�=;��7:��VA{����X�w�/\�3Q����ʲ8�gZ��{H���@�@�>��]��+�D����v������۽�kI�C�L5eD�����}�1���j���Ʃ���ל9~9-�$�O���d��!m[t9s�n�`~��3I��� \��������My�3�Zh2�\�̉97h���+�B�� ��qĞ�)nS�)�Q�a�
���$�v� 	^ 6�VM��QK5"��zJV�'N$~`[m�D���gq�J;�rŴ_�c�O�?������������3��x��J�c�c���]���	����훞dX��wV�ܰ�G�C@	��ߤ���a���rd��>:$(��"��֢g�p��Ad���:=A�� �f~�P;r��-Ć��+q��ck\,���7����;�?(�׆3�'8H����̷��|%!��zx�l���	�3Gy$���u[��ʆS�<"��ḵ̓G�/�9�����k QZ����n*�\g�����3\�K�,���6븲�/��\�J��8)�T�lq��3�Y�n�+��)9��.HK-{����]#˒>��&(��Z��ۍG�0�j1h�=�u�i��� j�������Z��`��(�0�6�e)��¢��;96�������/_�yw�f�Jx�]�N��廔���F�r�*�)e�@굏��P;�t�e2�L�㑚XB�e�d�(0t��u���i4�3�$~�?Ub���.ݞ��M얧>L{�L7e��j^谍d-�� �ܝG�d�&ϝ�
e��ysm�d~����&#?���d(]8;F%�JG�Y�^�z��j)�u$'�"��ǟ-�l�W�@ݵ`v��'+�,�O�:���w��fX�I�����~�8	������^�ÿ�qG{����}�bJ;�)S#�p��⛺owfcs/���.�%Y��ko�o��Ɖ�dL����/�Mױ�Q\6�/�UC�C<�-ԍ�K֣Z�,���G*L
I�7a�uF�M۰�h/�v��9e��2����8	��F�L`���Ω�����Ə���V�h(-��C35�WF.+���y�`���*+o?�䐚�?t}a�s!��t��m"�qeN���ڬ���R+�ɒn�EHn�z��*�����~�p51V!e7D�:9,�*���[�:�:A��I�e[9���i1k�|�,��<S�	U�G�;��C���lN4�rO w%G��#���r1ʵ�=�Eҙ=�3f$��溿2��[��~6��4��B�Y�Rn|��:����B�T.�8���j�'�3�;�f�k���T�{��R� ���l��0n�87d��dŝ�Q�����⎐�
�M��̲��ME`��#uhYx����A`Saܱ�KF�t��Ɉ�))k<�ɥ�P۷��<�����J���4���B-G(I��W�/����?�S��RC���'<���k��4%�9�J�B���{3pQ�V�h=��p�¶����;�ccT'�yn�]w���f�|c��B�p��hN�h/2��Ǔ�a��ۚ^s��@sL�
X9�Ox��/��C�Onư*�6ԛN�B��M��kASK�H�=	��Չ�Ζ��"5�^X=3h1����}"1����ԩ�_�'R���DQ��z�� �~���릈@u�Ύ��a �I�%�[�8Hy=J��l�g�#e�ZF�9;���qX�$:��I��������/����Q$�!�A���0�_z��G�y����D�H/�t�S51���)�7�6��uq���S���̷����.QX����+N����4�yT��AKZ�>�Bj"�v�l`P�eJ�����4y:Ь�7��͸�֛����!d�zv	fWt8&�����&�����Y�,��1	���ɬ*�Z�au��3��l��������'��s.��6@X�g��&���/�9�dl�ڙY�C��B}������;'��I��S����_�q|�ԅ���wl�&�9? R)�/܍_"CC����$�_ψ��K��5|		�R���683���7$��l�	��-P����Q��W��K��~	_� 0��<�O���d��� ���s�
�řP҈QoWp��^�� shS�]2$�|�����SB�H6���X6`1&�б����=�<!���[Wx���
�RÜ"���|'�W�FAM�o�r.�u��x�T	%iG+6��i@q��e�FT���;:�����Ȉ�p�O�ު ��E��ۍzV!�lJ�vR�^)<��-�\q�P_As����}6-�괄�������,�B�M�\[�E��=R-����z էy���5����d_��nJ��{,N������ܶ����N�.����^gL�3{-#�'�ۚA��j�	7�R��S��vW/~�Zm