��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\���V�fnvx��ÍG_;�ȅe�~�>���9�>��Y;�0G��g��;W&F�_�8! �%��VGsL=��ٯ}���"�CY��,26� k`Jƣ���W�A;��tk ��s-.��K�s���Ux�g.!zQz~��d��P�Xm$����m��u<�冔_ �iUc�gK&h���q��]�0՚�J?+N���G���)/�zK�O�!=�(�%��019^_���M&��Sg����˥�qK��z@� �ڻ-v@��M�cY�/�M�Ҙ���-]�/2�UP@}&��������|���k�9+��MD��C��o�9�P��	���U/�TJZK��H�EJ��i�a2Q���,P�$9� �-l��.�Ɔ��r�m�+pף��bQbm#�?y�3�d����{�j�~���aJ�Ž��I�/򻁻�F�C�62�h�O��O"���x8�����2Ħܾ�?����!X�1�ݘ�T݉�Iz��2��D��P�6��#��L�7/w�u���pT�\rZՀ��
��g��}b��R�]_���������)�$^��S��u�6DQN�S���~�Eq���,�<B^H�6��4�Z�ȱaY/ّ�j|9�U8g<�9l�nd�s���h�@aT�ӟ<4�Ӟ_�*)(��B��8t��s�=b�#�u֑R?�P'�7�q�����(cfw����L4��3���a��*���~6ߵ��wG|��P���R��$ig�}���q�G��,,b�ĸ��
4د�-�4������G
�aĹ�+>�S���v�yi u{�Mp?nx��[�(a�����@{���I�$���w��?�'z5�טC��*�G���J�*;ltKh��O4�-yA'.�����8/�a�;���(q���k��Y�u�u��aթ)☋&2���Ͷ3�oxȖv��@�[�0���7N�^�L=�U���0�_�8l��Q�c���Nj�g̠X�^�4� �����KY!�6�(��~�X���ICR8U���L�+�
�_0��dBK^�����R-X�]F?;ү��K���y[�sB�<JZ�=x�"��.��I������ߧʂmAW!�k���{b�
�e�Y<Y�
�o�@?�J�P�C�#r'A���IC�6Tv����=�� yn
7=&ǽ2��B k^�iL���|�)���@���]Z���r�?jF?�M�m���Cv���$-��ۺ�2pΒK�^s�t<��m-���ZW����
zV�'u�o��d1SV�@)s3ܩ;Q̤��<��O���W���ة�R>.��Id|���u糶�L(�#���xT���ǥ}���%��(��*�23� �ni`�bo"t^����j��u���"�^9�1�7�e�H3H�d��x��>`�&w�k��q){w�*�]έ� ������w���Jڋg�(��џ�0r+�������aN����`��c:���G�ޗh����
�``K�Jk�h��&8�]n-O]�g�\M֧'op�1�
ǉᐡ�>�!!���'u���]�*Ԋc�+z{�xQ�N��� ϕJ㻂�2�C�b�[.�}?�S{�BC?�Ma�kH{ڙqu�, !�5�p�075��}�i��FSs�5ݨ�3�/���N�$a�l!*�\��ɲ+L��<�߷�V̿#�,����.�Ǚ� gd�����(��� ��dP-�F!����W₤
_�3�v�r��?�Uei��;�w��fhC�u�I��q�c���d_X��}�a�����t^���2������\�/��3�>��9��YͣMO���*QF�9{�ᴡ�Z��~��c7:�̿+3nQ;v��Sr%y����u����<1�fu��lK&e+.�!w~�σp���aK(A�إ������2����Rj��u��c�+Y��unl��^1�y��������Ӡ��~z��ĵ͝�����nߦhU�]F�^������D��N�1=�$�%"�{g�?Z���Z��e��0�܉`r���o�{`l�G�<Y�&gHԇ�[?����kK=��2��?@���!]�a��ו�m��Z��.Gd����|-HȠp�@�xSwy�Z�B�K�=IFF�j��Q��A�ڥw���'�R	Ü˂V�=�u���D����T�5�[sc������*S���@y��M�*i�8F~ex�����a �;�v1D��͹<�9�M{gD�Հ�җ�E���x�;e��U��Sm��v�ܰ e�	����~}�>���¼�a�>ы腏HEVu(f�#�K���#=�ץVgک?̽��Vw��f������^
��n���,���S�nH�W{�tXQ��qC7��5j�RXI��/�����*��x`O�:�3��2z�➚p���%}�4��sT1P���4�3E��UV͗U��\vR]�	���VAD��2�-�j��By�|G��Un�l4A�!��|>����aXO��6��` g*H�L�@:w3�sg�����@��� ����6��eEA�%�= y�:�?dF<�5�DГ��t�ʵCO��-����"u�*2�k�c��P�r(XDk3�?�N��0]h$
o},��9#�n#��Y��5��:XxU����%��aXޢ�?�W�w��,��ޭ�������kA���rXX�2;�F��m�"q�?9]���l��ȌZ�Y�4����.)�/�<�i15���3�WJ��@D�.3ߙ|
6�Wm�����/�wvN8>���\_bGqtE�bOyy��{IF�m��=�B��\<<Ij<��y���B|�b��c��[)�:hb5����r�"Kׁ�}���,��*a
�霴�>D�g�
We"�v�>�Q]�2x��<%��{�tL�W����S�j�i��\�i8ޢ9�����oz��8��O�N�h����٫�TC��7g
G$rj�r���������z&D�1_�N�T����',���L�?D0��2m��Z7=��i]GRH�\���u粋�6!J.C���8ϵ˭��S�Q�$�ۥ�r�R��	�B
��1�V�A�ZǟN��^L���K(E%2���ER6��^�D��  Rh'�ͫ[h#T�� ���Qյ��#j�Z���\z��4�5n�E���܂S܊����n�E���@Y��A�1