��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>>�Htd�	5w��O�� ��dE�O�95,'��d	���aa�~��Zbr־�Xg���_�د�obu�Z?%�MP��������s��O�o��l:�a�o��
���O��HU�ڍ�w��o���.���i{�����VZ�+� ���M;i��R窑� o��9���	�HIH���$6��m�4�8���O�©�d8)�� ȧ���Z�s�&�q�Su��;��]�W~���Υ��E	vf�Zq��koɹ^� g��y�g:�:� ���6چH�66����O%}���nÕE�`+J+9&� YذK}��K�]�D�Ci��鉭�Dq���i�{�w[>	�S+�*4���DKB �]"�t:��ܙE���c &�-n��3
5����ܑb�s5u0}'oSc(�$^�Ѫ'��S�az��$�?�<žf���;��n�S*�=���y&G���N�,U����S ���|�q�P�m�'��7z�nf0�+/�(��F�����,4І ;z�" ��"����  Ash������x�h��[w'�D\ē��w(�����~�k�}P}�`kO�~}u0ZH�y��4�X�ya�b�ƒ���c$+�0�L�1ŕ�#"2o�({�M*ŜU���p��y\C���1=�(%��,(OSIp�2
�o"���]nU��������e�)� ��g��֔����'L���gs2q_7n���Nh���5C�\i2�l�ʾ�jHc�q�^Q��@��
I�Y��a)�;^��4���X	$��w��Z��3��D�-����i� ��MW&���6����b�挼V�kĜc�ܵ�x=N�ΈI��0�32j1y��|ҭ�0 �2�^8z3��g��(,!!�L��i5Qy������6���B�ӛůo�.T�ӳQ٧�#b�b��(����J�4��Q	c(�#ϊ|{]J��)�Q/��Z��NjaX=���F����I�Bk!(��[�|$j$N�4�O;��5�A藟�vXw���Y�POK��B~4�hD��z�1�]'���(:�xb�Nafq�d�����[T(!�y��\=�Qon[�O(M�ې�S�1!��z1~��9?i R�4�be�q�]	U���!�+z�ެ�u:�%�?_�G����Wk-o�S7|k��Lw�_�1g�`X�dE�9��ik���P��X����u���a@��a)'���f��#k8&���)8�0�	+����k�Hc��C��t+���
�2 �+ƾ_2Z�~�������Pl�y�UN�p�Gq�ǖ%�S/��CѩU�$5�pm�'���X�:�-bn���@���w`T�����"T	J��2�m*`��.�o�]5<�U��!���{�z�V7�1�""D�kf �w���M�U���Pl���>��P��-�CJr
�>�}��
J@��f"�l�Db��%b��l�O|���R�݊�y���oS���[��O��~d�nN���0�C怒���e�%�T�`����3�w�#���VW��a���.���[U��KA�p��R��_׸2$��_�]
ev����EÖ�$g{�S�RV���&q��(oeB^�[��*K�	G�\�b���l�c�{On��~�y&|匌�5���*��s��#sf�'*Ǐ�;tvpOo���+j5oz_s�։�0>�#㛳�ї��xS��S<aYq�����h(�͙lb÷��6�Z��EJ�i	�v��2Xi^��h�FB�.#�a_EE#bT��Vٲ������hg�` \��^`9� �˞��X��Ϩ
މ��d�0��}yLO;�r�U��ۚq�Z����i�#�-��YY#@�]	��Iy1l�:֜<ɔO[�- �.C@�U<�(ZT�9�*1h��$h�s�lG�W�E�9:r�o���֒R�L�t3�n�2|�-+�
�-R�����5\��n��7�)�����s�VS����cV��\u��I�qbK[A;o���r!~fE53�}��UaF�"K�	�h�g�����l��0��/�b1��в*��m:'��H��	�����cCyLCs�`Z����_�rmB��N!ϼ���P3ƿ���g��Vw+H��Ϯ�A�"�U���:7�}���xk�.2����ed"�
n�����M�2V����'"
�p����x�|�g�Շ��O�\�lQ��EaK��8)���g�Ʌ��x/��*��Wo칶����Og��z�-�>>�[q9�t��Kz@"3t�Qnͽ����M��Qn8�hZ����x0Ѿ�Q�X����b_��ME�<��-ay�6�����f�
�¡��=�vU�h�J����Q%���J�#��o7���7�W��?�����R��]�R�Lt^F���Gh��zj���������B����͡��F��ϑ�:Ymh]����7$��C�wu�NA�d��oѮ7!��u�!(\��,�B�|EN�-���`}OTt��߬�BSD�HQB
�nXt.��,dX��`t��1_`u��k' N\�O|X_焧i�E�R���t���i�J��k�AGC�
�X�s�}�0n���x��쳟H�0��v֯r|ٽ��w��
VwNH����D���Muc�*�H�d���k������'ݨ�*,l�E��K#�F�?��"\�`�f�OZ��>f����.�zcL�K�|e�����P��c�YRF����
 �{��l���ϸ٥�b�I�w3%�fv�F��#u�����sf��<�7,���n�l�����d�,��Fj�[�		*��֠� m'�I�D�*SX�P�)}�Cc2�W�3��Y��>�5S���cR��2���R��6��F����߼b��6��0�%���.gH4#�+��3���K�i�>�ǐҰ�]Mn�'���=M���bx9�F�ឱX,�e<b�ޖmeR�Y}���[ S�%k��!'�<�b�,Z,��FCp�=�B�M�/)p�>g\31�~����&�Ķ�2�O��Y��$�F"E�v]��7�H���7sLj��
�<��qy�ʍ[�[����2I>�y��[�[y�'c�Oޜ:��x:s~�i1�x�!=J�qi��+�Ug�Ǡn�X�-(��������T�B؂VJb��+TA�!�.{���h�?cʑӸ�s䧏�U�c��g��;��W+U����6{q}�I=��|
�U��a�̈Zj3գ�ΧY��_�／�[&�!� ��I|���E7b�}
�˖Q����$�����z����m4o_�%R1�"BZ��p�� 07kC�zĒo@yhV �tsl6W���|͓o�+��g�