��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�i��a
Α1S%� �uj?�L�3��TLei-3^5]E�$���e5r(��+�uG������{�����]�M]ۘh���/�ob�`e*���yy�i�������
�u���q0:�./o؎+ՠ�J2~E�2�r¯�h?y��k�c-Wy�EDS�(�<�jrV�`��'�mb�b�ݤL`4�Ԟx��{�B�I�f��̄VGX�nbeD]�ڴ��L5i�	�+�3���r祏�j�ʂ-�9��h���CA �˸uWa�-j\�ӂ[��^�d��'D���ج�Т9�9�~���j]M�}Ѵ�T��b���̶{�Nm�DI� �?�����A���?�m��[��K���Ǆ,��ᗥ�Ux0�������k�U�Q�πQ��L�m��^0�ќ�^��m3n:͢���B�Q���O>Ԁ�$�+�19;��~֬��X� ��KT�4J4*IfR�/qz�:�?���X��1���|7l�=Y��V��	��^f�w ����̫\mC.j�/ML�mZ�cճ�~�_Jh9��O(*���cw:8���>M�U���c͐D^o1��ԏ��rMB7N��XO��̯h����YT�ο�"�!<�O׈�2��`���]�����7��}�]A+���.9cͪ�a�&�x=�C���F.$�	���-�Uv!
,�{��I�T7��;j���wqH��h��y��b������)��Q�]�QY"�ΤD3r��f���VjB9<��L\I�3�mG����2W��"�9v��h0�5���J��kF��S Z	����V�e]�(W�=�f�T�����g'G֖%2k��\3�S
��g��X���]��G��8�T:!�Qi��h��NĬ4��l��}�"Y�u�'�񱜈� %�O�7-��y�\�pcYFl�6��*��0ft#jo9�=P: ���#�~�{��w��R���'�m��`�Q �%݀Q��ѽl�1b^A9��>7-r?6g�:��r����V�}M�=?� .'�xK�*��i��@�o�S6�O�Z^�@�dϧ*p��2���W�U��G�4p���ip�����MZ�d��/��u������`����=��VS4:�硶�8%[��{��j���^V>�y?���S�[Ԑ�=�b�Ge�6(]�/��1D]�Ģ�4Vr'���R!�{j�SY�����>\���#H`�����u D�R�#Ia �"Y|�> ŻHڒ�q$�>�n+ٹ�v��e��J˴�Qg�nt��e�g�YDD�7y��dE0=�c\B��%�C���A@Qd�+�
EvQ��\��c���f�U~X����Φ�V��?t��Ĉ_9T�"�,��݇{OȁR?į�T9��ژ���q��ߙ��Z,`��	���^���B;%�I�}o���s�t8�V��׌�p����-Uo�'��eAfYNa���vC��/�Y/>�4��L]8��Z���➵�9P�F��c�FZ�ezЎ9D��ծ�I�"4�z���Y�Y��.�f]��4����B�'˾����)}�@	��4zj*�,������LΠu׆*4 "��R=}��8��d,Y�),� M�+Ș��\��?�&�7Qe����󙦶���7�\=�������X���9����j��=��r���l���w���z�q�;�sa?>� �D����5.�5�nnݗ �"4��4��z�o�tJ��&!5�n��.�6qf�Z��O�Z��/�V�L>�٧^�z�d�M�����fQb�{FE'��X�A�#�l�PCn��#�X�"��s
�������7@+���0�$y8��2c��F�Q�A�ɐ��9�'{��~ʓx�}&13D��O\�=��]�����5��ui��Ձ:������0Rj�9
��`'z;��+��#δQ�p��t���S�{���]y�����˪�σ�l�{��U��Z�t唰S��.SݞY�o�L�}&�f:|R�«�o�0b�Ǣ=JD"C���?��q��zR�ȥ	��J`�I�ꡟs(���������e�����I�K��?�J�@0#B��c��wt;�o||ː�n/Ji��["H�=Yzt0A~ ��٢���J9��/iO�
ރ�;���ʄ����
g(�Ш��_|�˾1c6��v�ɬb��_�~�\ 4Rڭe�QRi�B!��2�&��l�r-q�W�|q�*O�	R�oiU��ڨ�)��6 JfS�l��s1}@��E�%lkIY�QU~�n_'��|X9��a�҆=��O����I�/S���4���46��)�A���`��׿ D&n�k���ۢ�FylF*�0t1�Pֿ�}���[��[,D�%%�U��y�Z\J�����>� T7�ӑ��Fq;���T��zFA��!u>�OP#|�b��g��s^))0G�l��xmj���k�ZC��3�z���1�j.�]���Ջ=�D�Q7�q=#�qf�@��s�7��Q���(����Ib��B��ָ_D���{�D�V�{���;p*0R�wz��>¥��]L�о�s�h�%Z�eui(���T���Hú���zk�ƮU]v:6�O�{^�Г��5���m��k���y�	dT���~��Pd�8͎k4��_I]VUT��������P���E{�b�/y���q�bD���H��m�BK=�Ú��&�2�-Dg��R������	rU D��:�$�}��"�_��c�X&��o3�\<�x�4Eg�2&9���߂)�j�D�U^#�R����a� ���\�g9���[����Aב�Rq�P8���3���]�=I�e���,�1���T{��R�]�B~�Db���=c)��$�����~x�s���b�f�U�W;�������ˢ�Zs�Y6���¼9២ї��s3*�
<���ժ?���I1�t����J�I4��-��莎�z(�{�0�@��'��S���)g��������Hg�!����<�Ʋhr&��ҹ�N�["P*}��VIS�3kz�ّ8W���eDK��3��[8�a6��E�$ƌ��X_�l]��-4DJG�X}��;�_�&�%�]+XS�p��H�z^���_�/�@�úU���Z�>N4��s���OÈ�E_%g;����D���P�PA^=��N��:�'1���QzV{L�[Z�<�/�㬆1�E����/�� !G4_3���f>Ԏ4��(A�E-6���å�{�k���Ka�\su���+FC0���ˀ�:Jz���k�f��6PN�z���vC{暑Z",�Tԫ�F�<O�W��Wk���h��%�RM���x���m��ו{�{�.sD�҂E���S��6L_W">�`U�����ă�8�	��D�wV=��a��)��P/��/��>���	M�2�M�w���ݳk�ޫ��v�o����Zw�^/�����!���_y�i���s�&U\]�@j+i^�	�0H�8��^��	��o���P8�U�'��u�~a�冽^�&�E��sd;g�J8u����c�ˢU�5�=Cʢ?�sy��I�n�}ξ���c�����!�^��揷`>��J��@�<g�Xw�YOXqKC�	�{��J=�1����׀�U[~��=����Ő_��ƌ��I�Ym�ݲh�
=�?��(��`��pW�]��cˬ�Kz��F /L%�hU��X2����%m1S�J�3�N�C�W��OO&��/�.V8d@��^��W D_mI|uOᐷ��F��A��S_C��k�'�Q���j�dS��~�n���.��ߐ'�7���L�ق��Pn\�M�~;^�ɜ����嗍���35���x��4�NX��˨w���Pv��x�kJG4�(� �&�8N�l����_�o��k���J�TT��mӛǜ���,H�'H�]�<�܏$��.v~m��*��0�م���y���6䏶���C'�m�E�Qz8���f,s��%]�;6�}��֏CaR�x�����DX��ͽrq�������� V��c�|�g[kMh+0��D�����s�h�HV?9�q
N�L��#�iu�v��>�$�VkX��4�O���� yxOUzy�N�Ʊ�/����'U,�6D�O��ZI(�ن|yr�ģ�zꪓ�ڇO&��B3J���;�>Qr���P�9F�l�V_�A�equq����tq����U�mL�Y��kt-����ǥ�����WfTp�f�u�-��7=�2�&�@U ������T�c������b:�S#R��,��@���Rz�<ղ���baDUd���Y��C����D��.f��*��xe��9o��JdB<n_�uI	)d�iL���z��;n�i1P�a�}�F-15���(��$�UN����Q�9����*@����r̺ә�k���k������O��,N1U�1�PK��T$��mM��S��MG8�߆4�S�t�r1��@E0�c�t-B!�Nq:�Un�Pt�9���^�������IP�gc�� ,i��eA/�h��|��#�a�B���#�C�2v��^��Xc��!���n}��_'����#��c
���s��%��Ǣ��8[�zh��ݘ�߄�;�E�u��o�щ�BW$������)��t4��n���3	Ɯ�HKԢ�ѤB�M�8�I� % `r�v��^�#O���T݁P�Vf�8�[G��#͸֤w 3�[�-0�9_V�2)jF���\�3����*4���z��)�w��9��).��2�ރ����`�)(+�A������ثlWܖ�z�jY@@��p��`�a�^�J�nϤzND��y�i��Mj��7�*x��c�)�.u�Mq��T�������R���Y.�䗑�cB�+�(-@�q*M:��R�fE���]���@�*?M��7B�,�l��~>6��)!�Ys�\4͋�b��Hg��yO��n[ۺ\���L�����{j!���)5ő2VE߁e&Lo�������h��%� ��P�h�&��!�H� ~!SȜ�J���,�N�Q�q�Z�.�R��x�v��G�/�S�^���"_>l%�[�[�&j�c�)�h.�k�ۼpffę�V����ͽ�~*g�����'i-ݰEp�ڂ�غ�S9��|��~|%�U�(gj�(�02K���		/	��+���ɳ�؈ڿ,?6=�T]�w�]9�9��!����mǃh07p��
�7���I�0 *47��^��1r`pP8�R����"8v&D�n�G ���d7���F)��(t*f��%��
q����H����}B7L��Y\05>� �[�%"���afP9._�s{�٭��ꫴ�s!��=���z�/�n�4�n��%��nB��]w�/��ݭ_�ɉh��`��E�jz`M�~3ٸL��yX�,塨M�N>���7�ql��x�=В3����X�6N܃�o~��?�b" �}��>�Z4���)��Vg��Ф�ar�/�@1<B!��4<�t'�^G!�� Z��q�H"����ni��~���̺Y����E��E�k��~@�<Sh"��}:&.NIr$�����-vؐIsj�����_��Z�v�b!��;i_iэ�
+j������)�(�iAs�z��Ua�j�"�C��C:l!+3��I�D
�@�h�*z�wy�:B��W�����X���ݹN��Ն��}��m@�뾠n�ݟ�)�7��G�w�~U�,��-͢@�t�m�z�]ȓ���.]a/L9�%�PVR��&V+Α�d=��Y�(/���"��|r"�:ᙴ
ȇ���f��	�<�~��4pA6	GJ��V�h��l���]��)��͚�5�.�V^��C�İ�۟�_e)�>(c�z(��w$F���d5���K>� ����?���E)�o�t	;�|jr�:�?�����fHhx�� ����"����w�x�ҩ
X�^h �-�G1����/reQ7S&�<i�{�9����J����:�Q��_d���lU$�P�s�0���[���4Ѩ���>�e8/UR�I|�I�����6�d�v�2�DZBe[�L�c��Tϗ542ȇ8�fa�tq�߻P���r�t���J����Z\Z�{�\���X��c��X�*����\d��?��@/`��[���w�L+ߧ���w�4��*/�ÍD�p�$]��BQ�Ѵb�I2����Ǩ��SEP'�~�����dZC
����,U����7�o	͹��g;�{Yc�<;�nǔ/-�P�,�<j�a�I�NJمm ��;*
U��48<���D<k�\���l)0�����霄}�w~�_��{3�1��tuG�kT�͆[:��V@`�Hҙ�3XNTR	G"��x:6���}����&\�Ϋ�~�,����X�1��w9H,+��)�Eט/�`j��,{ͨ�ھ7�JN��,SLqD��u��<O���wD�dk��>W�H��%M�v���	cV,�Qz	�U���岅���ւ��r��)Ix�:,�P�ey�z/��� �=Bn�׼4U���7��
!���P���	M��G+``�M����ǠAwq4��AU�wX��Wf&0��.ST�eix�@��@�bd������ w�)��h�D��bH0��(]�qq���8�;x����k)*c1���b�O��	[,|�#8��_OV0�����Gte���_�n�l���l1�!�1'F8��i������:������U��Z�g�n%{�	��u�
G��<I���Y��H�9gĹ)�2�b��iU�������)�^A��J�*գ�e�r"�L����b�:k&�u����R%�f�ӳB?;L�2J�8��dB���R�\V9~���n����R�c����,�ޤ�я��5>�����3���w}�2�@)��D�?ݸPq���6`�^�Yf�7-2M�U@<�|�It�D�Y�Ǌ�v��V�;3$3��-�7�I�!Lb��٫�8]�3���1d����]�uEў!��`R�Ǡ�Ҫ�%�v�x�3FH� �
G~}3�Cb��M�ӧo�C����BPq�31\�L$vk~(���i�05_-U�6kl�����>���Л#t<���+k'�L�u�M�?֚�����9Dq�O�G&a��|�F�"�R�kt���R�B�)����&-h�hs�OH�ǳO�9i|(3��-�Ƶ�K��[9�8!j����-�e��൹�r�/�|�R�ς���b���C�Op�E���Z���o�G�x��a�R����Ս����������V������X�WQ;m!������&����&ZҒpu���m͌j���!�7n������v��n�6��>n_��?בx��:�5n���U�q�aގ�U+Ҷ�r/S�[�^�~e�D9:��RL�f	��">�*b:�o|���k�}[Ļ[^�Gk���!�[�te����CZ��M��jڭD"��U=	�G4�J^2kt��ʺ%�l�I�+'�s�;f��� ���*PGUIjR�A�� B;O$��,�m�����?�a�2�����ؗ�L�`!\�qc��-��'I�|���sZ������Z-Q�q�`���DO��)]�gv�1��sUO=[-��t�vNԙ�~c)�潮`�ruol���8ˋR��"�7��/�����������E�ex[C,x��']�^x�[���6�QIn��K`Ԟe�k��[��[}������*HǷqޡe0C����)��ei����O����[��z�拗4��,)۞E4�/Q�����CR��\��ðe�_)U�7�a�zk>tpNֺKl;7�j�3��x�&Z4_'���nt�`��?F�uD/��7G��J��ݡ���$��J[���{�#<!H�\�~
;7l�ZBM�-�� ��A�Q�	^��KMWkjN��ī 	.�+9_�j�u,�H��������.W���c�ӿ�4���p�y��N�bjΒ�_�GZ��MaC�� wPW�+%�;߱��U{��*�B��2�!E�Z��R��vǒ6:�^@�#�!��;�N �ċ���3=�����,�\�}3Q�a���0�e�w�4F�6���#���@��&��Vb���E&����*s��-*�lT@I|> Ĩ���������Kʪ&�
���A���;hp7!���UJ�$�m�b�)]���l�(� �?�x�7SG޹޴�0�������*^ڏ΋�/[1@�-sF �Nu!�g)1�F�)ǐ�b���&�a���4�>�_�:9���Y�����y��Qc�&�g�$zr�l�x9�4�ej���翗���V����P�y�e�u4 |
xݤ�a9r_��U�[�I��2{�-Iii�{ϻ�q��qh�J*�tonJ����Y��Gu@P��f�Mh��!��e��M��Ť�&9Q死p�N�CtE�hA1�r�P��Ns��2��i:����A�ո���g�7��r��>��Os�$���~�zs�Z�|F�a�և��8\���Q���E��#栥��o�.��{�'�����s}�#�ܮA�IXp��M�Q���9�q���E(��z�@��j�s���R��K����pHS�4\A���Q�V骬W#R?� �!\���WJ��3w�z�We�Fs�� ���/�~L24g!���m�<:��y�7�^k7��LZ�!���i!��c�[y�����[
�|�!�(�\/��*�����T{v�\�EyB*�0��1+�,�w��	�&%�o�AЃ0}Y��u-R-�O?�-������:7!��zo�-��������x�P���j�v��2Z���������eɳ��dA���vjb��Wgm�F��!G�\�m��@��[�jQ���ѡ��Y�"����,�Y�>����d����ҏ��ҕ_�65�rĕ�4�?D����YW��wx�N����W�nOM<��8.0�5 (��⠝D0������ӑs�'Q�w��}�$�e�a�$f�p?�D�1�@I�����|cK�ܷ�=&�C��މ�Z_����rn���#ZD�xa *w��f-�|\���X���6��:,P= b�%$�8?�1P�׍�f��Q^��o����C������3`:\B���*{�o	��&��7���M5���4�P��wOPY����;�bR�GI���Po����-5��$}V��-��3��C"*,����Ci'�p�aR۾,����1���6����d�r��|w��b��(����m	�/��+�6 ��R���y-�D�l؛����1���.t�Ԃ�n*�}���kB�/��>����U
v�$J뮞"�-��Ɯ�]g��x\�^�,�K�`��z���wl�����i��J�=�z��R�߷\� �==���r̳��P.ZK�]��X�JB��K�������U��m�g�ɶ�c�E��3��=�����������A���$�2k+���B���a���*�	��"PDA�f"������ז��M���b�ʉ7��&,����#��r�k�O�Y�;���8�\a\��V�'�g���rq�tq�<���Pk8���cǰs�#,lC���AVZ�����4xm�I�[���s�����\�4����:�����'���}��*���^�\� ���o�E�*%�Ѣk�b�K�\$�̚a�� �_��Jppߝ�(oe��mG��3'q3��H�����Y؜&����s�Dh�R�(��#�n�P�|�T���[��t��� )v�cu��h�* x���QoY-Wgb8�%�7!⾃��
7�^g�d`LzS4�!)
�vX���۷;��v��NR��7�Heݡ{����/��Ot (���P8>��C�|`����M��޴�mM%n:4NI^!^�U⼔n^��t@0�@�|-��W���dq�I�������.�q�����?��NA���evD���/:��~b��JؘS�lI��L܉+�l��A͏��Q��Al�B~p���h�c]�N����Ozd. Q���Q4���ym���1<�W� V�y��Nl����?ܪ�������6\^�Y ��
l��঻���w���͚�O4����h@F��qFA���K��M�.�����߁e+|"���x+FhD�BJݩ�H�Ͼ��2�՜���_5&�@o�Ux\���k�|[o����#;'�Q*/J����Elr��
��V�ZT�~i���w��c���̎z��Q�hMu����Gc�tUB���0e��}v�w�طV�j�L��q�(�>�^`��� ��Vެ3����e�!�c�Z�I�.m?r�l�����2`].(�f:�8��@�)�z���'g�i�r�ݺ6�_6 }�O��e	�:�����1�J@[��_dk#f�� RO=��q�K�RJ���<�Һ���e<�}xx���u��	��e��f#dXȀ�ڐ��jj^�xw\z~:��T0����rUi���5�
u<H��5�j'��h�	!F��]�A�j%sԴ L�E��ߎ�V��9�&�
��mU!ߞ}��q��F��L��-}�?o �oz[H.(������?�\/¬��h�
�3 [�a��\|H]:)���"�x�L�����R�q�P_i5l&�!f���mx������o9��z��@m]�����\Wl��<����?��{+��.j����o��#��3��"j�ٹu�7i�W`���1r<H����o�خ�o��l���j��� ح�MH�f͔��>,U�Q��] �Vf|�>ג{�45.�U�(�,�	���Gi�]��Μ������^�=��q���8���ul����.Vqn��gR������a6~8�M�B
����TҾg>�a��x5R���o|���v�t��[�2.�(ߘM̖T����5�SB�&��ZS@�Z�����u/5pM�h�)Ќ6@Y<W�3���,G.�Q	�A�����71 R-���3Kj}����p;�%�A�:�|9p�HwD�ƀ�������^�W���*�y��Y)/�l��bBTT�`��e#p����A�b�Q��P��ˠ�%�����R�t��T}YW�gY�5��(�O���.���K���Cy�Y}�<�;��3χܑ��0��c���q�C���I;C�����8��I�)4��	�r�W O+U��A�M��;���׸T2���!Whl�8m,���g�����:�(�#�P;4_��i�ږ�FJr��"���'���+���&_�����$)�i�Cr����Q8%����f/xa�AS����L+AXqN���B��r˿{<��˳�g�G,�����	�$���k�cgY.^:�Z�����/��C^��)L�Ðxg������ƀ�#�D���)L�=���:Ek�
k|��LP"�̑��_�*���,�R���u9�]3�`���Hgw���l��
:���7�����$���>�$�J.�r�.L�#��Ћ�/.�>�2sʃ���ݖhH_�xʛ���������B�3Z� �OIB��}�u�*/�βs�%�`&�ZW�#�,�igPj��> aD��\D����' ��>�������X��	��"l���gȊ��-V�f�ș^�����n��'ho&? G�:,���z��h?���!�u?/sGˌ1[�}e�땏�T��!�^�'iI��3���������g
#��P*z�㿖C<�C.v���w�:3�#��)��r�c}�zם�~蕈�ͿݹY�͋\@��\7E�y%�-<��&�u|U6�_qI�?��=�^̜6gCu�0���w+iΈ����ǯ3�������<�H2��Fǵ�A�?Ƴ!��4� +n@NI�Z���ɋea��S���xb����ل.�ˌ�t�� �2��~�{�;-b��7�x���J��p #��j�7� ���uA��U4l%u�`����	jN\���#ܾv,'��{��i���Ƚ}���%!��o`ynUy�=_��{��c�4�X��,L���A�v&ٕo�!.bu��bB�~��Ë��� ���r4/���.ka�P��K�F|ںղ�FMTy���Zq̰�S�M)��1�3���`��,�ƺ�z��p������8I
��":Y:��/z�1a]њ���82�͟!�G��^*��%�M��L)Al����b-�!�G5ֽ�$��1覆�ܚD//�0�kG��Zᔰ�?E|�ޕ^�-$WN�W�_f�s#B����>��b7,�e������K�s�}���
�}3����U��E��C>e��5�n��qt��Y-�@�m�<���7\4�G(��	�{c�� &�sYQp�ޞ��A�5O��� |�?�i>y�K33�(���w�/-�NGB�p�/\F҇�����C�9��w>�;��i���&�m�=�#q�#l�x�$�� 3�Km�\�,{�=	���K%��>D;��
:%tf�WO����w��On��K����'�q�u����felR�o�����a0�����@�sm.fB���U�a6�Q��4�Z�~��*��jy��Xx.r�M&H�ڗ��&'J��YGɦ����=��B弧�W&��������G;}�v�W���K/I�����>d_߭�'�?�/v���a+)���[U�|J~�����ԛ�z!C�o0�c`Mt����i��=ee�(���:SR��v��N�	<5n���#����H�I���O�C�Ūƌ��A�J8$(BX^½�q-�_�˾�f^�Ĵ&��V,҆�A��������)vYM�M{�+�4W��C��D)�P�oӖy���N���cঁ��ܶ��%ATl@Շ��l��STޕ�L�Gل�y���W�s$',�^C�KPJ;_�R_K�L���O %>��Krv�;4Bx���E5���9�I� �&�~DM����b�Jװ����U�P¼%CM���,E��p��Zj�:?�_�q@��"�7__�����#'����k��=�I���]���`ăzb�v,U׉#��F��N!vb�'/L�������	�4� �E�^3�M�a3~?7������H�I�F�HR�;4=���RJ�e�x��G?U��Re;W'T%�eܗ�WZev�W:/����3-�|��\����Fo,��������=�1?Ϡp!;B���g����!D��4�Dr�x���^/ ��K��[��w��+F|�_2���8����ӻNI}	{5�|_�onO�MPQ!aO�4�z*����h���Id�g�S�K���<c�/��� lߋf`����!�?�oz����p��&��tD
�I:ѵ�8!����w(����k��̖�}��[ϔ�8�E���4��Gc��pq�p�K7�������J=��L@�x4��9K�����\�"XSU�@����^�m��BpDBaC�"��&g�d�?�I�T��A�� �6H��C.\������>8����m�f&R�,�9�s��+�n�2�C�5,l��%{�=T����V��I�;�7&���X�:���,\�+sW���.0vjRel����_]n~O���"Z4"��g���.�xv����;�)dᗈ��S.�}#9�JR�J*����tf=����������n��������c�6/D5�YV��|}����3Ա$��b<$+�%P���h�c􀝼&x�w���� �"Th���a��hZ�Y��Hh4G��)�4��"LŴT�Y*�k���$���Yٯ������"+-_J;��:]�BX�!�0�l�����1K�;�ݲz!��ۍ����t/�J�l�D�U������V�M�C)��ٵ��V뿗q�XM"�FH���d�n��jVHN����p'ϖ�����F�]å���2[5�d�<�-pو��(����OBx��HR:���Q�Ӑ3m;[�C+m��P���f�Ь�7��NƏ��8�)sf2��[7"d���F �;-:,M�+ ��F���Y�ʜ�8.����8p�ʟ����к?�p&-F�,m�=.��W&id�&$�e"�Hb�����F@�E���0��"�����P�4k#·�y���ހ �9A�	�m����d�A�`�)[H��<�E�S1�U疺����i�6��������?1_�L�ʁ����dq�ّ�o�� k��u��!jg���%��IL�h�˃8}�?:e��o���j\1*�T�A�k�T���_�D-�;z�5���MoIJ`��hE�#UN�� �QG���ϥ� 2��\}MN���G����Ϝ�/�(5	�g�
y@A��ת����"����_�>b��h-�������1eҺ,^��5B���}��L��z�@U�A�7����#N�̞2k'��7����;T@!]����	%��i�z,HL���eX���(� �h��"N�b+����^�����e�]i���&� *F�y�4�D)�k�ULl�� ���g�ۿ�2K$N�q./>���ھH�k�;���V��:3��(���|Q���~�of<��[�a�w�Yl%���>��U�wcS^�[�φ
y��m��Վkb�jv��=K�����X�`�RD��kVG_w�;�s��Sޓ ��L�����ڐp�p�	���(�}�uF}Q�%Z&d*�%��{��%���\=���J�g�%�B�u�{p;�*��f��pSY9]�q�t}r� ��d(��!��w,�O^MhQ`q� �t�r���qO=�Ӄ(!P�R�m�X�'
$����>�ZRU���J/8�g�"��`����J�M齋�z՜e�#Zw@�Q� �ݺClrZ��pjW�M�O���[�R&y���.T^>ŔU��\�?�`'�A�w�]S��,H�[/Q����7��c}m�B�UEщ*#�'�X3-�h���N��c�(#�;+�����������h�}�Ŝ<�rLM}���Q�go����0H�xZ1��� �{�Nқ\)`���ţtGq�x{T��:�[�q�?GҐ���q
A�j§�Fڂx ��ֈ�/������vB&�0vc�C����t%��Ì�z�������?��z�E���$Ҳ�\���Ϩ�t]�!Y�.s���;n/��c{�JM	��>G�4�󬟡N|t�X~_`�w���@ȃ��j�`�z��V�*��e�����d:�H9�R{_��7^��}��y1�w�S�yΐ�^��r�t`�����s����<�5��	.$K�,�
6�^�6�{&/�[��ܭmpy�+֥'����4�}��fv@K4,l��ʤ�x���ڇ0�d�� ӛl�D�`M��� ��6���6M����8z(�#�e�\���]߉��[���G�1Z&u�d��\�3��v;� Z`h���U�_>͟r�K��`Ӡ�JP�b�YD������u~�Ũ|�&���x=�ؑ@�Rڀ��Yd��;�tE�z�Hv���H�Դr�z<l�W�� ���nFQ��G�i�Q%ŝ%^\�糱� �Elm��'6"�	�}�ݱ��H��tVIc���"`�#e�
�%���Q�G5��\�.�
��J��Dx���Vj�;6�4鮮��s/\;ʜ8*ep���S�,�GA]$-<B>��Z��+��Ѿ�/|ċ��g'�+t�|jy̧.^,L'f0�Ԓ�_�9�Ϙ��c6����`I.@�2��h�p�q�Wv��v�b�y���P�^�<���[�e�k�7�D��k]�H����c�,I������������UxT���`	����O��3j�k'��vq�����u�$P�W�)Ź�� @��օ�r��_A>OUhۂ�b�<'ĉ?]�jV@���x޾�"���%V�'v�E4��熦n�}ij�|�4�׆���MoC>�J���������!4���9��	 �ӵ���K;�^�5�������1� �m���_�Mx���\&U�����}�j}`�i�o�oȅ�9ꡊ�������&�7���ݱ*oLlV�)��P��i�qcx��br��/r�X�"�:8�Q�T�2��FE0��׌�2�[��M��� "e�q��L�	�a"�\��A����	�傇�W�L�[�GM��H0qܖ��k>H#�qTWy�D�L������.%�/�
��k�<,͇��s��w� t8������m��y��vP�W$�!K���h���󤥐EZOy{������/!'�����u�G#��|�ˏ����3}o.^n�Z� ����F}�&��2�|`��*͟�}R�6��*D�����-P�Έk���G�(�sQ-x�yǯ�+��`o+b�$�����i'K�-E���S�@��E��
&[�X?kLhR��� ]��'� �'v�~�ltCo.�e=�.��C5�1�|�34�O�	*�6"�k�B�s)��P�x:�K\_�u�;ze:Z)w��J�� �� �H�ի%>m����p�EȞ�CÌ����R<�����!gE-��a�W�hm�-sY1T�;�d�!����X�b�L��|[�߂�.hϮ�[�e5ƚ�L����n޻'�O	fi%���9��U�v5���m�}0w!F�"������hL�v���G������%�[��
��_f��u�+��K[�gJ/i�+h�Zӂ&P�Y|�&~xxl���]�V�m`���W��$S~<-8��2s�j��:�Oa��,�%��2��d]Y������*/���BJ+�?	_���';��&#�A�П�Od]��z:�����0��njh�xY��r����	+NL�q���&�>�6/����I�u�y@
5/l�R��^�n�􅵦�֞H���̾fS~��X�'���{ŀ����иA~��f�!�M�g���ݠ8��ؔ"�oـ?�
b��
��G�]�jv=�&��! ����v�˙�x�fq$>�%�8��N����޸���q��4�6�n�����z/�#ꫡԑ��q�Ph�>�d��JN�MDֈ���-��� �8l���>k��l�������s<'yh~�?��uQ,�F�b�D`�}\���}���"��5tq��\�� ]/��.�~O�C
8��7����/�RIb��U�"3�I�K�
��5�NJw��Q$�l���[����a��˄����\FK���fT%��9
�X�9���;!NߵJ���&���B���1��d����"e���KwT
]����Y1���$.%�_
����wb6ҫ��j%a�Ɗ�as�+�M�?tk��~�1����{�Q��-���ӯ���]��T�{Na�6�ҀŽ�j�sf,#^��4��)D�u��3�_�Df�~�)���`���(5��6��7ڍ����M�~k�!�:^��h-�n�U�g�\m�r�<k�����!L�n���`v�s� ����b%N�6z:_�e����즸��]�F9TA�G��I{���8�ϔ�y(IPN�Eӛ�e�Y�Z��+2M2�<ꢙ�gհehC��Y t �����7�}�!�"��f�PF�zx]�G�/;\�ΌGk��Q���ЉKX���R�dE��g���!2n���P�\!�v�,�j��?G��7��"���D 9~̖�]�I�`y˵��:�?�:oN�|��Ѭ=����nE%�#�+�e���X�ƹ.3� `HȔ|���]+��O���wHR�;�x8�nC/WGp�B�ߺ��늧��� �갨:�Y����q�j%1��Ӌ��bǠ���I�0ۣ���f�d�F�*�d�Z�{"�j�$�Q&)ZA6^KI�s뵬;3�x�O���s��cM�6��r5[��x� b�\�ϴ)l��W�R{+.e���_GA�*�$��/}u�؅��;���t��	���r�&�m�_��5��g���}�����	&�5N`�Hxۂw�)(!�[�0��.\r������$�θ�j��xaF��0�S����Y���B��qGJ9�����Xc��1$�-B�Q��;�{Q�3��N."�|E<�
QDy�ENk���	���:��5�8܉�>I8��ٔ�8����ē����gf�vo��{a?-�C�sc#�fCP�$���ߠ��������$1G^>?�;<��l�
�S�):c5���"o�?1�L)�J�Jd�H*Y=��}�e�E�J��o'l�ݬ1��U�	�q�<.��T��������uF���&���B4Q4���o�(��#������.��O�zv���ہ�	�m�,��������E��G\w)���d���~��Lh����E�Ȇ��X&=�<s���������%l���(�5�\�e����|LV���M�]�M�k
�� �8Z�P�[\�R�%yY/`�� ��	�7\SҌ�V����p#�z��?u=���(/�W�Ԛ�릺kC=s�mv�_/����*rBҀ�!mJ�w�U@
�p {�(^�HV��?�*yAɺ��?1�P�!��V���u���)Td��g��B��tca��i�dP�Y��%T��n
��*��_�f7���]�Nnf�^��������]�!"ؑR����M�����,�J�aА���������b�E%��؛bh�m������8_ѽ�CA���;!Eb[uU���q���o�/��)n4�S+�f�����_G������rH�"hvw2�Ha{�{���$e6 m�[��ǳ˲.�;�,E�M��P������^,WC�)S���S��9`�+���|)6w��xte� 0��σ�Yũ�A,�����ӧ�E@ؼ�����Z�@� �|IH#*�¤�v.���$�nď�j�D�.@�M�ye��\�a$J\6Y�/��0�ӥ�������Q���Addu
�@�%�Vpd�8���/�d�gWH)N�'��SI"u�x�=�������l�i��Dr��B�s����;5��X��L.��{dl��������,��٫o�������Q�`�ܘ7��"47j�D�����J��T(֚�,���@�^��v�W����n��H��	\�W;�^�&�t)w��;/��X�2,��]�h���>��iE��"��V1��7|�����s�5�L4Qrk�����t_��,�H.�ܜK����^��R(J���/C��`�����\C*<��rR�NC��u ;�y�1ݬ�����˴����c���'C̰���ja���0�p����+�`��wsA�{�(R��ɥ0u�9^jgt��	{t��DB�[1xߴ��h/�iv��oK��G-A��R�+�Ȕ��	�2���t�M��ս��}�Ai��g�:j��&�Sq{H,��I�Z��O�1���1�U�������d�������$�,�I8�/���PWM��t��3�Ж)�E��<�)���VO�����OQ3�Jg��N��c����<����Hp4s7Y�sa�T�)�M-���C�Sp�[�s���*uP�tk��cHY1���7<�%��m1�[+�(��^j%J�ƪ��������G������`�|M&�an�WJ~�����V�2wRc_�xQ���ZW�
��:.r�Wi��ᗗ�X��-!H{a���¾�Y�1�-y �P�{s. �A�*~0<�W���ԗ
����譙G[e�Hʰ6���O����;×�Gf��Bke��u��)R;��GW^2C	�)�o�,�6���\C���'��g�l��"��]�~�7�h.����³���Zn��=�	�;������ɼ�#VPD�����q��F���75��㮛&q����������1���ٞwe�E����qs�T�*�U���w�x�}��I9{Q�TL_��S����rOa�ȵwƮ�1����
x� �C��I5�NJ\�̵eT(uT��m�k7a4�5��˗�^��u�Ѧ�} K=�� 
	�@��'�^&�"�b�~hլk�A�裱�� m3�ɷ�G���^��� �i���0���w&��ؽ�j_-�!�3Bh{���t(���������z
�\" 'ߘ�o�'7rCvA���+*�76�Y�<�$�f�:[=���]�^wP�qn�z�hs���iu����3d��+�OJ�:��-�m�]�)Rg��;3�W����VĄ��d�ɥ(!�v���a^z݈�/?�؏z�qm���$X ĺ�.��(��
�&M!ˇ�7�n�K��.�Q�O8���M{K�y#�ѐ��H��(v;��-�Șɞyu7w½�|wC��y��R� t�O�m9& D4CNQ}7����I�� ���H�]����wP�bK$�� ijĴUG�ji�4ks�J�K�uŔ�Ƣ�����?$�0�ս�
~�f�������*uMZ�=&�[1MVk�^��D=����P��S��8f`��B���Xd��25p�� m1�ߑa��.s��e����X�Ӕ=
�:�!�X�bܖ�u��/�;���2�.�-fEr;��[(�ru�Z$�6i�G9��-0�t�Fd&̔kf��1��i�Y<�yz�w�m�U��Y$h�i�ӭ�w�ɪ@�ǋX��b�����߳�<�{�����,�-�D������Kq����F�Te�enж��jN�L��^db��u>GHD��`ɯz�����ّ�*���ά"�Y����`<��j�D��d�"<<�~��-@�ʌ�c�L���q~�r B4+�c�l6��[�LN�����$�����+� �"Jg��~:�0K^3���ioT�������T�4��M������r
��(h�,��s�8��)^�_���N��s��C4��W�EɁWoİ��l.�9z��[��J\`*��kᷜ�Zn<\�ܱ�.nd���3^H����8�X���v�}�E�[A+�}���v���7����UV@EK�9[K6?�	S�@��ib��v�6Z��t(��;��fM��ڿ���.H=Un45�y�7�r�)��e����W�z��3� �(�GԵ;=j���\A�9c[+ �1�H��Z� 
���`�_�<7�c@��jO�S|��� �Mĵ�M�
��'I�-RT��c���*� |��|H#�D�v��zUCFV<���.��qW:��Qj?Ql/$�{f�	��w��B~hME�=ؙ�������lQ�Ǐ*�r\l����Ks�BR����/�NrwB��;�ی��8�c��j�E��>�R�~3ى��~t�PH��͒]�Ѡ�c�h��r���}�mR�O�U�O3�H��i[���^� PA�V���*$�YU
o��N���K%���Gu��.X��O��G���I���<�<,���±@��")��e��عR����~�a�eT-����ǚn�]�)N��!��5�!�!}�6/C������b���HK;n�������<ԮtC�+�����;K�8S̋g�ds�z�j�C�����K�$m�"�	Oo�z�8&׃dw?{29I�JR/k���jߚ�!�qB����3	tq�� 2�.��=���Mpv����:�����G��i�E/�������? �au��[E�V�i��7�����=Ș�������L�A�D@Mn��$^��y�.,��%��U�h����=�Q]����UoK��� ������ E`����d���vS^�=yr%��X'N��jn��<$��u!�����A���QeB�!� 4�>�
1�U�,)7�p:6��c����-Ě�΅E�y>E؏��jMn��ԟ�_ي#���l��kZ�Ȕ~��,�ăԒ "=�w�gfoݺ)�N3��u�����C���6���q~Wʒ� ˏ�6�_�jpT�tY���Y�?a�`o%ۗ^��Wb��٥�}[;��1Ś�rk�gأ�EUD-�(�gsQ2Tg���8���\B�|���8���)�l>���:�1��K��T���N%1��p_Y��7����A|`�����p�/�,��E���E;��Z�з<���l����&�'?AvFr��M�S|�W�LFK�\���:ش��H�	���=ƴo��K�8�O�o�%�8����&�����'�U�%�":��x>����d=M�Bh}�Qy�i}�d"�A5x��*��	� ^l#��˸�j�Pص����+�%�Сx�"3��́$���tT,-�j�%�~��h�Il`�/�ևW����V�t~�b��w4J{��8����n�
��g�%��e�k�[�3�o[�@�a�����= EL{��4�߬NB�����٧hع+G��v���߯�b?�ȿln��V�����@9~�D���,�!�~C|�,A���m��ٶ/0��l�;W(��"�HI(F�ǆ4D�
:e�zv�3�+Bڭ������Yłi該�kj�u$]TU�P�pX�}=��.�@��`n��÷Sxz������U��8e�3}�2������诎�̇�ѣd#��p�	�y\�q�YxWL���}c�NJ�@��Kc��v�/;O9>��:т"�/q��zPw۸8��:�:/�a��!�<�㩌R$�my� ��Q��I�8�l����{}�ڹ��G�������+Q e/ۊ1��W�w�
o�L�M�8N�����^���E���#�/���Q|
�[P#��,��c�����Ȏ���B�le$r��gI�e��k�r��Ċ�j����l h��ТaƼ3~2R����ܲ�q���#u�N2�sV�m�#0hEi��吏V������eiIk�Jԝ",���yp�'k�/o����7`q�̙�!#�
_�S(���Qj���2!;�G�u�C>zg�P���wR�¡C�8=��n7�@���1��1�BOPb���;�� 6���W�7z;
�y�:aFh��s�P��Ŭ�EC�#&�{p��	�B0>��(SK��ˎ	A!n@��j���ڪ��L/|�HdbQ��БV�#ZGh�2a8aΦ�T/�ڈ0�֑$ xK�b�2&!zrUҟ]�3ݳ��,�cP �Fǒ;L �
��Y;s�N�N�:��=�\�,�I;�>g�&�������ܩ{7��J)f�(*5>�F�`a����D0ҳ\z�)��r��^��)�Y|I���hr��+�"���6-Ű���ʽ-C��H�r�{�����+[I62����@����l���x����{sܭd�~%o^5s��NߩM�6��'m����w����0|-�w�����bI6���~6W�yM�:�k\<��|BV��!����I�c,��qg��|r�@X	�PH�;qFٰ�3A���Ľ��+��1�<��!I�Rb��c�a3P����H*H�[y�A6@^����-(_{��R�Q�����������CCd��uw/�sk�Nk�����YB��&�==d�-˗;�"@ęo����h0Fc%|v����d���i��
�]dI�1K9��>Gt�\+B0��~�>(���� ���l���Vû's�B3�@� I���A�)�b��)ۣ�a� �F�z�*<i�T�=wQ�ٸ�MkR��Q3-�;�d�#T�I{�8��j6�~���^�#f�b;���۰8 Ei	3Dk ޔ�k����\�B�ƥ	2뛸�7��1�����m/�RFdcgw�3�n��̪�B�:�
Z+}~��`�����s�_�`
���hU.�J��ޤ�-��
��8��4rU�Y�h12՘��*��÷�
�,HW�J-��8�����S.,G�V��p�~Q��P�_ܜi�)�l9�y����O�Z���Xk!�]b�]:b�;U\ď�1a>�J@���xv�Ԗ�R�|�t�쮫ds�s�N��dvKe~��g���I���y�9�}S>egԠoڥ��,z�s>���)gn]��� a�eK�<#� ���[���Z�����wT�Z�^�p4-L1�j���U@��� �$�=�CN���"Ѵ�$��G����0(��g�Tq��KT��T��lqsMD��(�ᜈ�c  >��*��ҨΊ8��%���	V!E��?��������x�u�Lc����'�����1)�82Ɇ���j���7h"�(���R��z��K-�-��aй5��t�D5 ��l�?�跩��k�@{�Y
V� �i���L$u�Ux2Pi���ڿR��R���7���o���6VY
(�f-��\��: &���sƧ��sY��/V0���w�##8���+�'�����P=ԝ�� F[�A��~�
���X�_]�'����t��Ұ�QS�m��-�i��`
Yٓq]��R��)ܨ((Hs2��k��Ȋ��y'�{����G�����斷WN5�8��� )����|� ӏ��R ���˩�׊��0��n�왻j�X�}C�G�G�uzS&����r���ӓƲ�ÿ���\$�V����Bo�М9* ��:�[�����t�n������R�լ_T� ���=G�q��uNb�62�E�@�K�q��B|�6��C���4�	oᩱVN�jm�ڵ W��`ݘ!�3�X��V|�P�����qa������#yX�3	P�<x���ww�߯��(�	��ݦr�m����9��,gQ��zT�!���U���Q��(�vC<W���?ot\&j�-j��q�o��)��b�F���}�pr]Hi����M��t��kSdv
�I���I�6�Ҁ;�7W�<�ET ��ߣ�y�A����U��a�i"�Nw��kix�CL��|�!M��֜��@������ɬGM"C��7B�<��|/E�n����I��m_T|��Hb�����C4�wu�)�z4g��܉�]���t`7���/F�t� Y���̢	���R���CR�Z�����j� ���������!$mm�^YF��%���Vx����D���sKpv�])�dڪ��팷�{���m���8�z;��i�J�����yhjbszV8
�G�c��'ã��!�i�6j����p�-�2+�T��5�':�{�ʧ�q�n�|s�K��%Y�N(쮮hݫ�<�Wp��B�g�I�[�W�����B�gO,�$8aϧ�t�/qXp�D�`��5N����Z���慩N�:�K�{�:'��B������9��2.�����ۥ#6�5NLp�H���.�YH44?-RX^����B�7�>H�DFǰ%/0���0!W������U�Ŭ�@+i��O*�5��U�|�	sf�%[0��3�ޭʀ���(���;BBz���?���e��}��?L/�?/��~�X�Z��x�疤�>��-�R����������<ԼuC�w�#1���o����[�`I�?_,%kd�'�,�TD��l��j|�x.��[�'���+3dz�s��n�Ƨ��;����`���yQ�)5�s,X_�@�w�G;�$[�?�ǉ)�-���9�	�!u�HƉ����(�����[�P;6�9ht]O�qI:����d��/�a����q�:|��\�n�<��9���m�G�ၷ5H�v![	}�;I��/I��h�@�տxa�R��ߘ��/E[�}�]1|f��K����_苬o���?C����˪~�4S'�.��@
D�㾅��p@tW%��e;G)C�?~�$䁹��gU���|0�����P#��Hr�GA�ۚ�{�jCcƵ�`w�8���#�L
d�K���b�&��;&�,�Kt�-�Y8�iz ��K�������ӻ��yƨl�"���R��7��*�uL@h����?�l#�u��u�x�;�I�q�����t.���N�0)�g{�h<v��9!�7���2&���m'��r�VG0��x�Hs��Z�_�N�|�n��&L �e��6A�;�
�E毝!~a�9�U`�g5�Rhr�m�]d����rW����_�@��l<oIm�7SY|r���,�P~9=�4�+tg�	��zI\mi��
�s32d~�ywS��z���e�Ғ��Qo���#̊�4lsz����j�%1ppJƐ" <`�EF~q[���Wf�5�b.��K�ʭ�?���;ါ��u�ZM]~}�Yt��gEQ|�FYl������/џ��#�5��B���5����)�Y���@d?0�Ю����"�Yo�hx��Y�\�1s��+�����AI��G}��� ��
�6��v{��-�@�zP���x�к� �b�(��<�D&����� �c�c� 1l+��w�#���u�`�&˲^��~��>���63�EݏV�~���n�|�M������Fғ�G�*��pa���nt,KkG�cPD�/�yvf݈�i�?��C\��cyI�Al>��jtDd*�nS]/?&|�j����Z�o� m�a}E~+�j��ʪz.��//J��~�;�L	������e���0^ӨD-�������K5����l��ْ�q��hsv�XQ�����n��)���>��,�$R3]��X���Ӻ`&$�/�>`�M�A!xa�.�R-
e�$�!���mN�#�L��)�I����(��yk���}֔[|�F=��F��03��r��Ǚ�L��_B�|�3�jp2ɺ >h�	�][���{�68z�ó��
�m���Q��hKOg�N��)�
�4xƷ�S�����q�t{;R�<[�2���!m7SzN��ga6p����]~>D6@2n8�x�x��*u�9*/k�M�˲n��\@��~0mN_�o�!��fY�=s�['�ӘX��|����E����c�B�o�ф=֛{*�1kU�?��*���#���.5.�������1֓�t,���P�v.^�a����Љ8K/j��dɰ��M��4e�|�Q�����C�5��ʦ��}��?���ID�3�4mQ,7�۱=�n'�Y���.��Ƙ}T��Z;ƌ�􄴎��}X�MƔsX��J�M��E�ǂ����Z@?�ﰍVȰ�o��4biav^���P���)"rLy@�ܘw�>����X�����9&E*������]����4D�HK?ƞ�����5��ML��G&%��9��(����F�<����Q���gO�yW%e
Q���je�?q�Ӧ���z�t�Q��=�-�5K�wI��t�H�R�qlԕ|�Ǒ��b-�y�hx�7��]����M�E���;�b~T��$%<_���ӫAi~ʀ�`\Nfp��������3����}|q�aT^$��2��i�]�vG#�|mE?>.ȸ��H�y9E��d
�lVzfG�^�@�܊?�5��l٥̅�������uxO����~�_ʫ�'�o���%񦛫�����J+�o/�\��9��`L������Gx��1��#Rv��w��t��5�5Չ��ڈ�-/��P�ac@|���L�XDQT�
�2{���2e�k�N�׼݆=�A-�X�v\J��j:���~��/`����n�8���lQ��Ꮑ~�@h��ző`�y�	@K�G��F�n-��OtPz�k~�#��`VtN�u����[L���?H�-gk��Q��
WC��]Jf^�X�9��ڬ�oU=Z�|�D1�)T��Q�{����+�#�� d�2zE�/�bŬ�xS ��Z"��n����)#��'5IFJ�?��{
�\��,~�<��'���[5��� �
�M�XxB�)
��0'dC��9/��u�����m�����r��t��-8R�t�]��a;�]ϥL=<kF>/q�4r��s�!tl{?�S0׋2���\�ar+$��!��q���1B����&��_	;�����(g��<�du����a��_B��
������������Di�{���f/��'��_a=��yI�r71��� ��t���#�TN̓�?�Q��f���|�1��I�2�/Q7[�H�9Mj�&}4�$Tg�#¼�sC���Q�B�9�s��H��$�����-7(CI��[4�V�a�+���<H=vOm}���Qˑ��k�|!X8���[���W���Ư�������W��Y��Nr�p<
k�s �(뙼���y���<���,[W��4��1@��='v�p2/������S�v�G"w�
x�w1��EuB��P����9�E�!��{�(Ԋ��g)a(Ǟ�-��T��Źl�=࿉�?�_	�4ު:}k֔��
�F�h�c��MR�m,�����H����d����6�]�:�^�m^����t�=T�ǌ/�ЏR���o�}h\X"��c�Y;��ѫ�ޙ@F`����A=�� �`�z":�s� ~O��v�}��q7��q��2>v���K�[Opn�EU���2�g
wb♑�c��y��o;9u9Ʀ�d����)�ozz��u��1�qtAȝ����J���Ɓ�^��, ���/yDc"w�l��3\2p��ɳW��h�yYU�>�|�ìd8�ƃ[�4�"̀��\C����q��&��5J������w�o��|w��5݄��w�#�N>�;TQ(�+ɳ�O@J	�,�s�h)'�P[�L��X�#��~ΈJ�%8� ���Rt��T��~e�*g�Sy�X:�6�|��}�tۣ�"E�Oe?;�ˍ0�4��8�JH0ꃚ���Xs����#�C~� �ѿ��)��W9�EQA�]M���\��>s��pg��BLJ�[���m��c�H��=٠�um�O�=�����[�|�b��S�׮D@��������b������U3�6���q�x $)*�1���eu^@�$x�e���l�XN|�< `8��Ydc�~b8M�.(�u����؃E���d��fje9
^�bH2L�/vۿ�8�=u�֌��\z��TҢc8VuTQE�22��*�����9�����l%�p�[��XP#��ݕ�U�a������"V&<	l)UO�� �<z�CCU[tU�Q)��+�:qi;��Sֶ�:2�c8}�Bj���q�O0)��z�!%n�K����ױ�E��R���6����N4�wE?�-W�z�ħ�*L���[̔�����=�y[륅~ri�A�N+d�0$t�Fa����ƥM85���[2bqcw�f�xֳ���N�"��W�����$&������m;�[��L��!�ՏJ/��Z3k�Z���m�xT����D���*�����$ƶ�w�	4�1�q�����)`Պ:�[�sk��(�T�©H��AҢy�-@�~hu���I<(Z�j�57l[��R���}�5�P�%tY�	2��E�וi�9��gl��M4@��q��r#2d�O�F7q�t�>*Յ��ƌ���R6�0�I��> *�,o�2vϗ�:,1���5"swiɃ|�o�62��dV�aJR�=7��2���Llj>�E�%�TM\&����z�x���vU�\�n�'"M	%�Z_-�t��i��ǰ��Υnn����Rta�d7�����r(��*�f�E;2q��({��eDnN/�u��K]<V8i��M쭹ޤx�����3�'"�	4|��o����,�ۣ:��O8��,7�}����!��ر��[�WQנ2��6%щl;К7r2�0	��b�Q��EBt���U��(�c�oOS,@^�k� ���
��^�+�Fvt����L^'�`5�?�N�a8~�쨠����9��`����&�-�X�iY��3i-��;c he��8`�Wh�����k}�}���M��v��̶�A�Ry>2�iڽ����_����LAZ4yj��.QM��Bt�u�o���>���m�<9c�����ޡɤ)4"y�C�)M��L�+�8,Y���
��d�kA������N�gNo;�Q�gc���W�\��bo�c�� /6搌����>��������ze�L��"���,?��������qF��wV8�F��A�S��	�(ͼܟ�����fb7W�`�� �5	�6��I�<a4lC(>ּ۱��;���!��>�$�Yg�U�'�)�f=�K�C�U�FSi��ћR�]6'��ŝ�âi����\�	�L�%��²7����y���"���!�x�������{���&	Q�����c�W�ǥM��:m;;�q��{(/������-��hyGEz���T���*��
s���Jb�G����s �ד�6}���Q����W�*`%���ub�#��Sj
��� :r���������+ 1`���0f�jב;ឣX��a*='ao@�x����� �1ȣ���ޛ5�w�Ӗ?��$����� �FI`��>�z1N��r�����-��A8�3pK�� �+�	@�|XN���SV�)߄����Ƞ��S��jt\Ʌ��Z��ze�[TcVb0�h�J����/AG����;
yb�IE��/����'%���_hݴ��I�c�A��˿��s��[��슴(Gn�%Tߘ��ds7��=ȫ���\\w��G�}7��|���F���~���@koQ�J���B ��w`����A��С�u��]I����	�5�{���j�y����}D��^IjB,���͊O~7v��nb;�E_�J4ˬu���� ���a���Y��wdcE�a��+��o��w;CRò-B��Qe����݃��D��ՑLaw}�Iס�M��+��d�X�^���2[�cQ����uqՑb�|�&rb#1�c��u���;�@���p���4�!i�Fz5��?A�YD��y�q-����p�"Ot�	�t�������^���2߱�|G���͔E��GF<%
���2�MEyNrrD�ۨ:��fSۈ�7W�^7�iK�]��L�Q�S��M�?~��qX�X���Ƞe/"A��cΟ�P� Ȧ�|��^߹����#����� �9K�.�G�O��m]��� ���鹌n�G?)J(��CU��~Z���V�Ђ�=��+����+W�)
���؆�D��F�ܥ��mN@9��%�>�����;��PB�2�F��X1w�x�b���-��0��Yn�).
K��� ����z�F+ךK���}[ZvF�&בn)6�<�����t�6��vnM�%N7t�k��G��QO9Ӂ6z�/�W~����L�{"jў�����!�M_|���g��~6"-w�p�X�����xy����ʳ�2&�r!GGq
��myb�Q�b�8k�&&��+&�ͫ�j�[]4(r0F�Xz�8���G�
�zb�@�ضL�����e����ꬖAn������w�ϗ���]��+��]'Ū@<|I+��t����+@�[~�GW�~�G�����\��-����͚<U��~wH�;G��*�[�:Z�!V����T7#�3ߞ���a��W ���Y�@���8v1���f%<���X��0㇝��ά��x�����r�LsԖ�D,P�EZ�_;AM����F���G��"4�.�R�C��}j�z�ԉvI,�~�.@|a˩ FY�!��{w�n��Q/�M���.+�<�멦%ֱ�5-`�_��cL�L�Z�vh���҃b?��dK��,��	��A�?����T�zW��5*�[�*� ��M
���FJ�U��mU���^
p��n�f��O�K')��7�
��׼l�i��� 5�4ݧH�7Y�	\��'H��7�z�Lb����LI<;N����1���鲲d���y�ꨯ���e`����qc����W�;��{m�ۀ�-Wm����g;C>�_�W^��3t�w�Π2�G$@x��l����Z@��v���j�5A�'��(��,��ȇW�����p�h����w�;�5Ә*
� �_I#--8��8�i�S�
��&��.rP�W*�v��-�X�>g������m�B��
�G�9�������*�$V��_U���-����Lq���gh���0�FRݐhN�~elh*��C���݉�L��0��%��m�� ���/��CR:����]�2�i�����$.i˝�#��O� R�B�R:��4��
�&��]��I���chV$͎ZT����S���g���]ܥwL�}�R�kn��n����n�š�{*��*+@���⛶WEs�d�H��,o=���c���R�N���W����fm3#0|�Ά�e�
k���'+����/ރ,*۸D��߶,�!�y��������-�YRBAU�Ɩ^1|	p�a��V=زg���u����j5�����?���Љ�Hv�i�c��1���we��㨋����U۠ni�ڃ��'TA�Ht��6X�j|.�]�o����4�*�!_� �������dۍ
���ɧ�]دc�x���?^;"�����QS�˘ɳ����v�w�u/m�{K����x֯�u�"���0���t��`�w�d�ܡ�[ w��y	�D��y�p�������E���rTp��1iP�Gk}ƨ���˘�XiDLѹ^p�Q3�6A�+�F�J��0�^���\v�p0,��>��$���/�Efhg^FLy�*n����h<'�*,��v��8�-^�׃~G�2*��	���H_`�5�Z}~H����&JB�q��;�g�TL��{��H�?0_�<�\vc�������izB�S'-ΥusI����M��
2�K��gN��BDk���W���?���R**�IB��E���2���73U�>�>�Zu�[��
��W ^���\D��P����u�t��ㅲ�k��=����a���a3��v��E;�Ϸ�X�<n��}�����!*?)�P���L󭺺a+�9�Z��9�P���'㮃�i�������|���t����=�3�7���a���&��~�4:�k��;�s��6>8�&kQR��~*��@�C~%��'P��,)�p�r���/M�����z|��!R�̉{���R��*9��%�w2��J����W?���U��?"넣s�F#���DJ�SU�{~��4� ;=ْ̱�	���q�@)���mEnc���_�^}w(�k��U-�R��\�H� v�n�!1�Ǘ�*�Kw�k57[?(l�\��<��� m翈,����}ޣ����g`��_��W��f<�E!��.��d���?����;2�U�)��DKh�,���voN�1�	��+aQ��4�{��z�{�Y�f����Z��θ��j��IP�ߗM���ު<W1��v����ۛ�ox�e�$~�~�';O�X�P�
�id�+��.zRY�9��J^�6s�/�.�g� �S��v�s�y8�0"{���]�A}CZ]��T=Ь��b8f���?��WCp����$�zb�T�5�>I��L9�6@��<�q�P��hy5�3o�c���P���qw���x/ÓH�����X�M�RH
m�AJ��ؕ�����p<�eF�9��a1�0����;xZ��W ��ȿ�*��m�h�}��+m�����i��Qg����Q#��9d��X��4�6�"�d�jܫ�I��}'r�E�ʹ���tcA��X��H��ԶL���f�Ew0��{{���)���<>�i�XNg��ۤ���UN=���u�.��ML��6ˊ[�\9�E֥񔹆�2����H���I�_M�`�<�I5u�=x9%n�BJ��4��b�]ϼ��0|�["���(�yU�1�8|7*�̳�������FU�nP��'�h��ٻ����Y�^�3�ecc�2gd�����K@(p ,�T��j�e)J�*N]�&�Y�x*�6��\�s3Y1��=�=ȗk��k&�P����ua�E��&���U�Nw芽�fsG� (H	�%�Z���K.���̆��wi8.���h%��!8ҩµڰ�5����~�l�c�9��e��/����@E�U"g�Q�,Q~��˭_��o�pP4�lۆ*\
��%>ٞʣ;���]���A��xٕ �
�@b�ٮ ���9P¤K�k1�q��,���0<z��$6���5��aQZ#�+�УZC^�b�\��q��_���H�[�T���h�;���1sI��]���xb��x�G����.���i]"u�/j���,D���eNR<D��w���k=-�|�0hcc�ʝP:*��r�[ǂ��𳳾X�i�,!��&F�=Qb�Iq�����C�`����<3�p2�`&� ���2Sh���Vx_�����|���~X�7����=���e�5���I�p-�
�`a�LA��m��?Ɋ=��������|[�YE�vo�vEDnL�'EZҡ�/�(f��V~�C�~�����;�ǿ".�ν��:#+7m_t�^��;��2H��݉� ��IL���S�k�䇃�:y�H��X=���:L��Ti��6�� ��H��^�����2I������j�0ْ�B�v����oJ��<�L:-�g�YY��]w�Ƕ���z`��`ʌ��c���"g�s�9���N
�D���ȫ��(���;�oH$�(��qw]lr���0�yB��>��JH(~U��	I� `��d���簱�I9��1CM�����q�P�vEO���8�r��_Q�:9���D�)|Yf|��w�����,�G�m�5ڮ� �k�,>��3G�qs���ܵMQu:pڲ�4\B�=�ɼF�fӽ������چ���׭c��,����L8�ė��H�[��<��\k|D�gQ��ҫ�GI��*��6$��?���}��RR���K�BpYzO�wrQ�����5��㿒�h�4���|?tv� sĴ�a�+}�:rA��������<#�wk�:�ņa�=��4�k`M?N�i�~��_wx�/-C��=�n+aD*b$��U��]f6��I´�Y�>n�-�s� ���v00��w*q�n���55w��<�,PqM���/�B��\�z{M��kN�I緰ż���A�e6�֩���(+��T,]j��>H$Wj(}�� ��;5�d��U\ҟ&J��^Y9�rY�i0h[��yW�$� !M��Ͳ�Y��x������@��muD�(b���:h�1�Ӻ_8\�*_��("Z����3?���X3;�Wq����R��03�������H7Ģ*M�P��K������\�&�5zA�=h��m�2���)�b.�T�ܖнE�r� |gī�_(>�%h$�;�G�O<�:B�x28��s�է(��qE������!r��|p����:{�VZ3�WӨ��R����t�)ܩ}�7`'&���h\N�2!�M��\������]bA-��\S�5Vzլ#YY`Z�t�Xǜ iuK|U�尀jS���� �e@zj��8Wu���[�"��QK�o��9��#�&#��XW��eF�"J��t�&T``���\h�ZUhĢ����.��~�3�����m�
3�E����0� ��j��Y��~�&ŗ۾�Q�G�v�:Χ��7z���([�Uݬj���|B�[(t��XPb��t�����D�Q�[�����?\����x�&�|�Q�pH5�֚¡���,H���8G_zbo���h2T�6cJ��\ ��H]�z�N4��r�>�ZCXѹϠ��Z5�P?y9z�ʬ�o��Ջ���F��
�c�+���3'�o�"��d����~wd�8z����\Qs��_/˗@�ZA�VvJ���鍁���)���&��AY$`��F�-f���D���ɪ�+Y�L��f�SU:��W �\�(�!ږ�^`�ݹL&�Vᓧc��9^�0!�t�L����mɥ�5Ljr���KUrI�o���׌�������ϻ���^��j���y��Yt��k3�S�i"��̥�y�Sg��S�H��B��A@�*���R�����A���' �W�MA��70|�f'���J�\U����M��!jr:~w��%D"ħ���-fl�7=��غ�8�ߠ짮q�K��
>��k��Z1���0�D7��	M����4>;xQQ��嚟��L��_E�\29z�𪬑#��[1i2N���T�i��h��A�����o��,K��d`�;�`���P��]=�����Ү�-��{�%��di��;ޛ���x����X4H��5xp��y�sY���:�@[e���J�g.~?�=�u *��[f���@�س��Y���
��1k�U�;��|�����a]'���`!��M��������T�t���r��0;@p[���"���!뀄s�4����Ӌ)��}O3T&)m{�[ʝ�3i3|CA�%>�2Mv�(XA��UH��}ԫ�R��d�ы��αҿ)��;Q ݧ9��k�2�~��V�]M`�)��E��A�p�".�ɝ䭁���?��d#TC�&�����X��Rf����QVw��}�����X���d�p�ܚ���-l��O�.Ֆ���#\��?�2���7�%�jmN͚��g����3~�(��k���S��P��� �M�t�ͪ)ԛ����JIU��״p.�0��q&��}���B��d����*C���ƃ$���ȣ�ZO>HE�V���VxH���������<KUi�����UA1�;c���V|-� ��V�{�"�������j�X$b�0}	��;�.(����4����F��~��b�lJ�E������Π�j�Xs�����;��P�/�e	wr�t��a��I�,� ����X"]x�@��
C���n���d+�P�?��`Z����S�4����?Ĳ��P��|oɒ��*��-XM���8�0j��@GVC!����|�+z�k������q$� �\8���ZQ�3����E���RR�;��0; �rאx��)�G�zM��p\MpAxI�R+5mS�L��qA��F-j��4�|�QP_�*�+�L�96뮟a���'g?��t�x2�W⃾�R��"��Ei�W�G8��������[MV��3�D$�k��X�%%��q�����/�S�-ܑ�E��|Tc_&��8�f��ݥ��}�hb卵���1ힶO9�:5J�-����
p�(om�U��R�S�-Bm��b��C��W�M�dPR�vK�wQ��W*s큃跟��!��!�@�;ٖ��bG��*�����&��)k�n,icIϩ�t�B��Eq�w�$�?V��(x�;;&�>!�{@A"��Ń�2|՗M�j{��up���r�YO���\�P�;F���p�����`��c2�z�H*�#>�3���ꈱ�w��(1���oz��l�s��Q��-���T~���ʪ�li�oq�����dD� ���92�}��j�5������{+�<�'NŐ
�� �,=���^�пyΪ˫��N��.�7*#�t3~_����C|�	n*ն���J�f����Q�=��<nx����-1K��aFe����z�k?%�A�/l6��+���\��~��j��KeZ���rWcK-�y�2|n#+����],p"T���U@g_n�z�;At��ʶ���Hv��M�WuT�TH&�1auƩe�<��UE:�KN���eRٽ �߈���}�
q
��Ӯ?���Q�b0���S"k��-M˯@L"��dt{F�>wec�,�(��Κ�v>�}��hQ?�JԁV�n,�\�c6�#j�}�Atn����)�A1D��̄M��9���U�s����3Dʠ�'���yqEr�#��7�ZӐ�ض��l�IA�����0AW"��\�=mԧS���b��,I������U�c�i108N�f��!�q�Г�B��{�8�b�e+d#*|м£���8ܿ����H��hT-� {r��J>�rl̚���%g#�(U�P����N���=�2��A/�yT��Lďi��j�u��Oȑ�Ф������MDJ���6E��
��;n=P�
\�4Y!f�ќ��<w��5��b�	ѠD<�B?���,Y*�����������؀��,���|�ϧ�5�0���\K%r�i�9�����FM1�~c��A���&����P���}��rWT�+ɵ��~��ߚ����p�a��`��u�
�&O��>;�G�ۻ��5|(������Z�l����#�Z)�8��8��Χ�Y�����ѯ���ʨ>�$ɼR�a��4{'�2-�x=h�"��n�:)/?P܂}*^��B�-�F+V1>�w�R�%���ֱ��7|�=7��澇	ݏ�,�/ өґ�ԃgQ�>�M7�ijd�A�l�@���l։l��46��J�9~�	5�YM�+~���AB������4��a��҂�v97i�Ͱ{��[	�ω����"�=�J����}_����~#�X�#+'�w9��ݾ!��D�MZ���wӵ��h4��V%�����[e�h��s�����v_�~��,M<4�|�K����XWr���`}�y��H�a��'mw"8�;�|�l��6�`&[ijADZ���I_�#F������u�`�	="`Zr|s��INs��dw�n��]l��B6]��3Vw��I|�`�}7\J�k���q��^;�.�؆GOD�~X/p��@�Qg��'��TK�4�댊�#!d��&�X������q�׼�H�L�j����/_[0���Kv�-���ܡN- �t)�N w��7���,[2�7��qW	���Y/�ΣА�峡QJ�'�}67I�~*S��;��H��z9�t?c�r�F�g�J�\�&v�-�����je�.M��Z\
���~���/S�EQ*Y�1r������I?��jW�KGb��I`�2d�d���]T����������X�����3|��_��B=��]&9���s���G���P� ~M�=*m�%�f�UC��T���*<i8�c�#Rhk���E69�����h@v���!�o�3���E��V�����7Q�#��xk9���f���
�!L�0yE��b/�dɷ��<AUs+w�xh��C��$����]����̋��|)�
���=�+qC��N�W	2�����v��p��-#f���Π4�T܀�ܙ���9�M;Z��V�"�-v�我��SL�����L�5&6P'ĝQ�P��̺�6�Wmu����ZjwV�F��ʡyݵ�����	n7|e���8�5f̡�Y��mc�n;��a�kFuA�����bp�R���� UL����+SNA2n����gi��3s�����_w��o�I�-�5���F�W*3h�����ȅ��U֐���8���( 0��@97t�av���(�e�y{���3c�֡F@��	��w���Xޛ"�Ď�<�z���xi��z\� ��'���\݌�4������<�'ǾU��O���;�'�]��AuF�"�-+,�ʒ�<�aׁ�v1�}*�,�X�cc�l}X��0Zk��i,�����WF`p���C��Z���%7�1L��=`/m�P��zH��J9ݘ��ޛ</3�n�.A3���� ��OA�o�:�TR�d�:�1W?aҾ{Ee�8����x�A�S�f[sxt``�~�~���5q,LW�h!�bn~s'����3�*4y��X�ʖ�^j]:�o�k�v�5��љ ��]�Gʉ�S"$�h��ֲ�o[�s���oX��:HvΠoTE���$zF��ل�+�C����=]�OD���S3���n�}�m� Av���x�;�%$J��T�0�٣�JV���\�*l�Z�|�T��A|́u���5�,|����L�]�{���eR	�&f��h�1�%���#�~��w%3���	�OG�w��K�\R+c�]V��~�-�I�s}��K�/O6�1�!�8�r��9�8Uw�˧c��TY\�����HxG��
z�}�������~̤�z�~\���~E�����h0v���gzKǘJZ^���~��H-��K�����Kx���n�����C�r�)S�ߖ��X<�;��?8�c��x4�8��;�����l�@D�����,a���x���KN�;v�T��@�#|4o����
��M�y�SG	��*P0�7�24����{*}<�3��x�5���r0������1�{l%�p)g�ec����x�Q�������BR[묋�ev���>=��cBP{C�Ud��9YTZ�lb#�IZ�捀m��G���EIռà�v4Y����L2}F%MI��$/זF3�G������w�v���BBxl�Y�+�S���b��g®D��P�_R+S�9z@�ڵd���cj�`y���B��Z
����M�)��M�Ep����ql�\�}k�@�B�'���[1w��vA�Y �|�XƧSE�3�����ܓo��eß�q���Iq�T���r��/����q�,�ɾ�G��Fd���o2��$�O*���\:ט�DZnۡ���wCx�6��8�����=*�%C�,�Lb�i)b9����;�0�Ӊq�G��K`��� 2��s�t��h�4qb����Y�2F�td��y+A�J��i�w���L*Ⱥ�j�Z�vu�wsğ��oi@=��'��CF��6�#���@/2ʃ��f�Y̐'a�^��T�&�_yfE�����&i袑|)Q�����'�)97fz�*B逧�w�l!/Cė�@��6�i�$��b!9EL�z��/V2	t����n��������ca!�0��)AV�^�&n2U�"�pr'����\t?V�����i��:�`/UE����3h-c2�e�0��p�#'!kT.]��\~�� ׬��\��0���k�RKx��?���)�ѷ���O8�zy��3'vB�H�k��I���fԁx��ބ��FZ��k�1	#�!���͈&��Z�	��K%B�-(��Q�B�_�.��̧� \����T7Ѿ؉.�6D�%��-����d����*�v �:�H���_o�I/�4RJ��I���lqBt ��@F�D́5���@%��[SbX_�,~l{�9�c���}�i��be	�r�O�ښ��-QRZ��<|�\��̀,��@����C��I���o��m��h �sπb�d�Wt$4T9͚LԧW�{��F����Dc��=x3N���U������qy���(�����:q��4�=� B��J@v:��g�v*�*%i53}?�����dUtp|J�v�H�����X�O�X{�M�c�����VTrj�,lg)B�+J�ע��t��[7�&D$�e�,���q4��R�O����w��`��(g��;�}[��/vN�G�I�J��d����������B|\רtF��]:ܷ-���,����Ar½�z-�k�sU�[t�sJ)�D���HT�%�@�h�6��Y��G�AD���&���ZG=(O���{A���=Y�Ŋ"x�c�n�ܲ������A�r���B�W(U��cx^f��v1`��ղ��x�r��yS���v׼�[�FE���nUPJo���Ŵ�w�P����%�f�rh�n�̝}ɶ��1؊�C�Y-��x����)|7���	-�j%P�O�۔�A�mz�+R�7#DT���DM����zʈM�H�����%aN=��w���E�ǴJ���'���w�\��X�X��Z1��4"c.�2��wy�u'@S�ϵ����+�z�x�.X R�����q;��h�ׄ%��q3ax����,��!Ḧ́j �ʶԐ�u�0W���f�{xV�{�s�Әͱ��{U�EV�&�̍��	��޲sD�]5��녗\�/&��P��ʵ�]�uf�$#EJx�b�K44� ��W��cJg�}nb���ƈ|�{�����^
Xz�c9��\��7y!��4�0�(*Y�/@�U���?tJub�u�4?�?�8����'oa������R2��3��3d�$�� ;��[c�9�LMt:� V�p]-����t��=���yo�k�Ix�lnj�6ű5l3}�T�N{�� �x�G�vH�B�+�wgࢲ'<K��x
9G',FN����/�$�c26�5i������C�&s���' 
e�R`�}j��BQsr�ٴ����)>�$�]9R��pn��X�¥S��:�V>��C���/sM�L�`'���(��7��Lv�@fH"g؟F,��5ÂOjغ̖�jO�!Y�(~0�d��~�QO�R�<�� -�]�^�6�s�I�:1�-c���3{��
� �~y&VɭïW��/�M��
�	��7ɝ7�k=��t��LČ��[�+�+���0�7/r�S�Z�ٖ
�0? 4��2尝<�B��~P��,ƃm7*�$���\S�)PQc��K"�JaO���\┇�����[j�A#Gg1�)���������1_��Rz7QTζ
�L���I��6�P׾�>���u��vs�׽��N����.V��j,w%w"�f�d��%�����?�o
wRX�̌)O��O=ñŴ���Z�]T�-�����9�QN�l���kJX6#l%6�g�0�����,�顥@P�~��Gck�� @�[-�]�%j�l_k�b#�)]�+�Kd�U�*~C�P���&�����<}���_
R��[�J5���B+f��@4�����Y���h�g�.�1HT�({ �*<�Es�]�<�����A
?%�me%p�(Y1X�X)tz��T�ON�G�o瘿٬,���Q�Q�n���䩐�~��
mRj�M�W�@͟w&ܧ����	5xO^%����m;A����2��Y�ޭ�]�xǇv���4�n���4z��F���g�I�N�y�i��[i��8�'�I�	�g2�4��'�-W���'^-K�s�W �{� ���qa���4�ջ��#g.�x��S.!@�s �M��;e���.8�4r�Ԅ��+�+#�2G|��k�p����x���T�Er��V0�NG�P*�Dj%�����o�p9u��i�6�N��F�{a����dϊ�Â��~h}\iO�?*Y�&O#�â%�L	<��D�%kC�}ށ6���ʶE��+�u�X�
��tN;Qa��l[-�|�_�"}�w��SH٣���T��FC؅pt��j��tKz�]"e.�+�}��"pm]|��䋺ڷ::��D\+�	��4�AE_��Z�ub,oݕ�4�;{���I<B��SY��t���(�"��奂Ó7T��9{ �;2w�\��O�"
�Z��@k<��mK=h9�Ͼ	�AnA���c���P�~Z"eNz����a?�¨�����5w
�!�@����q���o*?^Ѥ�:�"K�<&"�p.�R\A�QĔZ�T��P�3���u�U��`�N5w峎�sv��97B%���o�+�|^=�#xX��/��9��I�B[**��D�R��P�R��D�S�g�����6Î�J\lf�e�}Pp'^u�۱�:-	����[W{&m%^OۯK�u��BX/WPu���И?m��=9W:Gk�ρ��|:��f�d��G}��x	�>�Pi1�O����%��<�n~<�����i�������$�6�O{�~�P	��8�T 4���tP��f�T!�jqW�A�e"-�GC�e��r�*99��ʝ�����hm+v�X( �%���r��v�|'�>d��.�p�+�&�6��hA��E�ҙ2�}�[����k(�,�{[t����2:Zs� �?�����b��Yd<�\ǰrSC��<��;��i����OĽ�(@
�������ﴢ��I0'�&�ǳ!���W�+�
Ϻ��z�(tM1Y�9\�?S�r�ʨt��U0c��>���?����Ӳin�s���So�X��x�ɶ[�S�v�]���>�ǩb_�}��x�IFUl�,р#�Z�,4I�ᅤ��\�5�"���Y��FB�e�YX��nK���L%�6sC�%h�3�3K'��+i�p�y
��UB�7�_�Yf��<�r߬��:O����I���r���5y���J��	�k���%� �5C�~{�~���r��* ��d<��ZH ����w�C��֒�x���hy�vh"�	�{�i�R}��G@JTvl��t���6���~�g"���D��B?��-%�̲�r���ki���g2$�J���Sek�,�*	r1J�O[��s�+�ʩHC�8���)��+�OO����nI��l,
�PB&���8���t���$���I�W�A0��Jo@�5����e��/���)��:�Ir��jET���T]�:��E�MJ{|��E�[	�F �차 :aq�1�j ��
*�\�[hz�D���M�1�����ЌWߑl���9*h�i��������w�g�'ƇhI2N
4��N�.� �:RJ��I���S��Ȏ��]������ĝu7�q_��˜[s3:h�%�2mK+�͞���s]���N���P�zD�����:�R��ǳx��%(~ӭ%������#w�=A���Mt�t:����[O���G�W��c�~�	�敏�b�QG#��^ �������E�KM�غy�VO]Ԯ��u%���&��q�x��i��tB�q�����ksGu]{�.h�R���Q�UƘ1���6(�Bs�	xd����.X�wa�𑭹��(�A5�nn��U1�9DVG �֫���Q�^������l?�'d��'g��"��>*�4��*xa���_� �Mt�=׭���E�k蜧��aI����K7��½����U�9�6�&�kg�'*�!rj�C�Y�z#X�G!'JğJee����VpGm[O���/.Ɣd�j�F3u�,<�H�U��U�֝_ӳ�j�"e��F���9N<TVY�r)��Z2N��Wj�n��H�*�5�����D\���r:���RȰ7C$��8�*���!ƥ䶢gb8�������nG���e/K��Er��Y��l�O �"qy݃iVj$�<�nA(�@r�""��/���17�B1y�����$�=�4>/��Aj�&N�?���I38�.��n��	d��-�a��a��ͥ����M�E��=&/����j���3��2�k�So��� Ɣ$�xɆf��|t��M�p��7ۓ[�����,�H�3�X���}~ԁ8����xG�G�q�Uq����*�c|^"��h{>.{�?���PG?�᫨=�8���Q�5���0��y&seKLZ��q�ݚG�R���?�W�@���q4�4I,�1���c�e[ E��A���������7�!�O��j%�MR΋���S�`��*�ϼX�r��y`{�C�|�?Y�� `@�o��6�E�`~����*I�{�� �[���s/�Hv�8�'d����hT��P��k�(g��O��C��*2�>�WZ윀� | %M��$8�,�0�PKq=�,@Aԛ�r�3�����t�Mk�����$����HqRss:w��\7�h�Y����)��U�$��Yx�9�vj��1��rY5.�������&}t ��Aø��.1#��d�c�jI��L>��b��A�����k]��D��u-G��lD�/_�*Tj���9�e/L��KJm��.�N��(������h�~�_xRTqA&lq�2��?'��^:�C!�.� p'�\��~�	�1��w���>���	�pԠ�WL)�� _ТtV�	�I����WP�Q�x���:�쬣c9�g�'����ǠWc�oGn�t5l͎(�V ሧ� �$7Y���l��&@ ��oV���7^@!R��)�a�|�a�C&��kD�do�������0��Z	�ް1s�g��=��}#耏�_�o�֤ZB��6Y�ZM��`;��<2��u(��:��d������#�������O���&b����*��B'���:��sƼ
_-�
g;tߓ4����3���d�N� ��︥��7���	�*����Ԅ�Q�8�I_��n(�DI�?˜�AV2�N�E�<�`����<�z���V����Q{�zU@\�Fk���w��b1�����Q���3�M��'w�C���m��;��#
���U_���K�wTLu��J ������߯q.9U"��9���m����/�&�.7��t��=�=���z�ߟ_PSۮ����Jjr�׃'�IΥVfjt�0C�Kox��5��U�Y_50ɲ��:�\-n*;B�_#�rj6 �
R��|�$��S���5�,@2 ��*�G�S���g�#Q���?y�)�Fcб��KUn���Ahxz/'> ��Z�	��@~"�t��𧍫K6%�M�j�Ef����*�5�O����S�:M~�u�j�n֤C5��ǂsфt3��E� ��ː1nĔ�ɑa+��|uvo����\�L���$f'�*<�R��{�4���YP��`L+ nS8$��@�"h�� F.㮝MV�eI@u�.���I�0�E#IGe�0-0b,�!F��N�%�w��M�䫨����s�.�Q�o��.��=ε+��C�/���0����Г�L�mp��N����B��G?�nP�_ӭg�ղ!�\��e��+���8���trr�P��`4��٭k�E�EU@w��P,n��m�R�����G'��z���Ú\q��ɲ�-(L�m���̳� �{�mY��C�O�My�^1���sYz�-�䠦{��c�5y�%��Q���y��A	 ��Sݗ��&����ڨ�S�@��u�+���8�%�L�/I E� Ͳ��L���L��hTW9S�Up7(��`�u��S8&ۂ�{����+�]^L��Gj���=����y'���6̣Yt1��Te}�T������y�u�;�υG�-��( �����:�(�]�f�~7c��NdT��{��&�ix�16��`݂q�x��X�"�IҚ�Gk�өg���w��O��Z���(����4��	��Z���~LYo���	}GVh�:K���=�UXOO�DN�����1Ƅ��/��~�3ZF�Od���Ц�~���J�������\�z<ۜ�9' �U��.R�[3U*ޜt���3&�mL�1ޠ�&�|6�T��T~�?���;���F��A�H(���ӣ��ѧh93����� ���l݇R���E�ɴ묄��fW Ж�h�q6��Ti�Y�	�H����9kpK��Q���{\�n��~�%&Tc>�|B+9�c� @�n�tU��Ѐ�rQ��CN`�2��,-5���U�7g�J��2�\?���J��N���b���j�VpOD���/-v.��6�75�o��sZ��J���E�^�ޯ�Z$s�J����%l'D7�~�v6��D���aj��>KٯE��'15GN~���Mt�������8��x�,jSg�4����fr��XXĦ<�����l̀;%����q���Dl�!����)K��݆<v7�  ��Z�<dQ��B�7������ٜ(���YUc�H���0���pZ�f����!1c:d�J�J�W�U>���v'R�6o����C�H�0QKJ��@�L}l�.��o����phm ��ÏO���.�^Ps9�?&)e���1t����Zxo�8O�G�yG�"�
��O�^Y�{�nR6rO\�;8��x���r�Ы{^��s�dc�T$w��T��X`�ة{��χ�K��>M�k�ZAd3k�ɔi���4a5��	o�ǛVk�U0=3oիDA�~��҅���ɉ��ذ�9=J,KtN�g�U��+���H������'�%�f�~��'Ӊ�B�{�yVF��l]��q#r��>0>Qc�ٌA��MF��s�+��}�8�ƌDVr?�UX��I�o�7Eb5��&�� :�L�&��3r"�O�u���ޓ�)逰�只�,h}�G�w�:�x|�M�6���*�P�:S�q��#=W0�\2#�?��BIǳŖ��Y^����h`wox3&�O�T�Ja��^]L=�4ت&���y���1�q��2���**���G	�(Ggx��_���m4��^pn.N�)�,�R��#������-�׽�r���݆7�2\���+<8��Ļ/�B7���˘_�r<�;C����W��牫��O�V�)��ʁ���fGm1��W��KM�[u�ە�1^�eD��X�{9���{�������c����.>���t m�O�&�SnX鲌H�M�P���qN�pXv΀�M>�;]=1/䨕�0Ѝ��Z�ݴ��+_�� Q��,�Yp����;��?Z؏�o~$���궻U�F��jT�>i���>~�2�c��M! ��؛j�n�z?�A�ތh�<yE�y�pJ�C�y������"E�\x^��+q�}������Z�fˍo��L���/t}� N?�6���Z�Z�޵E}�s�Q�Z>tIo�s+��v���bE�>��֘?K�"6��/O;N�]��s�!�,�C}M\�Ƃ��F�j	�Q���-���4�'�;�5�V6(Y�e�k���U�PZZ���T�|�ӒG�E����fCA��Ԅae-��:����g)�_�~��k���nگ�5�v��x�ǫ��)�	�cY�#��"��y�&Jǩ�¿dVA"dp�vj{���5����Q�<xF�,���@=�T��i�~�]R�3y����ꔊ�j�)�A#{$�F�/G����q�l2�>&�1���#x��M�G`p�w�^(h'�B1 Yq*/�[��7�2��p'���+Q;56�������o��&O�������]���3���ڶV0�t.c���/ަ/=���e�+9�A���;���|J�a�3�z���S���-X���f��O��I6}�n2ԩ�[a�7��f0J�7�NJ��,�b���e>Gܣ�6rx{���]�k$>YE�V~g�#���Ja���`�]��-��"����>�� �U(�p
9+��U���t8N�H������m6p������3���c	+�=ѹ��cal9u}-�)����;�V��j��b��Kd����ݧ0��?��=�܈��g�rn������o�s���R��@9�U���P�G�7v�-��/�L���%�-�8r���Ѷ���#1,���3~p����G26�u�o�
�P�
��"ܯ�L�ı(�5�"0n����Z��r*�qAӃ���΄�*l�t7[�~�#D��\s�k��?M�LB�0](�E���Ōa5�m�c�R82�
c��Սg$;ȼ����
� �;
�,h�����!3Xx��N�ޕ�K$�,p���A�q��^�D���N�f�`s��9NyМ�H0��/c�A�x�D���g�Z�6�;��܁�MaD��m���Rjm1�9�-V���%��[����%�0����F��3qj��'[�QSg!;�g7���qH�헾���Z���E��s���m8W������F���³hW�����{�r�
��J� 'm�l{� ����=
:�U��e2H�c��k8ܲ�E�`DЇǿNaK5Q�o�"I�������ob��q��J��P0V.O')�bq��(�Ҧ��q�L�K�k�>�yR�]���>�˽Κ�M^6n
&uUV�������}�M��K�r���[#GNw���Ӗ�F�8�����1�F��7��E؈t�1�2GU�zE�	R鳃z���h��й�F	�X�k�qc�1�I�����U��C|�w����}:�4pA�И���=�����glN�Q�)k2����,�W,xX8�U��v ���`�ŐnR�:�t��w,-���lO�v����;	l�����zU;�+��C����@�bk�Y����9����n.y��/>��Bª ��݇%���uWܑ�U���-��U��D���wp'��Cr�0�<:�c;�� ��ȣ���]�t�ߠ���qV����G8~��éB�(f~��WZ0��Ƿ�#-����A�偔_��7RzA2�}��,0�C�?�.���JX�pD�p4W/�1akM��p
�l��P �Ē5���hMC6�\Qs���k�|��L���^��K�J貂�^<��M���κ{�U����?�3��R�H6샒[��[ԍ�Bn��G���=���P����t�T�����\5)��^	���,�#�g!�(w�,�o���c��^C'��-��`��+�1���}��ԻEH��]"�
o�ʤŜ캩X#��S6��-X#0��E���8��7zȝe]^V2��s���=��}����GXt���7���x��h�0�a��H�DTԳ���<s��� XDX�;	
RM8�K�+�{:��9�&d�:"�,�(h���9�#�7|���\z�ց �sy��܍���7�g���.�!0������RX��K$t؛'��������y��
A>":��W���ځ�2�Cu��i:��ɮl�v/g4h3`0��3	ڟ��U)�$W�O�B)��X:<XN���H��&=u���x&����V_�����iM��@�ZRkL�=@%P滚�HL��g!#��ǠwB�)|�[*_��7����CK��f��zC��tN����"�v��ٖե���I=F �Z�|��?�=;��K@h2�A��\��ߚ��#ua��f7yj!i%���ܜ��a�8�X^�?��:��W����':��+r3Lw��͋5���fx9S�&��UrpY�c�J fs�=rI��y�/���_n:�?�?٪YZ%��UC	nz1́}�VǙ��f��>a�P����Gm�a:L��E����G�n�p��' ���S蒱:�k��,�#��z���zV��A3�=wB��â ��~�����Xs���_?��ۋu�8f���!�jk�A��v"UDf�&�]d��9>\�() �R�9�檏~%��w�����a�w���ɐ�#�v��;���]#T8�=*��)./<�Ծ$r֕P���35<7Kw:=D�,��G�o�F�;�B���J���`�+�,�G/�F�#��bF\]$y4��+����Q���6/t��2��z���C�X����`7���t�0�yL�Owiv�*���� �� �����	� [��$��}t^�64��JZ�0$���U�~UUW�N�M�&P�w)�:�����e( �Ke�`��:�ϑ��gc�f�ݰG1{*Ig��U�)]����҇_ɭ���)v�a��)�-H��:{F��h�� ����-�٤0æ�Ks�G8�3��)�p��]���Ks�6��,!sJ@���겧�� F���[�6�Y�͑m�6��-[�!��=�bX������f
�t�������7�<������[b��P>��(�T�{����q#�B��u�N>����}����ݔz�N�86��.5=��C?��Q�
|�� P`�?��T���?���	3���ș|�->��V�P2E"��k����*����J���:r�~�Kh�Q2:7����q8�<+�n���@^�'L�- X|�Іo�zފX+��ݤ����J����zة��̌}��	 �-�;X�6�[�,hSAԱ&�@�`�ߎ{�/g�E�F�u}�f�����T��a3o^�<�..ȿȊ�ߓ�x�'�ܟe3�%[��Y�Th�)��`��.���y����}��j�S��meU�gmM)���+���d�ۆ�C��]c��F���������9Ǆ��Z|�e^�uBކ}��2z=ï~6����6�Oy����;���8�j��⌈Z;T:��hz�$ZZ	~u$��4��F���)�<B3~Q�x���I]
����pn4��,c5kU�Y�D�X�'�Յ��Q<�x����*�z���nŨk�u=\��k�����_��B`6~\�4����67K��Hu؁	;��Z���������G\5�U�(P7D��ߕc���m�w���Ī��2�� w*�pQ�#�sy;�ݼu,_|��*�R����N���#=&Ȏ��2H���8s���6��(L2�������(�qA�-��.�H|�������1u��K��p���4)Oa}U�w08�m"G=��B�5��7�g�O��I����)#��Oe?Ly��b��K���Vi�C�8���X��Q�n�&^(��`b�~w�ы�m�׏�W�Z-���B�V� ��RA��8�5���F�&�����#�X*�����[���a����Y�� !Z��3�A���UQ�t���;��ҋ�f��� Y����T�*�j��C�� w����8(c���#(�u�UA%�F������Ht�b?��s"8��V2d��K9��o��?xTE$�$8x"�P�l�3j�z,�uB���e�u,��yJ�Hj[U8��N�@�Da����!:���'��YU^��M�?Q���$68��4d4�y!OW�j���P�eaY��uu�{Am�iN:���tH���
\z�!���$�'�lS�j�@�:���x^Ҝ�*������a����3ޟ�����Uv�oF���(Re�ɮ7�{:��e2z��� �V��l��S�unM-��~1�����zD\kN�p�R�]��+�̏����F���@~�����L��^��
�W����8�L>~�d�Bx9��8-�$2��Dﲉup��%	Q�?��:)���Y8�����؀߆BunȎL(��;p�:a	x?�s�i�5� ���W�_ԗL�;5�o�7<n�tM�͗�j��$���'K�/����k�EUA��)%�'$�1a���]�ئ��c��T�w�Qj���2� 9y�O�K��@\M3�}�f;���cH,e)&Չi� 9��m��u871t
"�ܠ�6$#���p҉��oe)��J}�	���
��&/����c�A�H���9Օn����d�;�݃�j�1�W����?UV�]�m���徶k�c����ͪb�W|��xZ��F�'Oּ��ܨO�Z�9ϫZLd�<]&B/k�y����s,�`3y�^�� �I�f�|���4]ǝa�Ĭ@8�=�x��
^P�n��|���r#��Jƅ�:Q��i�;�:sߊv�-�#���a���|�1l�,������K�-�;?l�Ob��6
��:'�OD��#��q�W��y��/��� ��!�Ė���Sg9؆�˼�HCb��4Δ�&i��0��Q+&∯+gfӘ�����BZ��I}�+�-��s�]E*-����!>�I�$��#��B�F��(
�|�	&�V�ֆ5,��z�:nq�։]�G��cRT������R��J��x"��Cw~�t��0v�3R�v�u4��8z�@�%�+�k���H�N�˴;"���}%�T���a�/�et,&t�A⻌�2�؆�24HA��c*Ν]��8�~7#-�%�����S.r��%��O	��* �v���hY�"���k �j��!��l����EJ�kk�G��̔X��~+�GG����R7��(���)�&^�$�#�F��u�5
M�P���G-�����&w�[���uZf�WX��W�)���pE��ݚkܽHy+ؕ�GSB	؃�^1�8����n\�-�U_��{�^�%~]�Ns=)�ϛ;�1կBx�aC+8<.|,�f1�BU��{�q}O��1� �	���u���W��R�]fZ����Y��3,����w�w����z��n�)�;��4�ey��{�t�n���gpf�[��.�n(�w�oF�I�͜?|����j�}Dg��7�AL2Jw�ͦ'��� �kn�K����X�0K��#8�$Z�)�xס��?�#��<�(+�/��R{�R0����\�l��B*p��Q�U�U����.�N<���o�?����w�#�V@(�LTSL\~1"\<>������ԏghN}Q�j����� �i:���M�����e��96^=|u�(��k��YRu���2�-��Q�����������^�GN����H����M�td�0�UY�5F%���i��=�q�Y%� @�.Ԋ�+t��^AVc��8�����(M��b,���cU}2���P����dؠ�ǵ(�鬈���^hӰ��ei���G]��yz�Z69���j�-P����QG0����ɽ�Zf)M��h�S�g�*.���*���CSNQ���_6Vȥ�>F��5QX�ٹ�����n����VӶ+�*�����Uto���82"Cq+��@�ۨ|��o].N���m�[b����{�;$\Df�����w����U<wE��X�jĦ}��²1�kp���M� ��x�	7b�뢅P�%���L�p ���P�bc��%��B�vB3��q��c���>g{�lgi>�8�ر���&����40J����tj~����n^M��C�5��V$���KZ��)�~� ��'%�\ ɵ>��j�,O��UI�=8�N5Y��'Jd�s/���h�!��̀�1��b鲆�Sj�S�rQ��k���L���'��p�1h�\{��xgmoMr(m��ʻ���AX��5/��#u��ؿ�`t2ӑ�"A����Ti|�71�������,f3�o��w%@��:�x������	!������8�b ��u�9!��/,@�C�v1��	�ʴ�&Z�H
$ش��8Ɣ19��t�p����-�tj<H�oQC�oM��wN�e����g�Q�0��$�T2��n_�2t6��ƞ���G"���A��/i�ង눆���q��+-	/7.4�L�m�L��M=,���@b��9��Z�������B�8��.[W�`�и�ۇz7���
��Ҵ�:yn��tw��?�PpG�,w_vJ�")Ǥ�,D��6���t�2t��ّ�8;��D2��,kR����
DNݮ�T-��Զ�A�ҏ�i��d���ա��~Ȓ�	/���g�� ��r��!�BS`t����!N�}	u�� b�j�.P���k8�\���0�:T��5���o(�����_@c�;Ţ�X=֧�>�X�e��n*���
�=} �Z�"��������#�ԋp�J��y~O��W%H��+[p�-��l%H�g�P�a»���I�T��k�8� ~���N2m�w��ׯ2_��wC�%���>�d�x��M��ǥ_% y��\�a�vxg�f�Z�;�@R0�5uU�Əp��W�O���o�v����v�f��㿼o;��>O+ՙ�u��[DM�h���^�{L{��ò����=��nmH�l�0�����m^T�E/�etیP&+�Ӧf%�.�6��0�c��r���B90���E�����˺6� ��� Ѣ����mز�$]r���zM��`|&#L@��~ϻz�l����_�J;���������1��( -<U��^+�aT��YE��p�2�[�:zVL�Ə�������P����x�gI,����2�X�b�DM�~��;@{
��ڞX3��.h3v�sN��","V�]I��Q�@�����@������ ��G��DfJ�%�Y� ��Y$�����2�4 h��,�hj�/U�����e���s���v̜�{ZD���\�΃�7���d�2>Z���)<oP����)OϮ�ER�|���{_Z��q��F׮a~�ƥ�����Y""����?z�.����~λ���j;K��ķ�����Q<�լ�7�,�G�UC��5B�����g��-nϐ*
*�>���RJ����n3���V�JD���_BRm�Z�.��҉���h������Ew=��{G8P�X�|�/��k��ف
2
��X�������;�F��H���3�Br.ƙ�ڌ����v�����o��ɧ���ޥq2�4}����E��ƱW���`sа���;�D\܏��_I,��ȏ흧�"v��ܤr��y�E]X��]d6Ԗm�y_r辨U>��Nx3Y�m�^~|��-8(v�U����?�t<�}dq7#qJ�\{�,�Z��6oN�dw���\i���'���ڸ��Iu,cDG�4�V���L��yl�-c��@:Ϧ\�"B�hb�m����Ky'f �B#��[Ml���p5�0Kq�;������rH~5����T)|���-}�F�����S_�Q<C�0M��)Bq8�7��7�1�呚�|��bu�� ݪ�d6���m�0����]����d}6��{��}�y�����Q���y�O|wrw���R�ȧ�kl�Nz,� -ŏl��%ڳ��'�oN��ւ3�.8��u�F'֔t|
�}:�y������x��j�6�4�@O
&+흳��o����KI��oF��4����\X=����j��=�H�k >{19�>:���n=�yd	2��K��Q��|�{�"���l)���_���Ʊ��7V�9ܱ<yD�9%M�S���-�%�9�D��ce�ʔ���,w�:
��$��kn2�Ccx�5s�k�� xTIr�F�=��fd[˚uS
d���t�jO;��q�g��P1�� Q��k�����5�K�Hȝ��h��3k��-� �*�^��5�n(u��\�4�.�ㇵ3Ԓ�Z��P���9��}t����r��0�4iٕ�-�|%�&%gV��Ҝ ��SB�;��a.,�������r���%�fi�T�[ H��3U��m�ј����c�GUG�����<�w��Y��!��u�w���<�t�����7�a_�����mC^;S��\�O�e�H_v45�6���B��h
��_�T�rV� ��A��*����aS�(MP!Y �	���g�T"(��g��9&m���Dl-�\bq�ܻ�x����#�<���#?�i�Ϋ�kH�-41��{$�z��E��ANR|�:c�V�9�0x9s=�W���G�L |�7tT[�B�7z.�]�7s�!(\��$Dz�C�Mn*�pz���H%�PY��^x(��ͦcS��k ��v �.S؁�9�y���zMQoʍ6NG�9v�#� �y�eO=���cLE!%����ڡ���'���Bg�aU��^�H^��=^U`|��*6�kf��L0����L����re%TB3K�1i��~�D ;��B���q���0m^�0�T��%���y��⼙�/�����O�p~J��a�g[�˒�D�ub��S����ݠ>:�����>&��kF�غ{\�
���T�8`�2�˚��� c�C2vgVVs/�\0�����,�� ���>":��#^rSEF�����zt���@���:���?�i�{���U(�>����a�뵶a�u�a����V:��+��GQ�9NZ�U���nW�R^�y6���<ƚkumG��B�z#�~;e��l
xТ? z/�%+Q.�J�Fc:b��rI#���0�m%^�������M����q9���ߥ������� �ۮ�-,���i�|{�ޖG9�%�&iǽ�/).�Ls���b�`�^	 ���T� 4z[�&M�f_�Q3�6^�M@A����oY��娈(V�$ș�ﺆ�ʍ����Ն��W�:ˋ���(�-zH)�EV;T� ����2�����2rm��n���{S�?�/�\�$3��ٝpT�e��G�bCnݾ�5s�cA\�oyV�P��q�m�� �6�[ʅ�Ù?�	O���9%,~��&mh_cP�M3Fm�4�3V�28Y�����X��nQ
�j�#���<+���r(�(�c�S,�D�VG�_���NYT�TT������']	�U;�0�<�n�lG��R�{�i�7����>���H'�"7n�XBj ������p/v��b8����Z���8�-i���C�HK��X}�D[�^��IuDr��\/Ӎ#%�`���(��`O���kԱ��*����d졁"!}&�K�-6��lb�D4�[�,葓��:�BzI��d��F~/`#�}��t���yT[#kT�'h�����%���O�T�$��ɤBߤ��\����Z�/�MXQ�+]vVח��E�"� 0ަ��� rF2�F��L;����5�)�7��R���Z4CL�%!u�i�/O$P"�����q O�d}��e��=�ZDe��<��èqj_ECcŧțL���9�mP��aѦ�l��5Ƈ�%�e`0���`S�P9�K�����zq����	��-|D�F7��*0 �����+������g9_�W�6�:���a�\Ba":RV����T#w��-�A�<��:җ�T�Y������C��r
@���޺Й¡=��@����jq��b�y)� +�1���t�p�Q�5o�2	S�!0�r��c�$G�:�����GO�����UU�fS���`���E]3�������o?�%�!zp��ߧ�HZ����3�λ�<	�H�v���ʓ"�i�Ȁ�����I<l�G�si&���? �%gׇo`��~EII0XyH"��%� [aڼ��N�0m0�_h��V뾹�f��[>�0[��/zV����@"j��I��U�� �G.�쇤s�>�>Nz	&6���aܽ�\9ht��i~\��حa�=���Q�B=W��N�:]�5��2>�zmE}[w���1��lH��ϕF�$7�����:�p-���\�b�O��8Q���;����(�����f�g��C�V?�W�]�5�b���O�0�G-�B��}���R:Uɰ}� W4W6�{h<"~�D���pr8����Gc�XY?c~��۸�t�"��0=��>P�����N!}?����N��|��R"���uy��3�pv�m�y�7?,�mO�Vٳ4?�nV�	�5�X�Iz���E\�>�� <\���l�%WB/�.�æ�g��\����e�]��<0�)�ߓu�=�o�8/A� ��B�#h�4�(S�Y2���%�9o� ����$Mz\���E��t�D$"Ys���Dan4&�8m�n���i�Ft5l�zC���5b��J���y�y��-l���^���.w�,1��Q�"����*Ms���V#]����We�ϸ������I��PGKOה�'����u����>�2�|�'����L�=R4mW�F�!���Wj�s`HQ���S���k��#��/�Iu
�F�����=���{��R�OX���I�}-Ki��LM3��do&M�鱑��j�8У�X�%�������[`�x��ԧHH�3h)	�H}�r'O��H;�>�6/Tr�B�U�7P��UM�u�uWջ�EY�T�f�"p�?�w��a0Ɖ��qk�Y����s�� +P��a��c�$��6%2��Sh2����a����x'3��')�L��� =�*F�� �L��~��'����.l2�u�Li��n�ȩ����iK�����<#���䐸#�L�)�l�g�C��ކ0.R[pG�B��h�!e���7J�\=�{��OI��]m���Rβ>�/B���u��rX��	.���	�:=�������G��|.<��JD��������t6��j�	��2A -99����G�gd��L�,�J�����8�Iz:K�W�:�����?+V�l�Q#�5*�-4`O�X.������e��/��k�F���p��)���Ц�+���Qc|�L�8�-�f�[��M�'���jQ'N�t��U�h6Yf�s	Y�1F�!�L��o0q`����{�*n�o׷y�s��.抺�3�/�
9E�<�HB3��&牳eY{�Vw�n3�.��B����+K�U߭�Q����{��5x�
a���jI��{��O	 ��o<09ּ��.b��w��9�w�Ԧ]v��/&�����	N��z����ajɝ����HOC��mQ�X*��O?�!R�\�y�]G�z�0����?�$Z��w_4,�ʳT	N@f�������o���qȉ�K��%��ޒ)��B�T�!�0 D����F%�TX�#?2��)<{,�n�7��X\J�h�`��E�NN�����;!��&���[m3po�|�	q$Y�[tn)��Ʉ��en�&��kGì���W���S�a5,������CɀVO�sT-�����}P6�\�_G �V̐=��\q4��u�zs�5}�I��3�5�n�Q��Q^ޮ�2v�j�38�Z8��+h/(-�f�((�>F�</���R�Y��6������9���c.~��Kj��=mm�����n�B�ԃ�&Y< �p�t vY�NM;�b�rx�S�s@�p �y.��FJ��y�yUd��^� ,�#�����P�6��iĮ�`������fN����D�oh��WSa�Fqa�r=�ml��q��g�c��3���^�˛��g+�yѝ���թ�ȒQ��Տ՞h��`2�Y��
�Zsףq&0w
JBH2�G�o�E�Ɣ�`��>���Q��)��9�c}b4P�x-!� ��U;�;��Ja��?�Z��Y���։�h�o0W��uM�mv�o鼊5���!��r���ή8��4-Bw-o+ 5�t
��nߔR�F�fv�'Wӆ󵩙��चb�S3��$�V�ivķ�gYǸ��J�n�â��E���aaDB�ԉ ۺl+�gK�!/҅䉎�~�u����h$7�ZC��.ڝB�]���3�����1�̺]�U���}2]�\��d��%7k���;`�tl���\/�|C�l��u���7�{��cv��"p$Jh��V@������̥^���N��n})a��'� b�w3��`�$=�UG*xX<��!�fCzd� ��`�F���1ُ�Z�xO�����a�!���� ��v��J�J��6���+�7�PA�����}٫&S�(<�����~���Kv�r�J
;	��G)�(��Pd���u�E�H���$Ou���.$]���!�`L�6�<,ںJ肻�-���+eO�9�I�(���D�[�������h*Hi"�(�M��c���7�v����Az���Z� A�.?V�]� "P������Jϕ�t�|2s��,!���J���73pK�4�O����r�
Z�J�(��ڝ�eb�%;�򑨯^��)2NQ�0����
|��Mi+l_��av!k,y��̇��L��
�.F�:�s۷��-�o����&SZ���@B+W�,��z~��Y�	 ^`��2�W�����=����4�C�b�S/�1O�R'Tվ\Tț���IO/������O.!��a��;�E���sh	�V������:v�]��C#�;��o��o8�9I����X,7�I�q�#ؘr��"wQ�z0'_=	�V�_���n�E��l��T��2�7�k�9k_(��m�3.�WW���� ��l ˴{�ݖ4% |'k��5#2IN�< S\��0�!3�'Yq�B=�sU� ��:� Aw#�*�o����d�Q	�}\�
L#�fTu��} �cOY60p%b�\L�Y�/J�"暐j5��~�+N�h|`�z35w�e�&��1�O��cjm�d�Fh�N7�{�|��i�};�ɺ��*�l'�ɇ�lj�Q���u�,֖p�G��Yz�H���X��I{! cQ�ܬ��k����~lH���ϩ�d&X�xv.� ���J=�Ǽ(��~����R� �F�� �5Rd0�r��VRs�r͢�������a��x��G�I����I��3���?.�YT�]���bR�I ���,�a-�}kj��E�x�бEp���E�m����A�@��p�;�9��fW6�8�U�^Q�h��8���E4S�%L4gF�����B:�b7���6��BF�)�Dh������G�7f��{$�N�*�~F�K����%�Jt��h����J���Y�*�#�G $�<�*"xx�Z�tU���q��Or���7?m25�2���Yc\�РgK��, �G�� }����y����uȩE���=��È��s�*G�?M/kNg?��z���r���
r��VE|��~]Ka4Ͽ�-1*kt�Յ�L�:+ �@���8�����p����4|���B��>�f-^�.���a���2EkL3X$]舓Ђ2�.�;iG�гbEr�Hd(��!���KyڙSǴ>I�j�n�Tl����sW�)Ǭ?0�	� R�YS.hLb�f�
y�9�^�|��R�4���`YGy��` G��~Q����mar�7�Bk��	�=���vj���Q��>.C.m����&4���D�̤�싚J ��?$�QT�{>��^0C��2�t?CB�;�R&-�s;'=�i��1�aT����\���
D��e�ӕ��b�_߬_0G���;�*λ��
�͏�p�l�ȼn�;�!*�9T�j��Var�{4U�0QDԊ����>Y7����O�����N�U6ƙ�\�,�'�r5qr�U�"p0��
�]�)����07�^8�����h�x���~^�ht������V������K'[Dǥ�U0d�����s����zE2�&�]�IhH����¦�2��m��%� u�]?6�����wu�>Sq�cY�?M�ZE'7���W��=%c��z"]6�9f�u�$C�a�yP��|�.�
ۈv4?�;��R���K��{�]����#��2���"�������1������PP�b�s~9"u�Z�*�p��JM�&���?�V�TT�+�t6.���p���I�l����Ó͠���!*S��a�HPX�[��:��z)�)�"t4��.v����T�*v_V�S�N�#�6�L	�U�˅�4U,ws12���̌��G�>�����6K��/l���� �k��,��x�$�r�}�(�z���xj���b�,�r�IM�U��#��{��>�K����TX�O��h=�R��!�~��@ˇL߆��]}���;˄4<�E�m�ݷPW"'��7���Q�?�RW���y�v��������~0a�Bɔ�K4�hh(8�H���K�eBϩ����+��H>��D�ya��� �l���z)���d_��"�ȃ���;���j�]s�@�p��Gi�W4�٦��5��J�-��[g�G��Eup HM�E+�c��`pU�M��3(sg��B���s쾿��W�!��~]�k+�<I��Ys�=
ȿ�:�3�5^z>]�a��0�����YN�Er�'��}��-m�+wN}�xq�P�Q��M9>!���b��N��w��ˌ��k?X��2��4��V��Lv}��a���0������8 ���ت�N\*q�x�T�Sx�����dt��f�nE��IM�|��0Ք~r]�}v����;]8����xaN��R��m�;�3&f+�����J}d�?TC���{1�:�ުF=�|��P��w�+I�H���J{�� ���	����<�"����(J?z
�z�Tj ����4�.�.����A�Zc�'�=�f��1Pu���!R�s�mKCM.��hh��p�_0c�\h��@֣u�Y��<6�c����[xk��0M�1ш�*�y �`^p��6q��*��&��#���(���[��3@! |4�K�{�?��(�����Q�j�c�`���7��@Bn;��� �v�K �2A���./�?�<���t/d��Vv�e�G�Yv����J�es�J�� )VB���Xm����{y��jJ&��n(��F,3��
�Vt/��~,��IH�3Ȗwg$�s���c&+?[�-�]3��U�c3���tW�cN���Z���+,u�������mƶ��nYN�_!�0�kx�Ȉ�׹���_c���ξl�2L�#_`����OSf���x��	�Ҁ����ަc�M��d'[_i�����&2�SA3x�ܗR�*q3$qs`��-H�Eb����?e���t�����)\)��4{\��-^�ޝ�*%�	8�/��?�$.��6���':U���6͑0���\*��w�W:�gDڝ�؝m%�U� *���lTh��7�z�c�	o�Y��֝g����f�r�����<�p�6�m��|�%L�׹�Q@�i�e�*���K��-��{��谖�3� �^'���nծw~�1��`��O�l��9���9��S�nAg �;�gE-��2����^3�q��	�QLV�( ���N��#���'�]���z���p���Tbk���(�yہ !�-��	f�~��A@�M�i�i���fw��I���^��=�����td�2�ȣ�lm�$_h��Z��1	o N��	��a�,M�q�V�S��y�����Ŏ_e��d�3̱�irh!r:�V�Fط���s-Ŏ�%ft��,�4�b_��CWl�(Q���u
���IP)S-��;��	�q���߃	2���5n�@;m$
/�wx_�}�xA>�؈��grij��g�b��<�K��&��7L{�5vrǍ��͸iU����g�R��,��"`�A`�o���9yqDT�-��<)+j^F v�_S$�����y�%����o�@�g��FN��Q�X����0�0q��\�(���͍}៻YO?l3h��70����p�G���zB�*�Oq����8�@�8kʾvV����Rkz>���0�r�vw�p�������RV�lk��6�f����F�p5�=��)y��"�y��b�8�Q���62!%�'�MYO�����r	?��c/*g���)Zo�# �6���x��?5���p��YmZ@m\�V�1�ͦ�^��9�:��U��%t���qEs(�u���9�=��p�r$���k}ڥ;(��ʋ�)�9{|��K��:d������ס�3�[��xB�kUwk�cR����m˲�����&�c����ѻ��E�m3�����De'��~
�^�3�5 ����� �wb�EWPu`��%�R�O�-ZV�[��d����}}^���E�t`2�Duq6|0<q�F%h�y���yRtD�'q�@AfB]�G���NP-�%�g�*�^�T��Q)hڹ���Fs��ZC�&u���$2C+	�� �My�m�l�v:]�F߅]�rևa����I��%���Rv��>�#ı[%�:u�	K�3�<㏺N���jA1����bg�cս����.j��`1SSb6`.(���W�y��]���ާ�@c��V�M$^?d���8�����1���R|۔�����._�e69�U�4z����i:��1�ȼ��K�o�G����s;�4�SA�b���&�~)��QN����$��\�t�PmE^"hw��@_��]��m�z�B��1�����aKv��S��tX��*8��G|[��r�j�!��d*�f6�������'�ZǅǶ�z�J���A���2�)YGK�����-�)+��o
��t*O��m�����=�X�|�l
[�6@��x������i��p�B�~]���F��{�^�������;��J��M�_v�F)P�����)�q�pkðѮ#e!e5z�#2v��2�&���VC��B��ZK4�*����
��C5������uR�R>m�Ð��du�L�����	��˕ȑ�ݢ���Uq�]��7�/�G)���C�z��C�r
BJ�E�~�|�H<#�Wf�^i�`%���-�Y�L�j?QT���+�~~�/9���]��̈�?�������B�^��9E��4�H:K��$&$��?.�զ`0�6�E[5Lu�ѐ	��݌ࠊqDr�Pv� ��!p�-�DP��X�n�P������j~0��Xΰ�;��*���9w�9z��H$B!��[�V�t8��+۪�'����noX��d
/��8::a�=d,�+�4%�A?<#M���h�ѽ��]��{��w�Vj��s|�4Np������p�۝aa�D9d�(�g� m�qʖ�k%���$�B�2��uH\��A��v;;��)���w�Ң��{��ˇ].�:X���9�����r�!����e��qI�C�!7��$��T15�J�����8]�ϙ�T�@�G��Iy"(�0}�����i��<g�JϞ���)F�^��~�n8�3U��EP����, �]��,�}ڧS�,I4��\)��{Ǯ_�݃�B��^S�Ԛ��I�j�Pn�^�2�[d�q`�L�ݴ��%n��@�@hf��'��$D^ϴ��d�BPf�Ճ�p��dN���%��!�i
7�w�.�;M��I��hy��w5ZSΉ�f���Vk��_A	Bҕ�%YR�'!�9�r�y^fXfc�wnзܬbթb�� 	X�
��I�T��F���U����w��o�%x�1yJ�hc��'����=������,D���f�#�H(�烒��PF��y���U
-|�벟;�õ-�M$)	d�緇��J�%a2��l�L2	�}Z�5<��\��7�˶�k� MX���T�pHj����e��{�]dM�0�_QW������'�;h�з�D@B\L�LKn%�P�)�V.B ����O>b@����-�k���ޗ�<�Ԍ ����gj��Я�]�泵���Jf�h�7�^�P#-V�,F���%�g�a��z`
!g�J�w"�u���sqiN���H&��`�\�2�2������Y�鰽���$��@�wO�XI�O�����WU�Bw��Y��r�F���n`����*B%T��:�mXt�Ru�6���I��@����G��0���k7���[v���W����nO1B��$�á��˂^��y� �;�Y�������K�I�5X�M�G�$�L���S�6����Ѻ(�H@[NF���2�o�Oʀ@>�_?H�FN�h�h�@+�k.�,v��A�X�,_�f��������q7����gi���,�훢�qm���L"�+���k����yxqmɇCd.\:�"�v%��r���Y�[�+q�Uz�0Tf�JV�/}�^���$Bm=�nKF�^*��2B�ˉ�!���0��`TY(#'��x�uS*�S�(g�]�x=��UB|��\F�|þ�X&V�a�e��&@���G��<�a�el sH�����WV�w~��C�L�����q�8-�w�e9�]8C��&\�v��F}[�\�Ѣnp�(Ed��F�h�"ib���~�s܇a��P���t?�q�kS��M�bX�i)�Z5��:�g�w�v�-�t�����u���vƘ���+�2�Ɇ��s�ɘ�2�~@�f�ժ~�K��8{Ҧub���S��sjIKKw%�w@ �h�^J%��X�����/�A��[�z�x�yJ鏛R.%˛ٟ'�tf�L@9D�)t�<�	��F���pӖ����Xg�b7\���b<��� +(.\��Zw����88�F��F=��C]
�$@K�د��)��Ձ�7���C����" ��7�	,m~�HJU��7��>��
�[��2s�9 $��[=�PCfV�MB���蒄Hz�@_�	�Q�G]��|g(�{��ᗢ�'�
�ab
�.��v��-O_��k�U�!� j(�RA�pO�չԝ�gdX�r�l�L�M�8�+�3�i�]e��v���}�&t���+�������0%�f����]B �n,����q���X���gm������1��k0x骆�����)Z�=�h���V�܇v���Ȇ *�mh�h��а�G�	�a��_
�9�e���fmGc˛BcT6vK��c���#@�U_��Na�)h��kd,f�Cl��q2��	�?��Zon�&��g�����o1O�+�v������z�sd��Q/9 ��|0�5��������m�ۺ��j�������Yd�JկaR:C5�&�� zTH�,�w��uf�$���]<谢�Իa�J��
�m?�Ƒp+0�P�fԙC~���e���ۊ*C�"�*���骮���%�-���x �O������[RAd�����ή��`
h}���� _��ޝ���#�*���fl�siD�i��8i�|�g�S�H~{n�x�Œx��:�0JcX�k3��#/�m�wW}<琊\�'�M��&�:*�<_�J�c?�F��_J�Ň(ֳ���F捘����}ބ�( �I�橼;���8��7rq�9jM09�Sy��7`x=ڹ: �����z������i�)��Oa�vhi[���z��Sأ����ݸ���fZXE�ZE�%���T���s�����T������ɰ9�m��"��&5g�:3��1����y��#d>\d�26+�qZ'�������_³w�99 9�8]Nd�B���el�R�#?�hU�*v�A��{ָ�/k��N;���Y���Q��xfr�_W���4x�w.KNd�C�A���T�|@_�!�l��sh�p�,���D0���_`4��ET��V~!��aBA߁R�u�w��$�fς(���bS��GN���&1�u�&�t}�W�������&�Mƣ�����5Z͛�y���q!��8�k���t��ܤ1s�6"�xk:�w?w�rx�A.K��]�(�vr��<�kwt\��q�mUŵnM&-�`�ل�A�5�(� �]�v����2ly�V�g�;._($XsR˙W���������l���l����:=� �����ߊx���~:j�*��߭�^��z��&h��+"bad�eX��[3��pKy�
�1�mFP��8Y�"�}��J�MDGv���L�>a(�G񦙡7f�q�����\��b�0n�o�L���F�����/(�����ޱ|Y���?W(���P�A���ܢ�3Ɍ��~����p��1<U.4�?�fiES?0���xE��z!,������p����W43�"S=�cf�y�����տ]��m�@����m���kH�n���&��uO7Ggi��cg=���d;t�ݻMK�-P9'���M�������t8�߃����9ޓ��ށ���8�xl���A�p�-~�v�H��(��"ؤS��TG��*��<���%�  ��e�d������)#�m�`��J����0m䜙k�3ۉo�f��	@-�{ /�Gp���br�hܹ[fVYa> =>pi�+#��0`�NoĦ�OSq(
<�;��%��jwM�SޟMtgR/�CC,0O�ϙuGR4�+�}���͸�����$3�:�f�`�٣+ס;�Yz�Jݙ~�^iE]�m6���1\�G�`;Ä_�wJ�Բ���Jt�U	L�p�@IK(5r>6-��VT-\y�\j9b,��9OQ�Z$�AZ$����.�Ƈ�E��vw��v� y;ڡ�I3������f�g4+�]�B�u��Zp�c��N��
�� �'LK�KӒk��.���Ѥa�ѽ�{S���Y��=��hT5�:섹5 ���Y���'� �뵴$eU�5w��_̄� �Z����a���,��a �Q��\��=j��U�E6�
���;3����
 7�7�.ù��ǻ���.� t��l��em˘��U�Mf.&�;ӌ,ǎf|���-&��&U�X��
 ge����/��:���9�hu�JF"?��!k6�X]��FRHa�Uˠ婈�9���tl`hk?��\f|�X�Y4���u�<;�R�;5���x�������Ok�����Ӗ�}0�HI�P�������C�(ۧx��S��G�~ʮX�L�X#��ol�;%p���,���J�7c�d�����|O����q06I��R��5��-��4n����4�@Rp��|ўE����2�I�C��m+�_�� �Ϙl�����G�Lq��&��rЊ�-��#�[��6���'Z���P�y}���j�1�nQ�#sqT�?�C��	~Y�s�YÝJ��]��x���f&�­};�q��	/�!Yi� �iP��q�Q��1��ߨ���~^�Xb��B2�Ձu���h�O�*�9�OJOoX$����`x%&���t�Xc4&/TI���K�{99�s�b=c�o�|'C�h`�k�B��\�o]�����#}Ą$���pO)H�*�$�"��2��+��[SR����6��`���W������M�d�L�w�j���!t�=e{a�KC�v���b=r���g��\�3�!?a�[6�]�w����F�Z-�
���	�Ҹ��X%���ۧD��.��{�T�G3'DE�����F��V7� �őI���Ҩ9\B`��'�fK8r�
�@� �����I����:���,m	)��94a�2�ۼ&�h����5�C}ʨ㌭}��w؏�7-��+��Ɛ�+��c�U���49���$�˷10��µ�3�t^�|�i���@s#����j���!l�M?�J#BQ7N��d;t���m/�R�����Ռ���NШ����[�$�
���K��lJ���'#H���x_�����C�E�������*�*k����h���s�Z�|��x�C����jp�=���`�X�e�	;{s\���~��i�6�164j�h�qG��5�C���?>5r���x`�>��D��݉Z�DF�Ye�=Q�]A@54����}vŞ%
��>�F7S鷟Z�o��6�b+�O�S���/���1�n��J�+OG�h�	�F�����JG���%�rЫ1���@���u_y��+�Y��>��Se���;��I潎om��z<.
��B3�� ��Adn����.R7�!E�GH�F�
1=N�?��\<�Qa��ܻ����l]�e9�-��E�j�~U{�5�u��.�0��(Ϡ>BԠ��G(lLC��u�ߏ��ɇ�� ,�����J�;mp�XW'(�m�����-�٬����PS/:��2�rh5���W-�DX������>o�_x�W��Y��+z�H"�����������X�M��$�q�:(�f#A��p�`�g�o�rmp[Xz��^Xjq�,xqmsj_L�� ׅ%>�	�[��x3m��N#F�Nla���J�z�^v�ӎ���fS[���F�'�Ǌ�v�Ԅg��<�ԑ�v����ˌ��M��iFo{ݟO	�Ñ,��љO+i��������E��ECr��ϳ��n���u������[��|$P���5]�ӷMB���gX�X$}�LhU�_1�~���6��g_6%�,F�ā�b!��$��ߞ~ǲg�����<m�/��
�w�g~�E^�d�'�(����7��wWka�'@@��~q Q��e-������.�d��
���noȌ�ۛvpi��s푾���O�-)���|�/�}�R09��b6/�O��w
Ԣ84q���Ϋ#G�`Ɋ����Z��&Cc���i����0��xI-��=vf���1����}m�������ŏX��Y�����,��ag��)(�X��,���X?�A��R7ߵJ1�l"��n ��w���:�%�	`<%����U�!�Y���Њ��|#�.�[��ըn�R��Üo�Q�s���D1if���^�:Y9u�d�B?�
����ߤxn=~�����x>�HA<���sR���מB%���鏿��t\�����1��[#���I�l�����TF0#�G���Y��~����"����ݳ��I�O�8kcg����~)����h�Rr7p�Qjr�]�_\���ğJ�Wa��g�����+b,ٗ;-Mw�KI�ׅ�U�h��Q$w����I�ٙw�������*j�Q
�Q�^m��<������lW ^�؁Q�M�rc�`��rۮ�4�I�BF}�]Z�H�D�J�	:TU�`O{����~א̤������=&[\-D͠�. X�
��ʹ��C �o@��y(���n;��[�۬g];�N�V���x�,�,9��H&�y�'1n��QQ7}�Q~Nu��Qr�L�|��:���ym�k�!�U1!��猝��_.`s�[0�u��Hȥ�og-{�=�BO�i�
�&�J�O�P�̯4T��t��=o1v�}�!,lx\-ʼV� D��nLi�˙<�b�JM7w7�z�����x s���<�_;`�rv`�v&�Qv�U ��ǰ�2C->۔���[w�\Dp��o����#L+�C��I��ʽC��y�dn�%�_DnC!��V�r�P���gW�+Q�!��d��ׂ���ϸ�|qZf�gF�uB��g��QAnW�91M�cPT�đ`�QiJ�&��H��(1�r��[�͟+鸨��
L�;`(����s�PP���_ ��a �/��B4Dކ�0�x�cyŤFq�.�6��|?�MeT�Q��TI�(R�si�!��2���j(6T~ob\*Z4#I/%����2��)n�*H�/�h~�����~Գ$W���es���΁����m�[E�6N�6�_�N�HO9�	�h
ڍ��0~�Ӻ����e�HT��u�߳8A�j�ק����ݏ��%4���~�t�\J��b��FA�ߐ
�֗�ݛ��eM�{M��J��<	��!��ԛ艩hg�2Ah9���ٱ�qA,���0��s�D+6��jM+9x݌[&�׫����!��?����㑕;��ߤBf[*�2�yY��7�"��r./&��-Gù �т�J�=B��c�����$D2��sS��"9zg�P�7R��0�Ť�Bn+W�!��n��=�G�B����2�ԬtA�)ή+���4� m�rD/�)+r����E�J*�I	7�r۟�s��1��gY�y�.lG�b�d� r��&����ǭ���ۮ��.l�Ne�xP�~�Ӈ<y)V�ܩ��T��LN,bp� �7}qH� ���s]����j�i«�E3<��$%|l�|&E�����ijV�~������3(�����iP�X�G�Jր����I鷚��>��~|j&�&�:�^��S�"�+�Ot��^A�[�ͩB��#�A(�T=��XQikQ������� r�&:�h�Ký�h�4��iPp6c�������p퐑ER�:a�J�[���$r#�٢X�UԴ�P��l�Kn�T���@'���g������+ݛ3�F⎆0���Cjb��Q�Y�&�=�3K�xM�n�3Lݻ�#{?z3�"���(����|IDr�fW7�����A�1Db�ل^Cw�
.��P�جM��1���6�CNF��VIP�l�$O�Z�w�zm��&n^G�P��I��I�V�?d��q�r2��r>�b,m8�E���P?��w�n�����;������6�-ȝ���H��G��A�z$�-����9\�}���e�~HG
}>y�l��䶤^U�^��Ka��0x�o H:�-��tӇ�a�4�H�'h�*�_@Dd�h�����C�LE���ũ��م^K:���JD8�g[e���<[5����;�>�
��m�>lh�i�F�Y9g;�y�C�����/guED�Gj�~���.������&���/��a�-��p�Y��>@����0�(x��9)��O��=�{Ӽ��A�Ql�}x,?2�N�\�o��(��
�W!_�#��e
�D\M���f�|���t1l1##3��L1���:��5���<����p^���߀f]>���^���� �-i�j�ۙ �Mw��u��Z���UoP��nR���{A�iz �NxA�Up��ȥ)���um�b)Ai�{	m���(�9e�z4�Ź��d�����X`�{�(I�/���t$�����:>�Ch�WؕN�V�׍�,������W(/�)*e6	q����m��RZ}��q�U�h�̶nT�ж��7n=��e^�"�.1��X�F�Ȕ�C���>Ց.�0|�xT
-�ىr��Q{ϦW�7�e��A�ipq*�Gw���f�H��|�|�����,��iNj�x��-�}��Ŵ]�A�爬֖���K������P���i�	q�����������ʹ�hڅpR(>�&N��j4@��?p䷗�Nܢhs3��N����q��UOv���w%���[N��W�2�tV��׌$l�Y�$��ߒ9Ap&�~yx��ѫzT�4԰ A`Ke75qeפ��=F���M�r4|�Ͱs�m>G{���GxL}��w>`w�W[F?�z)w!85� f�\�������7�G�|HW��XT���ؠ�$��+��K�6f����C���;	�&#e��͖-x��H�X��<�C�D�W��>W6Z,�	)߬��|��xO������Z��{�5?xq� �M��?����ɯWHP��� �Bgo�'���-��6�|t��V���h�"�c�?�uȖ��#I�9���>Iso�{a~�<�!����%Ѫn=��)�i\/��&_%l�,���@�9���m��РWԄ&mFɲ���*�$*�|7����P�Bc�"��,����O�)��@�;�0>���y�����_�~���T���R�����P<��RH�aogo��qĸ'����z����8��t�c,&*��v L��˙�eSƒJ���)���42��ȟqCa�ԣP ����������@
~9d�x���8+Ւ>�����M�"��������h���=$�d�������@q=���9D�A�c�1&��j��y�	������l�6�ʬS��u��˔
��|�����z���{Do�p��#-!��[h�XuE��7E�C&hK�[8����;f~�r��� Ꙉ&v�T�|�X� ��7G���a���$7}��V�P�7����S�w�Q-�����R�n& ��k�^?+�D�A�V�s> \0S�� *�ve'�+=�ղ�*>���m\���Ds��'��H�����S_f����>E�U�M��\9?��īڭS�:�RՀ�c8�^l.	���8e"�:��c:������^�A>�'���L�C��>�&̞�C[��.��7��e�����e68ݲ3�'���ޱBi��rss�	�`L)$�����y��Q�/�D*�v8��B��Y����`~�q1�ْ�2|	tEe��B��_��kc�SD��6E)ݬQ;˚�W��|�Vf��P�3�+�1��B��Q]%��W_�a#fP��}LF&�/!�S�A���N�[!�9���o㄁���{QM��*>Z�@��B.*�N�Fp�s�����Iq����#\~������}���C��3ƃpE)c�(����b�T�9�P�WL�&3�P�.�F.���%*7F �=��#��	v�^0k���u�DBҁY49�L�b^|X�C`Hl~�c�
>(���=�}���`��Ʃ��dF�}�M�"�nP@���[�c�X�����n�����Q	��R����L��3�ja����o4�!`�FJ�`�px��6������/�o���`S�¦a�;�f�$����C�-������۩��)�.*)�׃�l�w�t	m�؈`���^\� o��֘J���uv~�V��6}w��%ټlq�AGҕV:�St���N�F���1������3��]ҕ
�bD̥�}��z�:^s�o�1��*�H{_� �e���b�#	��X�)|賿�-8sAK��� �������Y����ۘ��5m���P���r��&���}�P:o�C�������03-�ځE}�P�δ�	�����.&����B5ۛ/7Fl9.�o3���mbJB>Ɖ�L~N>���ay�E�7/^�Xm~.>y!Z�}��{݁�u)�j;%�m'�<�r!_�UN�B� ��k�]T���&�>���P{0������l����Eq=�!7�ԟv��r�v8�]��$�,����9�?�{�E:�:/q.j:d�Sz�"%�������\���o�ݫqt����n��ȟo��c9�lCNj,�\��B��WD�g���i�O���2�G1��a�hts��3L�R��U�pP�]�5��㰎|�^g\��M����h�m��\�D�m��{�X�Y� �Rk"�Ș�zI�6b/�IUe�n��l|V�I�����C:gk<���+fgT	�<.������<��Z_,9�G��U��'Ri�钹ь{�@�,C�ޮI�O�^�@���y�/�[�:`�+�*��2�F�k�s��ـa0�Ż[���Ƈ�� ���{�[�:��/�����|boV�<Ң�8�n{J~��b �ѨD0��o۽���ƻZ������axj�=��7B��b��R�4�3f��� 8��֣G�ld�N|
����ᅬ=Rb���F�вȠh�Id��ea�C߮�r��/��́��	��2@?�ȏ�e;A-)���OPrP������%܌ya`6P`�"��-R}Y�����2��S��YL�z�Q&�ָ7��x���Ę˗��h�ʘ�ek��.��~"�R��8�T�&ES��7��Q*�@\F��%�a�C��c��.����n���I[��!�����y��L��0��
�ia������b��[���:�Z�_$&d%,��h�+�hVk��8'�i"'V}n���!g�|+Y�`��b(����|18�Rw�ԙ�ݶ�۽�tD�I&���HZ�ϱ��A�^R�ω`-�ni�S��5o]��>m\,1,�3�~���s�Jl��
�;����	��(�*EJn��4���f9F�ݤ����8�w�:��#��n.�"���c�S߆�)�-w��{j��N|E��{�̡�S.��Y*�����O����I|Ї.���WD�N����Ɇ�0E�@+���$r��Jp�׶��u�x �p��
��+rR9�)F�s�Dr8�㾃��)��w#�k�oM&r��ş�P��nю:����*o���zl�o��	��e�ڄ�*�>`ZV��sȒI�;e�YW���A��*�/�G	�Ҩ5V���[B|���R�.�CVf.�{���yݡ�v
�y��%b^�J�?���&lԗ�q����W���G݉�Gǒxk�_�&�w�\�c������i�r�y���;ɷ擋�;uhv�t_�#e���f(�H܏u�IKچ�D�ۓzV|k9{!��*�=]h/U�OQ��@s���e����p�T��-�:��B�|H�N���4KU`��*=��n�5�~	�0Ѧ��*�?�ž��j��!�`����̚0�&
W�pW��"���t�#CS�T�P�$=O�[} f�f�� �عi�
����)F��*����cd�?���*��_�k|�:�mX��}5+=]Nu��o�M�TչtsA����=�**2���»-H"��{�Dyh�v���ݛ3r�>2�Q�
�&�Hp�oÁ�H�,x�U��`_�&���ƛ˔������X�A�M�0�;d��J��;�ۧ�n1������#+����+���(��4w�M���0?�IggVC����]�b��T�5�.��N��!�<r�ضJ6�O�zs6���f@z�z�E�Ț��V�9�x�2 �T�b��$�$`ۭ�BQ�t#�y����t@���E٨_)ԙF/FTع�����N^�3��L
1�aD l�����~K���Q9[�S:�>�Z�,I�>Ry��%�X�؀4͖�o��|��nm�7�<N�j�x��	��y�H�0o�[2B��en��5Z�bћu�{ 0�Db��Q����q A��[M�G{d��T� f)�,4l�ܐ��H�.��TBc1"�5�3jĬ�M��M�ÎI�షn��q��F����Z&6��{�ȼ��+�A�S��`=�sH^���*xl؟��L'#�_���"��[vgI��v�vv���S>��gIi@5;�.���\�2�2�Y�6K��.�Mh������'N����MM�-�b(uɊc�	��tK�[x�Ze.��ҷnj��m�h\�-�Qt�T7��#/>�mf�����r~3TmЋz����ұ�Qf���-YUy���L�x����a�C�5P���-@;
����)SI =���əD�Z۬�K��ܩq�nU�S?W�5`�1�� 7��^���ml��wt��5�^R��WτL�1�Ĉ~���+�X�2NF��V�=O�uE%�]{!-����YW�oU/�N��#�a��tD��Tg]R����C���}Z��lR���q�_��]���w�Mz�'h���q"?�d���4 `R��=��E�wiJ�J�~9��<��:.��\��2�F�\�úx�f�=���CvԹQ��6ȗ���1��L;-��a�*��b׶�F�ܒP��Oq�B��F�t�'�{V��dq�Pj�
9��������f��y��n�)��`n�3ʻ�H�*��P:Z�Kuu�Q����� |�p��JZ���T�d_U�tAju��ޗ���2��<�=ƳϨ8h�5�fʌ���l5�W��"_ʮ.���!�y�n���o;�]`��q��8�_��s�lQ�I!�*}�i�?�?
��X!�I��{z�G���)
�o��҃'�a"B��d(₮�a����AE��yJ��-��R���QV��(��F� fv"���[ڮ��w�t�Lsyڳ,k�4�g�CPl�<�s� �I\5�J��f͊�A�w}�bZ��M]vrU�z��]�l�����P_�|�i��Y(�n��(�Eש���+m+��!��]s��P��ve�nݜhe��%�I��͢2�`���-�OO?�KQ�JH0�pj��v'ڮ�Q�^x�hl�Z4��,�P�ʴz�
~���)�B�Ɲ 4�/^��0�;��f[�C�&��R��L1l��l�|����f;##)��x��5!��:�R�tlO􈧩&�D?^)��^S&��n593
MLC�w�G~)�F��9\�h���0��l�x ���7��h��BT��0g�]���;��+�e`>���񚂀3n��i�>��`#���YҼLd��e����Φ��Iځ�l��Q��& �?]��Ϡ�z̦�F��ԉ�l8�o���u&jq{B�h�&�6Ȕ��>ޘ9��E�����l�i����� ��	u|��������?tj(��Φ4��N!����X���x�
>�w��k�����Z+F[V����
�h��Y���"�wV]H��ۚ�g������C��iܑ���9�0jL��^ݥ�]�S��0��tуi�-8A�_^�z/OH�f��ap �lB�~l���z�Vd��쨇�H.���U&a{-ҋ���mh"W<z�(��Cg�J���&��c��Sb�4��Fz��6�i�q���Q@�7=L<�ŵ�>֝����QV����Gc��
X����K��K��ɟ�?�8!�.:����ߨ"�l�d��3�35a�s�@��h�CN��:c5�3�T{��=.��B�ԧn�>��������X_؇ ��/PU�bHZ�R�mv��$��,���у�i�֔>L=f6輎�/�8��qu���RAjE��>;SQ�h���]3+����`̻�}�����/S�Z�ID4�G��!��XF�pCq�R����::�"���	8p	:ն ���BJ��|6`M������`Z7�P
�{�hI�>Yԣ+��1�躕�Ǚ�H@ � �i��=)��}��F��O��ἝT����PK,���ױ�:�.A�Ƀ!Q�ư�ٟΕ%:(k��L�p/�i�l�\^?��|fa��b@8�aw���9��-ྗ+PNg^l٭�]E�px�	a8m���e��j�yF��L�ݢ��Gn�2?�z�TJ���[nd�������O|�QD�����ʷFʎ�S.��u#�-��ے�x��V����Q��r����Ge#ق�����U�ٛlO���/�MK�}����]���Н��)?J�����ܿ�`@e;&��!A5H���"�ζ�s�a�$�z9�K��LT�	�'���3�H�m�-�������@EZ~˦�l[����j��\��@��_TE�����)p��������C=N Myi�l�"p�����hT���>N.bM�H�c�i��>EZ<�����agJv/���uplG��5j~s�G�oB�r�7t�\���[T-��l�Tp9c\ٲ�e�l\8�x��=)Ż(��MO���ϳ����V�iVo�z��C @��ڢk��c[����26vg�&��<�p�X�V�)������]<��F����`�W�)n$��!|.b|DF�H6v�f�|���}�[/���U�m@�t�thDu��6܉O'u�����<)ə�>.�·����pjV��2c��vy�(|��?߳~j)B���G�S/��w��C�Q��M߸����+H��8�T�P]w@Tu�������L���w���տ���wW�gʺ�>�^���\��杌�.�~�XK��T���>��	�О�d���<f�l�.��r���L܂v�t���E㄄@�f$+����F�ѵ�����~q��4S�+���P�6���JO=��)���l��vΨ�=�⭝��Ì.��Hs�g�#2w���X2�D�cӶ;|t�z�Q8Ev�?L�N[_.��f�PAT@��ig�Y�D\مq�Ժ��ނ��Կ�^����uuԩ!�p��S��p'A	Զ�H�"��>۳��:������uw�Q8�U�W���C��˪�I!f�|�o�U��@v�G������i�}�����ȉ`:gzu���c��퐄L�+�	�������Б�Vv���/��y���K�n���6o�U�.�B1fi��s@����A���߬D-�NL4LS��&�kZx��@��`]������5'���X�o��BʝE#�s��4X���jEf>~͈�p�1����6��u����8a!aЃ)���b��G���މ���,��\�N�q��}��S�JΚ�Z�b�(��)�ْe)zȵ�k{�Krr !���G]Ko��j?�����#:Y��.���|�� ���5���`�{�KC|B�����h4���Ƹ���J��wv�1��C�Q���/0n��ዖ̡Rf��]@>�a�YSݶ�a�����h�":Ŗ��No]�}]��!�b��Ӡbf�{����z�8]�x����iz��H	���G��\i��V���$��/�?�R�y�?b�L�O~H�8M2�?d���d(�r�mE�e�ğC���6�Fd�'Ic��_�5��Ε���b��c{�F�S�l���d�����|�gG1�gȻ��8F�=,]�}��o�:����#wa�A�*�R�=����%#�p*R&L�UB��Q8B	�����X2^����/E5�}AD����7�Վץ�k��Ԫ�<�3r<#/VryDҪ�-���O�K�>4A��q��/lY�x�� ym_��YP�=9���&���ړWq kX8]�K1��s��﷪3�O�|'sE2��_^w ���T���pΫP�p�f	�� b��e��H*d`��v���u�H'�gHM�B����}��F��u�b�[�Tޮ��&��{�}�*�j�_��b�)�	4��G�i�{v�[9��ֲ�U�����T8��_�"C���:���k�CO*z�=�;�%���W���~D�S�S�NX�`b�u�H:`�n��d��	�H�A�y�j����I�&��)�����0����
�[��� ��k�Z�ݦg�TR�~��I���	�t: �����H^�-D���9�'�w/��ԉ\�g��})��S6��o� )e���?S�k�+il���ND�}��m��,��>f�.M�T�ZJ�!|@Ȧ�ͧ�b���c���ԁܗ~��(�2Br)0�L�����\h1�Kr�a�A+���fq&)ѷB~Rϕ�43��[�����$n����vN�=o�(q�?�%M����r�J�ٌ8�u%U�r����S7m
�3���MH�g�T+�خ�8�����������^���%���r�є��/�]^��F:�vչB�:������o��1ԙ*5*����
�U;ѧ��Ν@����OԮ�P��yN���S��J�`�`���@�yib)0	� �)�����@���{�L���1�/���rʅ~.
����F�7F7�6w�eoWV�;�ͯh������5��N��邾5�Ob\�ƹ^a?��4������b�i�0������_"������5�cG_��@�&�RiB'����M"h�*R�e�k5�9� ��3�R^q#���������S��	Y�y�j
��\�����d�(�&����dV���ѰcPdK�l�K�����.�p@�/�*-����~k|���|X�]����z�xY�r���f�k�ڬQX��<"��G����ţ��
B�l��b.�C0��j��%ّ�U�^Z!�Ar��BPC�o��zO��9,�S����[��=���Aq������Xn���&��Ж�0�;#1J���8K��s�R�dj��k[�H��t��X�~�y����2�M��1��#�T�h�,��_���`A�󑌀f{`*��
�Q�G���+0Ih)�Vo!=��$S�Y��Qp����$��z[��᭣׻���K�D����-���#4�bA&�I׬.G�Ȕ-��sW��oe���9�����|�SɎ8�Q�H����2�n*���̐�l%��jC�O����j5��<��<^�dgp�cp��
|�k�/+tE�ˆ��ia�oz�"�JWX����."Ϻ��9o�1��<����y�5I�L-�a���W���٭��khY6��!����<����;E��~{�G����jt�6�P��g��
��8�ߺ���~@�}�%%y�;4�aF^�c�����ܢ��9t��ȏ��4z���?��W\��{ݸk��H��=�w�#�vA%��?��?k��A�q�辅�N����yr,K�
̡O��ru'����9���P8B���w+���5N���C�������8�x�8��ҳ��4F���B;'5�oشy>�qb�ek���G���NI'Xr���DM�*��ڌpĨ����i�@9�x���ż�GvlOǷ�ߵ��':��3��`3��T��]��xǓ�g�]`;�تH�N^�y�7��,�R��:�V�兛5�0�^jL6��A���Vc �&�%�9���^���BV�>e3�����k�r��lz(�/<y-WK�g���I�b�)}����.p砆j�AxT��Q��b�<i"ޜ�}~����������<��*�8��*q0��^ֈ��mm��^�@�5+(	�@m4��L0W]���,n���S.x4���m>f��~�.m�5��2�Wȑ�<ooM�ƶ�;1O��o�K�R��<�M���4]��$ {�y	�����7ېf���(i>3��k�?�˄�{�{V-}2В�:��9���h�92���	�k�ත��y�P���C��<�''f��I�l�"�5����Q��w�
��0ӊ
Sx�+L���j���O%�F�	/V�蚦ڳ���l���W"d2d� ���y?O&sl1otWJ����٘W�~[�J����D��Ng\�p��Ip�j�+�l�0Q��X���iv��ufƕ�ƾ�1K�W�����e`�6�ym~��s�h#z�0�B�/q�x������r����澗.K���\�{҃|~�WZ�3��RC~�^�_�)��I���0{�L��	F�]0~�[I����Ǣ~p�NHs��g����臶��G�����ؽ�@I*�y��oյ}0��� �}W^�b��ZHY������=��ߴ�4��|
l�������m�O���^vo��{tB��;�s��?dy����X!}AS'(����1;�;y��~Z��8sn�/�l�7�3�c�.����U�8k�O¥��RS���	zK�LKSOs��yK��/��q7Ϧ�ݦ�0�v��Q��H���Mζ�/+�6td~�5��}�	�LABU`NS{�g$��\g�oC��'�J�&i��Ʀ�Y��d��˰�ш�Ay4}��c�S��~����yk�0�9.u�1���տ2�f��5ŭ&/e
��U(m��;�Du��֭A�S�at�\uoL�+�O``����W��i���zZ�CmC:��Xy"|WK.$��,uK�׭�j}��'��)����p�3��� e���Z�q��bn�Uk��X���:P��|C>��0�Q�cX��������K(��GF��p6In������B��1����Y��|���]���MNw��>�����������S�	^��8Y��^G4�b��t��d��^BL,(����@#'����N�g�"K���/�`�:�FLN�m�?	l���F�l&,T�����F���˱Uy��A�Qꗸ�o kg"����!h�����s��cV���^TR�ڇ��X��2�!\��N�$�P��~�v)�e�Z�4j�~� �˻?�D�X)[��X�Ѹ��\�Q�|?��>$�>]��S����,�{�'z�J�ϵ�> 2)J�>:ݦ���*�%f��S!�Bt��-_~v#�h�flGi�`1(o���FCu^���v�L���+�E��~D����B���5�d2m|[�y92�������Z��h�X���i�K,�����p����Ӯ�d��[�]�dZ��b=����ġ/�┺1�q?�V�o���%�;�]<Z�>�Շ�����f��Z9�Ɔ%㎠A*0��G��C0��>5�nb��/�A�I��[��y�8׳�n�.�%�����!^6��zl���}�W" �����t�X�8�o�°d�(�u�2uR+�{�.� '����퉓K�3�ΎC�b�d�I .]�>n�Y�(���S7|6�;*6��!;OܘP��BNu�^�Z�e�� �U�~Z�Kqu�ԣ<�Cg�t�6v3@˛�M:�ȹ۝����q����? �� H�"��ãjg����I|@��<@�<:������L�*��1�i}�- O��`�SdO�ްl�y�z#���=�!�͗����Z���b����A�K�䞚����S��Y�������ٚ�K�d	��yH�t�➺��o`k�>��ʡ�.%lm1?A_�U��`%ἇ �[�N�۲�G~vov�R�|s:w�>3��Z{�!UB��Ĵۏ=�2��b�!�J���X��N�9�����^^<���\1굝e�GW�L�WdX��fdHq��Y| ��;�LW�K����`���jD�%�n��ɓuҨ����p�m�m�GaɌ}��J<�M��{�U4��|����Ol�`�(���q�
p6˶
�AQ�:P� jF�x<2���������C��u!�dT�n���ĸ���Kuߖ�ĺ4h�Mu���[$Ч���#��Fu}r�!�¢[��oW��$)����}&���<�����pQ���l�э�կ��I-�"~�E��F2�C	t��R�m6+����%���$�3�'����fI �N�M<��a�l���	`�i���GM�@�3�Ⱦ.��e�%5M���6�u��r�-J��럥f�%��9܂�jm'I��C�`����^�h�M�+����4�@T���!k�����b��x©���s�W�TU�"�:��|�`;�-������6Ɵ�?#�i+�U"�iW��x1��.��12���@�<���ִ�w���F����ƗR�8�j��-�'�UsVmW������p�&�n���*�]�f����GC&6���N<L-*�˦o�%�/K�>�D��x��;�1bh	�@7�f�>�Ct6�mT�d��w1�{^1���8���ku� �"�jT��5���1		9������p�2k�2�����6�jm��qe����$V�g^�W�t�e�dA��ʢ2�K��ke�-a9�.��J~�Y��*}u�rU��#ه�vT{R��'�N���Q�R:(�e��ܪ`0��gZyP�v0��z������){�c4c�I��]�oN�U�X��LK�-!�mi�0<���I�^˓�u�����@��HGn�
�wL�1�CB֢l�l��Š��3���τ�u5�i�Cs�����0 ��X	��Ό���Y¢��V�K�G5�A�,gA�2�v=^D�LJe^lp��V�ƓjpgrSn��?��g����ȭ��*L����Ωx@o�����^0&�
I$��L�~qjפ(�@ȹ��=E���uݤu�0��W�Pfge���j�.�[��X�tG]D�d�����ŊrL���ɒ�@�\��S���ߗ�(���W����&��2^��{�e�1���Ś�8V!�j�����d���A'���.#d�@��吭C=k���0�^<IYlL��
��" �2}ܒ�$[ss�9��N�����~������2"����a�3��*x f6X2mG��
�^�Q$;[}xLT ���;U�f�EE�/1	D۹cl�N,ߗ{s+@��Q����R�Q�ӼH��96��r.7i��D��d�g�i��G�lP��i�~����	N��T���7�>ߪ�nʮw����n��$���Pd+C���)G���t���C�|�K�-�ꦾ�"{7&�M�ca8��9׺4�,��
���߬�~:�e�1��tI��Si���8%c��1k��O���?m�H�+Ϛ(�7�n^���O�I��u�k*��ӹ]c��~O⮚��jO�l����+ŝ�+M9'�*(0_nOu1@��h)G���!���L�vk�2���!F!���5,�i��H�a�UMaY14T���C9~�$�c�߱b�T�Ⱦ�X/��(v�Q���(��ì��r9�\�X��z������l�0�X��@H���n�� a\�J�R�o�@��ǦD��i�ڳ�����b+���f⦀�℧��>)��BI�o�^�<��A�y/��6�+� ��U&�}Log��:��
za��(��'��͉�1�]p�z�+�ώP
���� ���%7_���.�G<1�� �AsX._���=& �V�}_#��Ѽ��v�8zD�*�?�\̆��aцE�0$J��sлՎ�X�]	���M��ဣ��F�k�#J�G�2<�1�t}�g&��;(hOo�#���f>M"gu�N0���&Ij�RdX����q��X�AȘ���x~-z����'f��N���8�fE
��%eKソk�LC�ÈJ^��np���b1�K}�R�L{�z��A����-}�_*��l!
�p_tT���:IK>}���Wߛ��l<P��ѝ��m�\��hyjWm`�|n7&��xo�Ұ.6�aԿ���
�H]<W�|i��Uq�sF��t�[�dE�>{m��>[ߨ�k>1��9����v��2���X� �����F��/��W:֊t�rM�)p/��S�$DV��b�,tz����w`%����Y�7n�ۥ�u�܉vO��_�K�.�Y^�ڭ�T
�'�������	}Y�U4����,aE�M�%g�������u*����p5N�8L|�7�J#��E��Av Y��Z�4���$X�;���؉<����t��%b��ɪr��c@O�b��B�:aʔ}�(�br��Q�J���#����`�{2�X�c(����W���JpnY���,0���vSm��^gC��f ��A��RY���w���oؤ��4�_�t>�`�w�t���k�s ?ٸ���+B�'��
���w�D�j.R����@��w���I�c;H{�f�j�ݹ��ZB�(����[