��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf��4Oᐢ��\��QOVl7�_��s�q�I?�ϳ�������Q�����ffʣH��c�)?d���i ����\�O�W귓��C���Uk�@�EN�\v��T��N9�
�X����م�x"��XΫ��<qT��O2b�J��7Q��K�j���8g|�X`a��Y�v����eȍ��6��Q�d\bx)�[R3¼*ћB�L��P���4����zQ���� ������F���X��BNCk �Pb8r>8RX2�p$�p�u��FN���q��-N}�)hZ�D��>~<p�E��*5�5� H\
_,��e(1�cIm�`�$3!Y-���7��?��@��vJ1���o����])ȶܓ����S�h�X8c�Aw���ot��(��@�G0��u�Z��zL�>5�d�"5�e��Q ���� (�����Dh�X�P:V�3(��l�^9�	���!>�3��"VƁ����;|������̫-�ɍJf<�� ��[@{j�H
�DCp��-]˓����xĀ���ti�<2�e$�|:����Nb���[�~�vƀ�'�nqn^(�	#7�`��R�o@��qE!�����t��Ѫ�
��o�y��{��i� �#��s�\v���֛=��ڽ`
Y���v��)p��J�����ʷ��o)�Q��U�QZӷ�V�����,�G\f�PӶ%�6-B�zOb҄)<ӟ(��:t��j�w����*XUၬ�u��C�W�	g�QlQ����Et�(���)�� T9x��bZ�˵J��5R=�~Ѻ�,�y�pʧ�7	}�dsB�Jb�9�,4E|�Qc�'�ؚ��_ӌ?�}[k�����v��V��L�y�[��r�oI�(��P-:gZ�ki���������<+�H�0��`����F���^��=��
�!e��{���/	w}���S��92ܫl�q�x��M]���u��O�]T�j�"5̱�����L�u��x��"ZFx7��~Q�|�6J��<�����c���	[:�W��1qr�ꝍ�eg� ��NI�`������>`�]8��$"W2L����������,����X'�O���������,B'
զ/��L����@ClH--<�e�!h�%�z3[X=��$߷F�4k�z�1;Iq�3�%=ԷL�iJi��\���@�ϙ�q��h��w�5�ӛo����xj(�0W;�m��J�G@�d�f���\��=���%ş3���7;u����B�;)yE�2��&Y�#���F#-I�A<|;Ҫ�3�@:�oɂ3���--D�	K�2c���z0T0�I�����)���{�+�*"T�3H�F�^�	(����gN�}��y� X�b��4� %t����Dv`�K����|��L�0�����v�s\T?6���1�Z�1��s�+�-���$�������wD�ۓ�-	��H�-�|�O'd����H��\ʛ-��Y���]h��rn�KQh�U�s�f���e-{�]��Œ�M��AG��\��O����Y��`���#��Ӑ^l�*�������Kڻ�W3�YH�J��zs��P,J���1����9�.qU k���U �B��Øj'��ѿ6m��pO?�/�(��Q�v�u{a	'	���C�s��g__f�jS�O�崲9�@�Xl�Fz�$A#uY}u%�ޱG��e��� �Cʦx�CI�3kz:N�.͕l����'[��H�a����ʢȸ�M,%��[~9��#����#?-?�I;�0/grPZScu��>��
��-�ɳ��ݻۧ��-�`sUH�O=�� ��$�:��^b>��"����0�cPr�ɤ�ס�\A��\H��S�O��o�ʃ)�=ӎn��X*'���C����C�gFZ��f �~ﾷC# ��l�![ ?��^\ː��ު�я���D�w�����~��^}��vr�B����M*D�v��8�HH0�@�8���s\���>�|�8����?K�@��'5�l������������+�x-Ǘ=����B�����)����=�]"K`���\[l��J�H��H�P}�z:�q���ўWMfo���Ņ�5!�!wKy���hˆ#���H��I�q�t����� �"Jy3�k���~���@�:�'^�kϧ��^�l�E�bi&p�Jo)!l������?��*��P�~E0�n�~X+~�<���f��"��hd'�jc�'"�F)\��;+����E�e-�������*!{�ݏ
X'EN�zf��}�^�gW�l����d�-n(����4LX�}A��*�-�0 p���k�(d.m�۴O�p�ߝ{e귈SG��m������fK!��0�R��0XQls����R�Z�������*�	��&�����]Á��K�/�c#\��
��j���J��R��|"�m�b����d�N��5�i�K�\#���?��ϐŶ�q��2���P���)�S6��	��$՛��Z�_�A�<��^;�Y�ѳI-Y���NMs ���2e���H�,�������	p����'��
�8TA��P�/t��O�#�4����	�ٶjI��C�|.����\��Q��g����qR�q�%7!'�����YR5U���3��M�+�L?G�\I0љězo�q�^)n���c��gĹ̕D"�Ѯ�afX�������=zg�D-���i�1ʿ'�*�s��[�Id"�X��=a����z�|���QPajS�R	����.���{O�����]�jC�۟��.(���� �|-�#%3�agpOjF���Z�.��_���f5�7eXY@3yAZCg���)᪽��J>�㊮�"�%���y�(A�y4��lkY���83R⹯�D���3l=�������6TUz�t�OY<!�&��f��Ɯ U5�&1Yc�i���nk��Ɂ���	��<��R�t���kW�����Ҁꓘ8xU6��NC��,G��	U�|#�	L����K=���V\}�j%��x����k!��:��e>}��P"J�4��r��Ha��m���LY���>+M��:`�Ͳ��<��|�DG�f�;���8�D}>��lW���W%i
�q�V��X�.���ע��
�s𤻰^���/Z��f��mke�e�n�k����3]EL=���g���������}	
㝒; `�����¤yP�=-�n�]ڎƚ�9��٩H�O-�5hKv� J3n��n*�ُ�DmI�21/v�G&�K��hͷ�&�G|=���M�����iN�NK��ޯ_h��m7�5��6yH�o;eH�(�%�J6=���>*)�����V�L��>
�=�͆��F��j�UD�d��%�{`I,��zՒ����d���㎛(�A`?��l�l���)@�es?����߲>$�=G.�m8a�ֽ��	i�����SE�ߢ7�$Y���α�s���Đo�����;Rԃ��?����2-�C#��;jj���z�HbM$�;���Ջ�J��"���#ON�#�t��X�s�X�~��eM�k�Iˠ������Q��}����F�1�w��K���͊����O��'�F�BV���a���z1���Λ��</:��݂>e�G���eU`�S]VJs�I]�nZir=�R�&;����s[�"Ѩ��d��a+�m�k+۠ک��#!D5�㯨�	�A`jU��¨7�\sooS�t�n�-�xR�R�I)<ha�b�P~U�v����ti�@ٝXh�Kڋ����㇝��D�c�_����b�D(u[ඛ��dZ�i���<|<�	[�V��B��7��?ϙ$�p�5AÚ�)�@�����b�<ϐX�kH���}�[��b��}���&��c�.`
7ʋ&K��zʳP��Kb4�F"^���%ڠ�㶷�KF�Y���p�<LH3�@��g�����Q� �S٬�9�PK�Y��@��_,JG"|Q��K��42;�5	#��n!��n,Ӝ�	�~��;�6��d@�gA��y��٨�0��7SmAi<�6�����Kqex�&���ڦ3��b@���}wA�]�x�=�&Og'z��X��������� �7�M���/;��|7F]]�=w0-W��RZ�z��N#�&Jԡ�E1s��͓���TH�}��
&���ҙ{�{����zS{�2�ג��\gR�5������cӉ+��Y�1�Ԙ�$R�5\հ����C�,��,�����@S���1�����9NU{������[�\��n��a� �#a�1��#��ծ]���hx������O+L��nC��98�?��3���s���qs�*#��r�.�ְ6O�..��r���nbhG%�t�ز��#�a��TN	��S>�-� �fy��۰q@JJ�����W��I�,Z��J�������v�����bI��M.�:��BF�/��D��@%9I��t��"�����\@,Q�@�{��wI��7�ݢ{0���a��W�e�?�52�u�a�z��0�H�W^��(`r��T5N)]�������m�ژ�{oF�g֞oe/�����x�����R�-4J�cu��:�������$������R8Gc�g�$���"�`z��(,�ފP��I��@3 3����#+��] ֏�(�`��a�2쎬��Ͽ�^�Oֹk���D� ;{��o�{��݈D}�����zg�d[ԏӶ+���+?�+�[;����)��ɨ�yY�W �����d̼G�^o� ^�&��dSop�x��Iҕ\g��P���r�^k��7���eF���<���P\�w6�r
�u_
�xB��
���z�f��'��o��HQX���0��¯��1����E"z2��#�x�m
#Ǡb���<H��?Z𑫝�i�]�u5�Zf��I0��$��	K3��$�h��~S��� "w:������Q��４}���A,���D�dcr�c�yh�����qa�f�+�F���'@��3Yw�S��/��W|޳R|�@U:`7�#�����}\	r�i�L��TU�~+��d�Dk�t�L��T����A2����V0�J�RP��¼u�,�U�ӳ�Ǣz
��/�s+�M�,%�Fʶ��r
n�v�!3&���?�l���KX�Xзo���j	9#
E5S�m{mea?i�	I�[�^�`[��}�}����9�]��[�����EG �Ut�xT���Ho����*/ob�#K�m:�&�sO΂�D������E����BZ����4[Kx�6k���uT�SŶ�3������C(+ӵ��R��T���x'f��2S�/�,�D �qc`�	���u�~����?2k����j���ę6E :���T�Ը����'s!
�l�l��D��LF��%�<ݪ��3)��̙*�9��ɐB���]�4��F�2�-.7��*�oys"0��Gf
�5����h쵞C�Z��ٔV��v�,� u��+Q*�+z�m�K���OVj�{]
���xj�|�*�>��^D�P;,�%\j���{��}k
�b�o�����UN;�apV`�c�
���f�g�&:C'���}be34`j*��
�ͣwZ�7��}k��A�z]U�=<*0l|m�o�kH��/�����z�xvԻ��u�{DC-��0V���{>�
'u���o�E��t^�k���������3�����2-��zƫ�W;�!� �ʠc2�P9�膜�9(KT)�y4#����l����[��z��,�����q6Bi�~���v��+�&��۰���n��;r����$H:�����@%~�m�P�M�F�܀Q�����ïg�ɪW���s��o�k(�o�E�`�[ɧ���^���ft�R�Ü���Oq��=��\���O}{LWR>B����7�E�`��dX��hc��4�x�7g��VR��Jʳ�,*��y!ȭ�.%�X���}��d�{Y~Uz��0�˰��Sl���W��Z[i���bB��-�_𽚴���:��q�8��x"�V}א`�(T�f��L!�`�I&/�jt�}�8>�$	��a	U��.�}��UL-�d4ܮ*K�\�*�N:\DMJ`b�{�Z���d"㍩�KQp�S?p��ek�0ِ&�J�'퇫O4omz�)`
���� �M��R��&0���:����
R����o5��%k�����m�@zљ�z�/�P1-V̟��E�ab5�j��6�Ƞ�����n�D>pzo��s��'�kӍC`�f��
P�7v2�&�!�veb�/��r���?g1��ǖ9*i<����C���w�I!m6�G���w�7[�Ku��z�d�-�H$˃B�w^����j���f�-�p*͇Zp�p���WI�����q��J�^z��^�AN�WvW�	�����71����HR߲UW7c;br�k����Nad��Z,�#]����;W�f�a�"�*8�m<���h�c�+��@��M`��`p|���l�r:#�q�*!$����HwSn�S�{�)5ۮOFFǾJo�&�����%! ]��y��B4)�aF���eM��Fy/�2���h��La��1H�U�}<ɑ�����}Σ�j���!E����2:��89�ҖV������#���|l��ݡf�:Vo1�]��W �p,�q^���ʺ;߈�h�XJYZ����n��}�9�O�J�1�Uc��S�Y��H��=��z^��Z��*�N+``�n��yӂK�z�X�\!�	��觛J�F���4n����.X���"u����@�gvH���!.�2�m5��|��w9�ɛ���J�|���h�����P )�5Ă�.`�C6��n}dS����򀜠�#�.*�:(�P T_K���b_�����!e����e>!��ǁMl\�wѫ���؜��{i�ӻ?O�����u��h��=��H ��XȨ8R��-���ᑯv$���yW%2hj�ܙ�BΓ�z3�
O�Gc~X<���Ʒ3���z�qtL���8���:}s���{�������ǐ4W���Z	�i��r� �$䲪�׉Ɠ�y�L�5y�]Uǵ��f�����U�\��d�YM[�q1K'>]��4+lKI61�X�6h-�u�uϸw@��/����Ѝ��Bt����此�xjO�ɦw݇�uQQI'Fo����[8�8�X��g�W}����c�q�7��PI�A���ݷ*1v䲈�e?���r�mC��|A2���b�B[ ��)Z�8-�$7���r8��7�k��j)�4NH��بw�����4{��کUNKĢ1H�i[��>�}����`)P��$Jɀ��.ip,0!� �h���os��Mǽ��1�w ��j;K2�\U�}�׈P��,�z1-!=����/���1<v�i����fZ�	�@ �(W2;9�Gڋџ R�:$�e�9�O�=@��8��-����6�s�8�`8���)�kgX��E%=;z�Ӗ.ih�>(�ɷ��� �v%�x��<��A-�l��n�����{����4w�!��������6���a�ψ�f��$�z3�tO�S��|���R�Z��
������ZќA��Y������(�_�t�\/�s$Y���޺�R�`ͣ.�������i*k:����>f���[B�-�oR���/���_�мmey�i�	S1��><X8^Ϭ�r�Tګ�����Z�cP�F��|{����.���@��aw�
]�A����Q!�<8�YS�V�"eh���P��C�:���V�STަ���G�g���=�����0!yf&t�@n�e`Bh,r8��d�~<� �Ȅ�D��R����L�Ik�����TIm{_�LQ�?����Q���v��?BV��k	$�����z�R�#�>�r��%�w,���?��ڃ��l��=�}���o�Jo��q­k�t��t�����N��6�/Ns㹛.6����D���F[�"Ǆ�?�E�R�/��S�n������VR���-�F��A�����[��n���^��1_��\�����|}-�����2����� d�`�r��9e=�R�T(\cF5ҋCP��%ɚC��S�!�N���@��S]�q���r�t�����>�d�3J+�
މ��޸�UY,��/��N�d~��P�mk������=�3~9��ٞ�%�;G�����8���F��O��. � �:	����}�ti���;`��L�����:.��ʻM�!1�p�
=IZ^���� "�C�
��d&��A>$(�Cq���t�DV{HI� В�FR�WRoM*��gъ�ԭ^=eA���eI��\����h]4S�^�X�*wul�OtE-v�k2���雷޾_m��1�Cƙ�=B�>h�������{x�[��8%��q
��0+��حr�'ܺyr��z�,XNF�iF��F&8��{�-O������o iߞ�J�TT��*���z��a*�=�F�5�RSČ�쩰�?F�:!���y���~�ԍ�P�Q�zo�2י��Mj�!)����t@Ö��+�Ƽ�ҕ���iƏ�S���v�ñD2���4JE�	��$��a��fN2ѯ36��#�N��t洸I�;��J*I�G���}Ì@}����)v��wdY��'MA���j��ި�,iyaC���L�:�$j�=������� �^�\u������;�'a���#ړ�,�3y�Ɣ�) ��UP���h%,�	Ƭ������9��F��*���D��^Ƴܠ�ƥw��-�|�FRb��QA��@V�̚y�g�pA��(����_�e������KY2�'�j��q�,;��ɧ0��jѠ��@�O֗+tt��#Qka�#r+�gP��2�a�4����V���Oe�Dg�m��9����������	F�l��#�`��03�>�㔪����w�6^��F���=�K�с �n�����T R*	�'d�V��z `�}�~
�c�0�$	���k�J��c*��Qr�}}���$!�뙖���l0(�fq��gJ��9�k��QρP�}�J��p���H�a�Ӂs1�%�لZ��wK����؅��T�������"�-��b=�0�0%ODn��A	-�G����`�F��,��Qr���a0T__J�s1��\=�������8k��	P`w��K�'�t*_ɉ�p��zG��+��6�og���h͐o�W�>ªV-?"�o�~���6�&43�u�V#k6��,Ї!ݥ;,�P�F�
��S����)���VjyA�c��\r���Ue�3P��@�cEW��Őp�kvE���Uc5*$˔��(�7��¨�u�[!�R��[����ʞ���Y�r��g7A��8�����p��	�J��O��9��qFK���4+��Ɉ0t[?O3ݣ6&�T4E��2���.E��#���b��X\�Ui.cNoSF�xym�4���_��B�k���m�(Q���������D�?�w4h��j<���4�q�;�$>i�s�˃]���7���2�>e/����{�Z��){�1����u$�s�Q�Sg;��k�+�.��cjo��l���;�:mQ�;K�L)n�A�5;م�]s��Ѧk��f:*EH,�7U�~�XG3.L��~�O��_�j�Է$�&$�f�`� �F�؁|h2�h���_����w)|�_�ŉJD���.X}' +d���J��mG3�FN�aI��8�￈М�v����J=��Ϫq��9Eufe�"[��>7�C�����M,�ߝ��wM0�k�:����1d�3���ii����	;��t*��>�������U@�d����F�.T��׍[ͳ�B���}5<��	ѐ��'�P`�/�)�gU�����ზ(���P�6�75��Va�N/����S��}������ߧb��滊�M�=�զ@���l`�˗���o����>��׃��z���&%��Dl��{ġ�t�1���M�ꜽ,�>�;um��-�-��/�6h ��-;�Ы����x@�$�f}�/ W�S�uU��a�T 3Y� �bc��B�w���;�k����ݮ`��8|O�]�m�s�_=$���pT�[62����5O8F1�c�K���ѭ��-�[!I"\?k��]� �{����~Cg��)E�I�u, �swk���%I��Rͺ����e�4IdĖ�b�=�]T0�#��eJ���c�ۜTG�٣x9x�����Q�3��'s�`Sk�}�aU61��h��B�)��X^P9��-Ӷ�@?��H�դQX�mE\�o�3vW�r����� t(��*{�^����Ջ68�p'�!�l�����c�~Gx6��r�HP��s8-����!<����7g�)bJ�q����
Z�f�s�����'�]UW8������M�;��LΖ�H��[��k�>�"�ƤGDؼ�G�r�� {e���(�����v��p����!/=k2"�ӽ�D��&�"�6�L�N};�`5z�e6����<7J�w5Is6�����x������J�*N�b�EF0Z"�i�,�	_q�4�j:1�����W-�]����c�6���Y�\�l�]�5�O��\���{`�s��k���V=�9�XA�,f��"q�]	�ވ�@�u�������; ;�`膽]v5�'� n��~�u�>��΁�O��K�͋ɧ�$ld����i�]l��ρ�tD[��(r����%��	�7c ��m�A{��Y��J���i:(.y*eZ���%�*d��x�\nr��X�h�ӆ"d=f�x�瑶���Ұ>#�����?��pN�9j�rh�,�#	|���7�P�M�O��x����i	�,J�$8A�6,'g|�Ahl7�E��r�hQ�ڝ�Ύ������n{��X+^2qh�A�\i����+�c0-�D�
p���а{a�Z��ԜB���6@D�_Dp�V�%J$?�k� ��όJ�������!�8�Bw�h7mJ�M���K!��7U�!,�&��[�
�_�ܮ(�/*U��>e*�35�EY�/@��?��5�s$���U�
v�Dg.�7\��Dfh��a��oNK����*��3p����_���c�@�0'')́^�v���[.BvJtSVԊ��L@S
O�z�|m�}���ap�:z',S�{Mk�¶�ٟ����T]���95[��K8�I�-�yN�����v^�����eƧ��'v{���E��ܽ���7�)4�5"����|�#�_.����m��4U=��1�/�Xd��4����)�V�J�?1�V����ص���A��ډW��o�a&�1ޏ��1�;�!\O�v�O'sI��h�N|�j�쩗0�_tۆ�U,%���[%C�
�'�`C-�w�M�s��].(���JS+��)$C�0;�5�fÐ������	�᯶L�_�N��d�e�8���:>rġ7@#E��?�j��s��X�����cc�I�9O,�R�����ߖ�� �N�}4Ƙ����@��+�0uZ�J��`~8�$:8{�gq�(\�+�� d+��͐Gf��R�3)���:�E<x��s)��/;�ԣ���^�>BR=v<��`	\�T��n���I�ɚK|5g��h J y�PbJ�����C�Dȭ�Ovx�Qeb:��oޢ��LE"��\|ana���h������Nd�a�]��W��cI���٪����K�2V�' I����E�.��{��\�dUx�U�;j��f��P���ݔ&��a ���]; n+��;Dm[�<�$DRu�ye1�P~���z��d
vh	�z[%н3ҎL��>�m-��Tw� �]haK�U����@�tMK<?$<��0Y�&�sVw^���LB��k�b�{����)���+�$�*��}�^��U��q�C0`r�WoEI��:���'�C����%i�0\����kۅ<?ݵ�+Q�x���9�{�6p!ey��̒*�h��q,�%=�ol�����P%)����{6{���@�B]j���2<�ν �ђ�4�9�#m���W���K#[b�?�v��t<j���!�����^�<�-A�dٜ�$�u�>��Ee
]첢,oC
}���M�����
2�9:ߴ�ʨ/ǆ/sTm��K��[SF`����u�^v9�d��B����`� }�O6���z>im�<l_���'�����&7������c��!���ns���"*�O��g���}�5����Ű���=����r��/z.�[d�!M�Z0� GC��������JI�^�p�Z�K�����#�o0�@L�V��y���\��C��,9���V'[�~�}���Q��O6zq��'}��j�CnՏ��v@=�����N������F���v��e���~}
3F�������E	̒��>(p��ݎ9QC�&�%AW^gY~�߹U4"�d>�y4���V>��)5yl����B	�LH��[RT�M����yJ�Q/�\r�#ea�ĚՍ�2��j�BX��m)6`f1�:x�uVl����|�_\�3�����=.+^ܸ�"�_#a������Ml�Ԅ�Z��g+dc����rVD�h��L���>����v�ק���r�s2�c�������xI�������{L,���asݎ�
]�7�»Le�0{N�����7�ld����`4O<L|v���d��_g������^�P\{_�$��q�	��Ӱ�du��D�,qi/��� ���҆2VK�r�ue��[B�ط"7��At��(�*��j
.�S�#L��{e��]��ݞ��fOR;���:��dL�����'�ug�z,�bF���X�̯e���`�!j�1�\Z�G��j"�,:�i��+�Vɲ��s��*�Ƨ���'�'��։"@�>н:�.�ܟ��LWʔ�!����&Ly�/P<36ߡG���+Cz�^��k�p@D	�D� "'�`��#��Bw��q怒	�_(�`82]�D��T�g����^|�/XG��bU/.$G��WY�BE~AD-/fP�9���ȉ/��)V՚n�T�"e�A���5[�%����Z�b#v��q5��4vu�f����ς��j�4c[�
�S��آ�k��,oi���szpS��8�1\y�Z�u���>Y>��G�U1Y�s���e�z�F�� F(��v��K��	4q�?ʦ���,�����	�Zf&����J��&�	>���珃^�F� ���-��W����Ƒi��By��Q�g'��k�J�u���%hb��c���B�	�.��_c�g�o�A��6GR|G�~Ǿ���'�,H���XV�Zۉ��N˹���KHZ?�0�`�/4�<������LE�^�m;w�l�k.�u�U�H\Ӟis�9�:�i����Y�Tw�K���󴚖m���?��Lu�P����<��<j:9��,����aA�0.���Ǟs,�N6""�y%�֖�ޢ�8J���5&bP��
/8���ɾ���.{��dŉ�S��2�E@��/=je��r��5����Pd����>�-}�]�w�;���ǲ���:qup��,bCQ�艥}o��#i�`�\�6?W�ܮ�τ�Ц6Sz�V�E)7��U�8�^�=�QƤ��2��T)�3�	 [ɐ��^쯪H��ؿ���
�R���H	�zyRܯZ2D��[y�muc���f�̙\�[c��o�h��%[(�=?x�������\�&�`�!U�/ߐ,�Ű�5���LF��0�+���E�kҫ�eǬ=2�1��ų ,K��2m�g:=�K�ڕ/+L37d��e��pj�֔�(U�>��MW4-��o�J��q�>���1F���D��^[E��]�	�l?I�Qߍ�V�uU�F'+N�F�Me�,PsI/+7c1ҬF<�7"���x�g��L[h�>2FP~��
4jTe��R�`���ƛ����;�����G�qU�� 4#���l�lm�vy�!Y�?�|�x�`;�9#Y-9�2Y~��s�>z��Ti�N�E�&p|aB��!_.�0���/�8l���dY'��id�f�Nw�����N�v+�j��v�|_�HC؄3�9��E�aU��G5ep����F���h���L_��%�4C�'�W&�e�'�T	��Fx�QG�����"�G��F׮d5�:ٵ*��l`e�N��+ϭ0%O>w�rw��9�')�U9φ��c����]�C�s<ys�{��߈��<pxC�hw7��
r��i��'8R65V��Ux�g�n��A�&���腘ҥ��աW�1��f�I[�Eq��î����)#
|��u�A �~�Ͽb�ޢ(�˹Cl�0�������.�� #���d��[�ğI��S�Kc	�|&4{r�;:���k֐�q�<b]:O�"�S�[6�
��F.�uG*H�Іu�v&��=('���䡦�������-,X�WR��pJ����)^c�!��xO(g��X����<3Pƪ��~��Ocz",�.E����PhJ:�Ql�?Yf�ͯ/~�W3�i��UʒL~ɨļ ���o��U=oTJ�<c��%d�DfOK�@d"��.����wW�����O��c��tz�1Q��?ʎ@�и�Vj���O'�;�;���x��>Ǎ�dR?(�qy������g);�С�H�:D� X�o��~¢�T�:{��b}�x{b�:��$�q-��,jҢ,����>���\=Q�����>���n�*q�}��=�b�N�t�[�s�D*�|J+�(Hj�
h��/�kc+ ��яP�O�a��"�xOPJf��V���:َ؂�=���s�_��B�F���6.-	�J��!y��y*��WxV�3��d�{=c�ϩVM{2;8T�qV��G�vc�j���G��X'�B� �v|փ�vp]I#��V�I+����#SF�z�qlq�,�����xz��׿-�B]_�㯙2�d��YX �#� � ��%����O�3dd��(H������`3f�*�6\c(�w#�x��h���I ⤻(�{�Cul=����f8�_�a�m^4t��D���K�����>l}[F(�[[$�����99�/��d�k����M��!=�����'����Z~�C50��ud��������Vq�V�/�L��)`6�$	$���_��J+q#rd��ěP&�jf8k@i���ή�C$ꁞ�.#�!(B"��q;i7��9L��.��S�.�I����`��k�SK��m���޿�ʣ���u��\�A2�ʇ�6&c�ǵP���k���PߖXIy��e���E ���Аs��W�QHMx�X�㓪�AAq/)���(p^�a���u�9ك�޽��,��ύ�,~���B
m�$4����]�`���xVn�fُ��W�b)�1ӊ(i@v}�5�Q�c2S�#z�}�\Q[	�!P�y"{������/�
"���Zo��j|�L����p
\�y $�r6�i�C��	�#���f��8�-2룛6=�ew4ѫ�J쳨�D���mi��=Kg����8~�	��k��quAɨ���aQ�D/P#��1�t#�+�.�I�ݕ9WEUt�����?UB-���N��h1���T�Ce�������P�tT��֏`��b[~?�Q[^h�a �7*Z��.����FtN�c��O���w̧�:�������&z�:z�{#h�@:s�S5}}^��F�e��5U�uz���R{
��re6@��HP6�g�GT�K���[cs�
���� =�� � SW8�$���jI��_�;���?Y ��<h�DVH� 9�b)���Tմy4��g�u���P�����*�-w����/D��_1�NM��mH�k����n~ߠis���V���,7��2`g��M� ��W�v�L�K?rm�=�\��M��rt��f�D�)"�<W��{��������K�I2&7 �������7)]�c)ßd���Ys�췬kV�S�Q��V*g'k��*�}����A��Y}#Z��9~|���Hf6�Z��|���w�=������:M�|��q�4�[\�*���qtA5(�[���yF}'X.&WPK+__/t�ʲs��L��:� ��O��5<ʓ��4W}�E� �ˠ�ϑ�w̲�V��c���!l*����Ll��	w�jcN���Tm��d�d���v�q���2ku9��ճ�4_#�����X�6�/��]u=�cXLv�0D���04	�\\�f#�˛39-=���������w��I������n���bD%9���<q�����d��W}���(�}��Ho�}��l�m�'Ô����U^�r	�����׳���uM������s�pm��=iW������.�ȩA �_^B�W�q�	*>�4p�;/Z�o/"�i�9�A U|�����Mk-;MSi����a������T��k��wi�Н]uX�@�.���P�݌y��AMIW���5t	RC�����H�7{�C�Q&i}�����_��4��7("ڵ���O�&�N���a=y�'��X��C�A�-�9����1J�ɂ��]�둗�ғx��'kF��ȱ�u�+��qD�g�#�ȧ��?�'��V�J�-�t�Za��^��_",I,�-P��� ���	�}��ū@K��y�7&rR�qy㙰˵O�"�ǰI�3���I�!���N&�>P�2�0Q�����}t��x`d���N~�e�P@�}�?����̵�{Fh6��"�I����&�H^�u�E�%kH0����*����bQ�ۦ��S\A��"!։	�b):�Km���D�p�-#A`��K��Wn��J�.M�����	m�{�5��-��9gw9'���Hh �g��a��%wb�2�q(k��(��O�4��b�yP/��x�Hϛ����e?��V�@R���/�F0]��`������{����7 ��ܳ�j���