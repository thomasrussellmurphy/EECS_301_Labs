// megafunction wizard: %FIR Compiler II v13.1%
// GENERATION: XML
// bandpass.v

// Generated using ACDS version 13.1.1 166 at 2014.04.18.11:39:30

`timescale 1 ps / 1 ps
module bandpass (
		input  wire        clk,              //                     clk.clk
		input  wire        reset_n,          //                     rst.reset_n
		input  wire [11:0] ast_sink_data,    //   avalon_streaming_sink.data
		input  wire        ast_sink_valid,   //                        .valid
		input  wire [1:0]  ast_sink_error,   //                        .error
		output wire [23:0] ast_source_data,  // avalon_streaming_source.data
		output wire        ast_source_valid, //                        .valid
		output wire [1:0]  ast_source_error  //                        .error
	);

	bandpass_0002 bandpass_inst (
		.clk              (clk),              //                     clk.clk
		.reset_n          (reset_n),          //                     rst.reset_n
		.ast_sink_data    (ast_sink_data),    //   avalon_streaming_sink.data
		.ast_sink_valid   (ast_sink_valid),   //                        .valid
		.ast_sink_error   (ast_sink_error),   //                        .error
		.ast_source_data  (ast_source_data),  // avalon_streaming_source.data
		.ast_source_valid (ast_source_valid), //                        .valid
		.ast_source_error (ast_source_error)  //                        .error
	);

endmodule
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2014 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="altera_fir_compiler_ii" version="13.1" >
// Retrieval info: 	<generic name="deviceFamily" value="Cyclone III" />
// Retrieval info: 	<generic name="filterType" value="Single Rate" />
// Retrieval info: 	<generic name="interpFactor" value="1" />
// Retrieval info: 	<generic name="decimFactor" value="1" />
// Retrieval info: 	<generic name="L_bandsFilter" value="All taps" />
// Retrieval info: 	<generic name="clockRate" value="20" />
// Retrieval info: 	<generic name="clockSlack" value="0" />
// Retrieval info: 	<generic name="speedGrade" value="Medium" />
// Retrieval info: 	<generic name="coeffReload" value="false" />
// Retrieval info: 	<generic name="baseAddress" value="0" />
// Retrieval info: 	<generic name="readWriteMode" value="Read/Write" />
// Retrieval info: 	<generic name="backPressure" value="false" />
// Retrieval info: 	<generic name="symmetryMode" value="Non Symmetry" />
// Retrieval info: 	<generic name="delayRAMBlockThreshold" value="20" />
// Retrieval info: 	<generic name="dualMemDistRAMThreshold" value="1280" />
// Retrieval info: 	<generic name="mRAMThreshold" value="1000000" />
// Retrieval info: 	<generic name="hardMultiplierThreshold" value="-1" />
// Retrieval info: 	<generic name="inputRate" value=".05" />
// Retrieval info: 	<generic name="inputChannelNum" value="1" />
// Retrieval info: 	<generic name="inputType" value="Signed Binary" />
// Retrieval info: 	<generic name="inputBitWidth" value="12" />
// Retrieval info: 	<generic name="inputFracBitWidth" value="0" />
// Retrieval info: 	<generic name="coeffSetRealValue" value="0.010203563724686556,0.012932756030581471,0.01512270704821752,0.012068446880155199,0.003213435218133443,-0.009332425643292215,-0.021305432522186026,-0.028075493490979247,-0.026904015056020802,-0.018467932378731518,-0.006711281658122525,0.00303340633084108,0.006770326514160918,0.003935988141761719,-0.0023589087671465653,-0.007154869053087672,-0.006535131179731438,5.722228328130816E-5,0.00943594651043356,0.016571088393085416,0.017673176350322166,0.012565585272318096,0.004926811471388852,1.1774704104413707E-4,0.0017842044969155876,0.009464328670584035,0.018567270470924425,0.02309719489042789,0.01939796679160803,0.008705625414294073,-0.0032745920106467025,-0.009704965648003959,-0.006984173007706431,0.0025990310743164856,0.011775136788602385,0.012537755725159869,0.001318046980699057,-0.018112527768242032,-0.03615682427373677,-0.04285950013607926,-0.03433605823292291,-0.016238486474526796,-0.0016361231295620945,-0.003843469911322044,-0.027853422758449417,-0.06529532175930496,-0.09643614482306025,-0.09904895527969378,-0.060062052609500566,0.015982320586741032,0.10654735047658259,0.17964623721832346,0.20763643437223353,0.17964623721832346,0.10654735047658259,0.015982320586741032,-0.060062052609500566,-0.09904895527969378,-0.09643614482306025,-0.06529532175930496,-0.027853422758449417,-0.003843469911322044,-0.0016361231295620945,-0.016238486474526796,-0.03433605823292291,-0.04285950013607926,-0.03615682427373677,-0.018112527768242032,0.001318046980699057,0.012537755725159869,0.011775136788602385,0.0025990310743164856,-0.006984173007706431,-0.009704965648003959,-0.0032745920106467025,0.008705625414294073,0.01939796679160803,0.02309719489042789,0.018567270470924425,0.009464328670584035,0.0017842044969155876,1.1774704104413707E-4,0.004926811471388852,0.012565585272318096,0.017673176350322166,0.016571088393085416,0.00943594651043356,5.722228328130816E-5,-0.006535131179731438,-0.007154869053087672,-0.0023589087671465653,0.003935988141761719,0.006770326514160918,0.00303340633084108,-0.006711281658122525,-0.018467932378731518,-0.026904015056020802,-0.028075493490979247,-0.021305432522186026,-0.009332425643292215,0.003213435218133443,0.012068446880155199,0.01512270704821752,0.012932756030581471,0.010203563724686556" />
// Retrieval info: 	<generic name="coeffType" value="Signed Binary" />
// Retrieval info: 	<generic name="coeffScaling" value="Auto" />
// Retrieval info: 	<generic name="coeffBitWidth" value="12" />
// Retrieval info: 	<generic name="coeffFracBitWidth" value="0" />
// Retrieval info: 	<generic name="outType" value="Signed Binary" />
// Retrieval info: 	<generic name="outMSBRound" value="Saturating" />
// Retrieval info: 	<generic name="outMsbBitRem" value="7" />
// Retrieval info: 	<generic name="outLSBRound" value="Truncation" />
// Retrieval info: 	<generic name="outLsbBitRem" value="0" />
// Retrieval info: 	<generic name="resoureEstimation" value="1000,1200,10" />
// Retrieval info: 	<generic name="bankCount" value="1" />
// Retrieval info: 	<generic name="bankDisplay" value="0" />
// Retrieval info: </instance>
// IPFS_FILES : bandpass.vo
// RELATED_FILES: bandpass.v, altera_avalon_sc_fifo.v, auk_dspip_math_pkg_hpfir.vhd, auk_dspip_lib_pkg_hpfir.vhd, auk_dspip_avalon_streaming_controller_hpfir.vhd, auk_dspip_avalon_streaming_sink_hpfir.vhd, auk_dspip_avalon_streaming_source_hpfir.vhd, auk_dspip_roundsat_hpfir.vhd, dspba_library_package.vhd, dspba_library.vhd, bandpass_0002_rtl.vhd, bandpass_0002_ast.vhd, bandpass_0002.vhd
