��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\���V�fnvx��ÍG_;�ȅe�~�>���9�>��Y;�0G+��{���Bɇ���k�)q�Ջb\ǜA מRĳ�x���YoP�n����΋И7/�D�8 ���<�u3�����bz�k�j5�7�a�2aGY2����*�ˎ ���o#<$X�u��!ԉl��������^�2�k��Nm���V[K��Nbkr�&Q���x�G����+]3$����*|I{d���bY� 媋,��SJ��$�I��3lkk�}
i�������Ǹz�$�;UF��v�q|��x��H���m�}e;@��9�:l�7u���B�ͩ���zZ�~��{�^DY�'��i���͞�I &T���Vy�b�{�ڰ�Cn!�(�"���sf���K]S���8PǛ�}�vQͻT���``��9ع[��MŜ���'�J$>�%���a_�����re/��֖W�y������{�P^`"��M��ɥ8QdL%��;����m���Mg4����`�!D!m��ެ6�'�d�]*�K������_�� ���`� ��	���､�me��q�H�H��;��.1��i�;�}u�rn/�9V[��$����Mfm�^)q3	0�^�L��'�W*���Ɛ�(Z��c�?�*C˱�2��eiF.�x�^�܉�S�1�w��4��"1����z�E	o��p�e�!	�i�Oًg����\-{ń�Ԣ�������W�W<9(s�o��^2�sӣ����6�`��y�iO#
B���7(ky5�bU�fm�6*�>-1�u��b��8My���hj ����tp�F5�������q7���Nu]��,�niK���Y\����2P����c/ܨ�W�Z����	���4��{�8fj���iT�1�';���c�j�C�*���E�;��9�5���8"�z����~�^w��ݳ�.�DD��̗:���r\v�֡sZX�gb86ǀ��y��}�M��\��W��/Ob�"�5_�G�=c�e�D����H_��U�+(��xa���:�˼_�1��4\uM	����T�e�:%�Sd!��I�@N
���}X���h�B�<��>@�X �4$M�j�B>�q�$1ޏJ�����s��G!ܫK��--�?��8"?�Ԯ��Ñ5��x��5�:m�h��]1�,V�h��N�4_w�y6	�N��,�*���֝���3���b�r6���kB\�b�D��;g�P��_�b�nE�::�@��ƃVfg�&`�Mʱ,m���}���nl�� ��>Ԟ�8��z��-�"��N�[R3%�OI��9ؗ�Ƀ�mj��7�4�3�:����S1�Xw�
B]�$L�b��oH��E��ZY�h�	���y	&�����x �P�p���*�{�QoR�-��(hOi��/� nD�)}'u�O�%I r����B���̏��;���q�J���K��~��6z�ڝ�&�J��0��e����N��D��.�_1�jD
f�k��H)␚�>
��'X��)��t�#>1