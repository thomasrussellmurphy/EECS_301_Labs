// megafunction wizard: %FIR Compiler II v13.1%
// GENERATION: XML
// highpass.v

// Generated using ACDS version 13.1.1 166 at 2014.04.18.14:44:35

`timescale 1 ps / 1 ps
module highpass (
		input  wire        clk,              //                     clk.clk
		input  wire        reset_n,          //                     rst.reset_n
		input  wire [11:0] ast_sink_data,    //   avalon_streaming_sink.data
		input  wire        ast_sink_valid,   //                        .valid
		input  wire [1:0]  ast_sink_error,   //                        .error
		output wire [11:0] ast_source_data,  // avalon_streaming_source.data
		output wire        ast_source_valid, //                        .valid
		output wire [1:0]  ast_source_error  //                        .error
	);

	highpass_0002 highpass_inst (
		.clk              (clk),              //                     clk.clk
		.reset_n          (reset_n),          //                     rst.reset_n
		.ast_sink_data    (ast_sink_data),    //   avalon_streaming_sink.data
		.ast_sink_valid   (ast_sink_valid),   //                        .valid
		.ast_sink_error   (ast_sink_error),   //                        .error
		.ast_source_data  (ast_source_data),  // avalon_streaming_source.data
		.ast_source_valid (ast_source_valid), //                        .valid
		.ast_source_error (ast_source_error)  //                        .error
	);

endmodule
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2014 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="altera_fir_compiler_ii" version="13.1" >
// Retrieval info: 	<generic name="deviceFamily" value="Cyclone III" />
// Retrieval info: 	<generic name="filterType" value="Single Rate" />
// Retrieval info: 	<generic name="interpFactor" value="1" />
// Retrieval info: 	<generic name="decimFactor" value="1" />
// Retrieval info: 	<generic name="L_bandsFilter" value="All taps" />
// Retrieval info: 	<generic name="clockRate" value="20" />
// Retrieval info: 	<generic name="clockSlack" value="0" />
// Retrieval info: 	<generic name="speedGrade" value="Medium" />
// Retrieval info: 	<generic name="coeffReload" value="false" />
// Retrieval info: 	<generic name="baseAddress" value="0" />
// Retrieval info: 	<generic name="readWriteMode" value="Read/Write" />
// Retrieval info: 	<generic name="backPressure" value="false" />
// Retrieval info: 	<generic name="symmetryMode" value="Non Symmetry" />
// Retrieval info: 	<generic name="delayRAMBlockThreshold" value="20" />
// Retrieval info: 	<generic name="dualMemDistRAMThreshold" value="1280" />
// Retrieval info: 	<generic name="mRAMThreshold" value="1000000" />
// Retrieval info: 	<generic name="hardMultiplierThreshold" value="-1" />
// Retrieval info: 	<generic name="inputRate" value="0.05" />
// Retrieval info: 	<generic name="inputChannelNum" value="1" />
// Retrieval info: 	<generic name="inputType" value="Signed Binary" />
// Retrieval info: 	<generic name="inputBitWidth" value="12" />
// Retrieval info: 	<generic name="inputFracBitWidth" value="0" />
// Retrieval info: 	<generic name="coeffSetRealValue" value="-0.0053835052795455475,0.017457594967310367,0.0017682548052020955,-0.002746624734616668,-0.0039803354564860284,-0.00425329886609632,-0.004181204887671317,-0.003872261192041397,-0.003304498064728045,-0.0024399982725885,-0.0012860823219235612,1.0586232607250154E-4,0.0016363610327956022,0.0031571959051302505,0.004496485230871312,0.005477931663470896,0.00593614294035735,0.005750192684917203,0.004861474113543832,0.003277125622238054,0.0011012299658650494,-0.0014846593361374611,-0.004222236843786738,-0.006822786236491282,-0.008929134580193546,-0.01028762215466291,-0.010556384427359953,-0.00964452310263456,-0.007441753249432458,-0.004030444150626832,3.342324056203246E-4,0.005316823654384976,0.010440697069758044,0.01511301541699726,0.018747233570988373,0.02077062004486329,0.02065805759302448,0.018019127788853746,0.012647298028070521,0.004538224771975385,-0.006100723844520582,-0.018855627407234236,-0.033103853346400605,-0.048045978870335834,-0.06280729185346626,-0.07647962604955479,-0.08818521422642893,-0.0971552041577995,-0.10279919383146127,0.8952874797309053,-0.10279919383146127,-0.0971552041577995,-0.08818521422642893,-0.07647962604955479,-0.06280729185346626,-0.048045978870335834,-0.033103853346400605,-0.018855627407234236,-0.006100723844520582,0.004538224771975385,0.012647298028070521,0.018019127788853746,0.02065805759302448,0.02077062004486329,0.018747233570988373,0.01511301541699726,0.010440697069758044,0.005316823654384976,3.342324056203246E-4,-0.004030444150626832,-0.007441753249432458,-0.00964452310263456,-0.010556384427359953,-0.01028762215466291,-0.008929134580193546,-0.006822786236491282,-0.004222236843786738,-0.0014846593361374611,0.0011012299658650494,0.003277125622238054,0.004861474113543832,0.005750192684917203,0.00593614294035735,0.005477931663470896,0.004496485230871312,0.0031571959051302505,0.0016363610327956022,1.0586232607250154E-4,-0.0012860823219235612,-0.0024399982725885,-0.003304498064728045,-0.003872261192041397,-0.004181204887671317,-0.00425329886609632,-0.0039803354564860284,-0.002746624734616668,0.0017682548052020955,0.017457594967310367,-0.0053835052795455475" />
// Retrieval info: 	<generic name="coeffType" value="Signed Binary" />
// Retrieval info: 	<generic name="coeffScaling" value="Auto" />
// Retrieval info: 	<generic name="coeffBitWidth" value="12" />
// Retrieval info: 	<generic name="coeffFracBitWidth" value="0" />
// Retrieval info: 	<generic name="outType" value="Signed Binary" />
// Retrieval info: 	<generic name="outMSBRound" value="Saturating" />
// Retrieval info: 	<generic name="outMsbBitRem" value="10" />
// Retrieval info: 	<generic name="outLSBRound" value="Truncation" />
// Retrieval info: 	<generic name="outLsbBitRem" value="9" />
// Retrieval info: 	<generic name="resoureEstimation" value="1000,1200,10" />
// Retrieval info: 	<generic name="bankCount" value="1" />
// Retrieval info: 	<generic name="bankDisplay" value="0" />
// Retrieval info: </instance>
// IPFS_FILES : highpass.vo
// RELATED_FILES: highpass.v, altera_avalon_sc_fifo.v, auk_dspip_math_pkg_hpfir.vhd, auk_dspip_lib_pkg_hpfir.vhd, auk_dspip_avalon_streaming_controller_hpfir.vhd, auk_dspip_avalon_streaming_sink_hpfir.vhd, auk_dspip_avalon_streaming_source_hpfir.vhd, auk_dspip_roundsat_hpfir.vhd, dspba_library_package.vhd, dspba_library.vhd, highpass_0002_rtl.vhd, highpass_0002_ast.vhd, highpass_0002.vhd
