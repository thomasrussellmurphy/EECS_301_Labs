��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�uwC�5�b ��ϴ�	+�
Ct� "�J~���z����<
�����'k�z��ߵ,d�.��Z�Ӝ��2�x$ҟdL��h��ʔf��#
����;�;m�ȋ��[F��E� &'{=u�3jg�b�)��LA�u/5{<	����[�Dn����à�@��cO��IEo�y~�E���ސ�m��X�i[�6����؛�sP�C ��������?����<��$�2\���sj��܀�e'�\�;l��<�&�| 
��]-1�g�u�@�ifW���%�zhK�N�?�
|��9���'��#��h��o�j/)b;fi�g�����Ac�x��o��������L��N�t��(Rw8C�Ħ��!#�%|E��i�]k�PإI4h����a����9�� 28��+�e�q�_mN��o�?��� 苊��+��̵M.�z��1r�-���H`@�wEf�r��'nz��]
�%��Ȼ�{P[��7M�������n����ނ\|~�o[����S�^[�8'U��C������벪[za67"Y�Y���J�ol?ɨ��.�Y�����^�*z��}5/7#tE~��|���z�L�}� �ܐj�YY�#h��7?}^׈H43�] ���L��W�<����:U��l�;U�ԛ�����R�G�F��YPD:,!dUJB��pZ��*	/�9�\�|�o�ۦ�Ĩ%�֯I��}ם�O�째I6>-����_�!4�^ �h&��B��� :���8DU����r=mӋ'��	)?����,I=��?;�l����m?sҕ��K�h�"�0^t��M�K��m������H��	µdZ��aβ�w\x6mM��SH�'MŜ��A�uR<���/�왎�@,�x"g�e���Ք������_�f��} ���Lō�����J����^���~l1y�˚� ��Y'L���~���VO�^�>�H�F�h	1����O��_
�U�}��&ᾞ���D���JcP#����Qw(K꾐~�O1�-!�.}�D.�T�8��7<����l���[N䘵L������a�)���I�W 7��0�^  F)i?�]{I/�!l�͐�j����vk����R�Al�~Ǟ>������H�3L�Vw�
��,����/<W���<	!��Ͱ]
��9�v%���D��LŅ����52�_��s�+	H�I�Q���ė�1�C��jN5��op
c�������@�;+���]��n����uPqM~�#��G}�h�V{ q��H�6���)��&Ly�)�;��Q/��aޠ��S[C��Am�vY�%�(q��~�����k��(�Ƕ�tl!�*s��woŐ�w
B��1�l�q;p[$�����3b⯢m�ӛ�D�7C��<5U�����۰�����S_�L��,�ަ���{)����󭳐[���`�A=�;s4UW����
�@_�/%�"��������"�&4�l���/��H�x>��T���H��Jk���&��9)�cwW֭�n��J T�ƒ��.���ӿU(B��6�aU�%�ؒ�$�Ӑݜ�`�T8�(N[�j���>�y����P:�f� p�>bg�˷��r�;p�?\�¡x�q�ZA�8YuBY�SѸ	��e��}:��Ԃ��������>�z ~�����#N�2��t�	�"�Wu_��}�ǡ�� ޼�����i��Q�^x0�*�D��YN��<S9�=T�ɣ��Mb�/8'���-�W~���8�/��Ҟ��z�����kڽ�<a(Ȼ�]v��S
�v�u9��Tm)Yr0Lۚ�@^�Nx��q9Q��hם\�O[&�;U���&�.b��gAA�P��Y��P 1�Ft�]�'g�l��Ga�k���;��Cy�߇_n�ʢ��R������d7�aȊ��!\���^�2��)��1�P��
N�?Х��� 	�57� 2o&k ��v��u0�G��`v�H0c�cW\��_��J�ҙ�nJ�V�Lზ�ŗ��(���Y��62W��:�Ή��A-�u�"Qti2+4\��z������=8������A��lJ}��)����u����B9�up�,��7Z�*ܾ�Q�N����@�U���Cq]�����Pܸi�m�)� +�@�;6b�~�L�A̚0'��o'�V|�������	���z4�g�����3*�tv�Z0�����P���Rb=O����le؝Ȫ��'B 0u���c�4��l/^%������Q�#�q@�l������d��d(�C��2/���U	q1Dno�n��8yN����{n�_��Ƹ-d�V�l�uI��,E��pݎ��ϝRq����*
gh$?�{T�:��إ[ſ�F4��=�
*������ʖ��zI� D��f*{Z�g��A	�P��wFg뙪�ިu��:y�D5�ǾA#�Y���>��I@��p)kգ�JT7SL7�E&�rzwoF�O�7^�UU�N��q�>�E.��"}���ʋ��ӀP�h�1����G��@�Л�փ�*�+�F�2��C�'�J&�`4��oB��]��n��񇕆9Y��@���`,�c���[�Sm����TrAp��g,�n�EbEG_�.k��7�2��wl�����x���>_D��3ɴ�9Ӵ�c#U�j��b�6E|Ӷ-�������4'�*��Q��u���c+�F�_W`�������'I�I��R\;�;��������Yk ��8�J���ݥ��>���²����P�4g�l� 0Bn	qB$YH4�Kӯa�elH�GC�֨���NU�s���Z����Q���[�ȍ/���˕�?(�j��#m�@>H��ə����� �.���P�p�I}��?N<ҽ\�z/�����N���A�+��#�S���0�)\����}�5��j}ؾ����J�<�6O�T��*WU ���ۦUwտ;no����*��[#��f{�,��n��:���_�ظ����:q���Ⱒ�����������O�r��6�|Qeǂz"R�v4��]�����R����0C99]���5Ϩ�q�%>g��(PG�/�s�����#��Dj+�XǷu��b�N��7��RD�0����"a�К�!\T@�>G�:ߒqn�B����V�9�,[�_���m�@�*�\p��Q%%�
n�8���utJ�5T��[�F.���!���������IW�B��ڿ��$dD� m�S�n]ӆ�ܬ�0�K"f�#�:AˡB�bˡeOx/^�c\��h$o���԰��$������I��p����-������=�[%�'�5R
F�9?l{lX�0-s��qVъ��� �OL�`�/.�k@@�_�$h�OpU��w��qKl.�+Ѐ;�$o��z��3���*
��̺��ʥ+>d<?Bnșԅ&[#��(=c ��+����%q�!�Ϗ�.�91r��\N�t�aZ�me���rh���H��K�B�GJz~��Z��W2�#�w��Q�
�����~��=�~CIK/L�EV��K�5&U#���S�0W�A=���#���@����E�U�E����ǐ��03Zw���BDn�H+��A���-IHQ]��O����K�p�]���Ʈ�v��k�ר2�v�S�6̿�.!S{F�`��&��G�Q�uď��~þ	8���d��;�����s�Dv<.��1�EH(XwEX��ua�px_W*��gy�ހ�Y�/�ȋ e������L�-<Eͺ�����^�mt�J�*w<��  's��`�R*�5�s呝��!S;���G���Uvt��&�0���j"H�,�6�p���?X�LAM�,{��B$�U��x=PQh>�����b�z���7[/�"%�?�/�ff__��@C�? %�c��IY Ǎ��<%�"��z�^�`x0�ݝ$y{@�rR���5��䡔�w�O<% U���{);<��	�NŻ3ܡ�T�-�9�q��-���.�x�a�H�o	����FB-���2j��B�׍PnCϯ�жMA�����Y���$�r~=N!âuc@i�p��D\.���F|΋�� hӻ��"���K�"V�տ�W�A���>��w`�����Wv�}o�7a	�6,K	wשs���C몼��Z���R(�3Ȥ]"+ѵ	ia�.a����ߥTc�����_� ޓ�5�/��C��S^��U���y���lz��u�#�o���Eg�?d޳��Qo�A�h3��N�8q�Q�KXY7��!�D>QS���t푥F{�V��E�Ӄ~���i�&���p+��x�w}y[Lҩ���>�`DQ���i��7�a�]�2|��㍡FEs���A[��8�%}l�W&��Z޸g��}�<�&��@S���&1�[PBsG��U�z� l�ZhO�'P"V0��u�+<0�J2�cE�;�d[��4��D˅�aQ�Q��|4ŀ(�Ο���9���O���
~�/�Q�O&+%9�u�nj.���A��]y��b'R���jBf5���0g�,n�*�}������S;D.Y�'�<qq7��PttEi�����1ɥ=��+}}U2�_� �#��5��D�OV\��<�[��)��j�s'���!)���C�Z_�axyz<^[��,Hs��싽Z�
�����(�x=�w�'vf�l	�qz��!q���:d��!��z�R���@��t\ג��GZ��y�LQ�#C�aQ�k�tE�p6�z��E�$��3H�G�
�BƬ|`_��Vf��ZP�d�n�m��kr��+�g�������b���w g� �M�	���L�HfG/JQò��ݴk��F��"��#�!)Tk���||�:��-��W��7:3�9��P�j\���q�~l5Eb@�e��<@;��kM�┺�y?x�_��Pcu�)�g,�`,�����3Thⷘњ6r�f xq�Zԃ�s���ﻊl�d���O�'�!�P��t�\u6@8�e�����3o���WM���A��6%���Dsf�F��Uj߲�D�/�����܉%��ؼ�-�W��N���/Ā٬ns`V�`�
n5�i�*�.^Xi] O��.�Y?��)c��A�1\��%�O�E��Q�k䤷�\t���|@�����(��S�7ISLp���y{]M���>�;�)��֗صlk�ힴ��c�����^�u�������b�=c�a�#�R-���)���mi�wU��"�amB{W?�h����ee��h��ԑ65ea���*��<�<`�.?[_5��6�CJ}i�`�x���3�����SU{,��b��EE��R���E�
7-,z�8ఊ������+�isq����?_����я�"�Q�.�f�ӢUC��`��N>�a(5>��e1p��o�����W�U��� ����@GL{�Gg#o
�Ę_=3��6�oDrg�L���c1U���B8��3!���ұ������F�=�(���E��6�Q���D�@��u������m���͖^b�m�yy+QJ�G[�FPm̨�!�L=Q�"��CC�n�K�X����Y�Z�nGgR�O�࿉Wļ>{{��*�l�Gڂ�#8�L�X�������0K5���m�l�Nׇ;��Ƒ���{[�eM2��0/Զ���`�>N'� �\a�=����aa���u�f-�P�8�-��b^{癌��	\Ix�@�L`l�֞̊N #�.go�*k��c����"����I]�
��v���v�"�J�;~x��h�W���8џ�\q����S^5�<�l�]�W<<�_�A7�u[~�zr�&���+1 :���aЁ���(��y�C~"�s+�?B�)%�*�]!y��JP
�$�T���$��i}������,�EA]��&(Ls�hC�P����C��k>��jgI�t��G܆�������(6�� �(�0�����ѵ:��7$[:h�R�X��K������˿.sW���ar}\�-�O՛�MI��$E\�7�H��|��K:{3�Û��hGw���F� G��Ģ�]�}8ĭ��<;����W��?ҁXᠦ� ���]��,�Hc44�w���B��'�R�v#�F��&��Y�f @h_�q����սi��=T}��l{T�T�w����*��ݨ��N�+x*������c��v�#]3[�yMj�p�9jM����.90�jEu�����rǇX��Z����Y�)6��p�uc�p1
��p�찓j@���:�LP7ZGk�S՛���Eq>'|>/y.��Ŵ��q�#n?���H
�B"�W�e���*L��>:o��Kаw�+�9U�k�G���({d�a�s��.XIb!��д�2��8�31�n���!�ؔ�3����j�r�"��n~$?`�H�0l������B�wi���!�݂w�͗�Ó
>[�������ϵK�M��ab�A���s�o\ӻ���}�}�й�&����z�{u��f� �]g��]5��Hd�_-c���X�Uf�W�_���a��W����x��u�A�n�.�]�\7�����XhV�GH���\�g� ���=��Q	NWW�%D��fߕ n��Y����خ+r@����Q9�0�<��?#�l��_[�Ix�lN�}@�)�!ٚM{7�`�L!zN�"M�$@�.�[&'�U�����!�	�-R��_-1�wY�|>���G���:�B������ŅM�mn��m N��g:ߋz,�pL�x�g
C��TS�+�<
��!��ބ���(3"@#�=�H��0>�����X�SMeq?��\U��Lô���u��;���"a��3���J��;R�����+��G$d�hѶ�����뮼� PV�)����@,тJFs��n�Pd2��������.�5[�K�=��H|Kp�G`%�6<�Q�n6�7�h��+䲠^_��������+sCS��"A�ۤ���.���4��q�0x�����8�þ[w��nB;�$����'��`�/�zDNŊ��7�,( hi�h7��U�3��=�_�}��@�̧D�q~,_���L3��Q�Ϩ6;�����k����I�����Q��W?�z��-�# ��W����c'g��<v1����B�\}�mv#qV�����Jo�1�o���?-�br��U��s3O]qU\=(��4h�wDK����-��!{`�Kq�>y_5Ã:��"�g�R�Ϟ�]�Bs�ƀ���$��#:������Q�(ª�M٧��WD)����J��/(�Ί�W�e��x�3�w7�i�k��8Aױ=��>���=��QU�]�!Ze�xƈ�)\p��#ع�4�<�21�⻗$΅�m3�������fM����̇%��5ȹ��C��=S�?⤋~��?��ϊ����t� "U�! 1tbE5�,�x�+p���#�5LP`6RelC%��v m��)S�|<.WȄK2)>J돫�I��bC�5)���g`�xm���z[˱�$��AM&�.�����(�5�0n餍��T�s�㻑�R��������HX}��圾 �\�Z�*�t=��k'���
�x>��&tvF�!���|�'�?�F��e���:ӆ�P���T�W%w�bz��uD0D@���hl*r)�����
-rh�"7q�YZ0��KB{�}R�:��g!QO�Y]��SP7��-!���o	L��6�tW[G���d����5T�����3b�cΔaL��3��JH@�S}�H3�0P��ߟ���Oٍw�֪�wQ��bL��U��}M�ezQM(qB�;���R%�6o_!u����H��O���t���)l��O<��R�$��;7k�ҫΡ�F�h�j39�ڪ'i`�^]!�T8y��������F}�߮\�rc�R��ك�Z�!�K�і5�Õ�p�<��uu�( ���o��9S��sL������E�g�
�|J���g����
N"f������3V'@=;\�@�r=�V���eF���m���H"��'�_���E�7'c{�P ���+
>]oK�~CV�C1B��»�T�F��'���q��.U�)��p�0�Y�!�H�������d��oۆ��z��漙5{$M�K�G��� �~nz&�W�o��c��*8/ݚ��P����aU�� �Hl�U�0 )���AH�1Zq�-*�"@ϡ���k���)�"k���a.�����������U@�S���#����p��/�����o���~*�Y�/�C�C��L;׎����s(#�8 ���w���kv�x��q���Zʉ0��5��>O��^���)jDp*y�@S��@���$�A��q�	��-����:c�>~��#����eٛ�)��a����8m��Ԃ��^c^<eDb��:̣Ƈv��TY#ߴq����	dp�u�D��4޶��ҙg�-��g��3O��=7���G§]�i��t�{"��C��x��	8S��z�<��={bT=��mA��1��W�jt'1j�lM�[E�!�Gā���F��#��#�=Xn��?f�y^�ma����:�����6�/��+�&�0��
�`chµ���$�.]M�L٭}���>��Y���֨�7�эu�Qd5�p���p������X�Q�]S����+��$p��|+�����L1i�L����yO8>�1�I����������_�4j�Ƨ㪵P��Z�����װ(��?)�9]*�U���|eGJ�uq�pk�3e��Ek����|F:V���p8]�q�2\���N��`�u*��!�+gZ%Q�_W�$��j��C:��yQ�*�P�<V�d��!2�4b9t�P&.,i$������A/NS����j�-��*�V�-�r���+�U�%�'
��XRn���.O-�T�-_|�CM@+͢=��z����.cz��4�pF��#
�����������H���jx��jWa3�wM��)��$�QӢ�-��q�qC[|���o���~��#S�.��L=n�'�+�k������|��N4X*�wi��-�Z�p},W=�6��_*���O�7<�Qc���ǨB�g��x�A���n�=t�S�<�f;gx`� ��Txg�Ǽ�5�k~C�:����<�\�����=�h�q)����"���	S��nz�jO7�B9X�GXU�X�����T]����'{��PA"Kjor���e��
���%?j��L����Gj��* �ӎ�Y��Pizѿ��g/bJV�j�ڟW��t��%�����m�C�B�������p�N��;�L�xˈ�����]�y��'�o+VJ��yf�}�\>,�E��]�Yo5�Z����
ѵ�F� �Hl���"n���R�i�p�̙�c��z���:�,zՙBԗ�
쭳�'���gs�Q�ōE�Wn��(m���\F�Z��~��\��4>`H&��,R<�)"M�|����4j����b9��7�zN�7��B��@߅�����& &l�&�%KdH��lyjM�n����c)x�8���f���ʾ�mDUHѠm0
ԡӧ!�	:�J�ܱ���)L���G*{�I��d�t+Y۝�!�tH���>��^0T@��o��Q}хnFהUv9*l�πU��&@�ᗞ�@-�ҷ��}$��P��p�Q�f
�ȩ��3g�'A�1B��vv�:���Vp���$������暿>֖��v�mʙK>4�V*���yIx���>_���C!��'퓾x��1���H����T��w��&��,�Hv_�$�3i�������!Ns�?���������(��	>� �y�e�;���)d��*d�v�"/B@9���
�k���Lm�c�K�y����ʢ����hyc�8�Ԣ�b�2���w}�
I&k��>}��0;Yu�*���H���ucר��Cl�D��$��]�i���Y��1��u�E6�iua��S���Ô����=%5o{$v���(`�b�d)��n�� Rnf��78�4������U�U�X�xq�x�ŕ{�˝h���O��:r�~���M�S>�tHP��x�҃-��P� �A��7���`��k�ڷ��ž袬�jj,��L﵁U�H��$;y���F�C�'��M͉��S��Й5m���F�K�{�#����Te��|�J�@��	;S���K���5+�"N��;�swk�Tҿ�ܝ�����_ɱ�K�λ�T�_��礠�4��d<��b��b[��7I䜹	���ed3އ�P��^Nө|��'P�=���*+��e IY��*�����D��]n��mמo{!�+��ƙ�<���Ј;c *�6K��W���S ������;��eqL�)X��P�Č���ïT�B� L�N!���@�5𞫤z�}fp���_+��S���ߌ5&2嫵�|��L�0ASlq\`Д֌Ƴi����76ɥl����v��T]k�����2��AZ��h`��r�߅��eW�۠@�."�S�J�ȁ���	��2�2)�P(Ӈ�z�|b[T���D���ꅭ�'���Eh7��,p*2�Ғ��rF�«�xne�v>�"���N#޸Ӡ:�|dB�fH��;R8c�7��8��"���G��N���x�	�o�)�ϓ�:��%*��(�V]��������,��	hъ�D1���R58̕��?���8mS�pD!q|Kn��48���$R�$�fUk����ިZ�5��3.|���`�-p���d�T%�F�����xj3��|�Dh�1�{��ΖuSv���Q݁�����X�C���nrN�	�V��φ++�,7ڵv��Ӡ�o=76��B�TA�%�@<lkՍ9���O�*��#���]��\aΡAO�wW:�ќ���&�sbE]9���c:�'�6"ޑ���~���r��R	��=�l{��Z�_V"���T�6 ̂��~����t (�nO}�Y�&��E�E��QCS�	i.��ф/c�g��m��|]��{��M葵T�ǋl�>�@��b��wͧ�������߷������3��q�6�|F3�z�\��ShI���lyq� [}�a�gWY�vk}��U�W\q7�q�L�Z�XJ������|���.�M'�{�6ؗ�e����D%�z�Y�?(�:׭E`s#f�)O���\�`lLYv>�e���T�ӿ��P�9�����$���F�A&zqD�I�dgY�T:?(߿u4 lhZ�����NK�0GNq:���v��w͠�[qS�]Qk��S��PH�$�؉ܫ���{�a��ٝ�WРh�Oil��I���pq�,�o�6�IH�-	J��r��53`�g9�D]�<P��ȃ-������?$Z��	��Qa�g~��)�^�W ��訳*5I��T�Y���m���S�A�_��.R�Й��9v��je�?a=ԅ��[�| U��Խ�q�I6[_@@"��IE�N8l�,!S�+X�����b�"���G�J"C�U�:B�	^g��,�2ZR?���.�$�8жQ�o�'JQ�9J䚃�ܛ�`���{ӥXH_������S���L�TM�hU��f㙇�����)1)ڔ/p��ˁ��Y=�WO@�N[8� �q��M��J���S�hBa�-�s��B=�w��ƍ��m��F2��U}�d�0M'��\5WVE�S�h�'��~%�L���``��Q<m8C
�;�s��0�Lmg)EC�+���6�l�|�����WJ��W��
���w��5�j:~�CZ��2��;f��!�ߊ�py�J��0���(�x&�Y������i�(뽖U¶�X��1�'
A�I>�P��9�>�^i����m���d˿c�ƕe�%za =��<"����ۃ�ꞝCR9$�7�എ��t����ڦ���ɂ�Hh`y$�҂� y��}�lj��c�h��B��Ċ+m����L�͒��J;4$��׫�����ڇGI��|�92�I�ȯ�=(�:Qы�p����W�E�~����0:��H"�G��>��;۳p` ���y��V�v����8p���މ�襤;��i���q��h[Oh\�[�6g�]Q�*3ھR�k5�!�}P�i@�e>(a���G���Y�9�а�4`��2�k���y��ʘ��h����n~�W)�@Xgu5�`h��F#�Q�?�oˉx;�Y�Dľ_s�(=�F]�}���^��s��e!���~�6���_k��-4��_(��0cfyn�x9�>;Ͽ���K|�\4e�C�x;3ܕF �y  ���Ѫ��BC	���k�C���9�.�~H>D[�����K|����؆P�I�|�z��8Y�V�7�f���$�^���G�ڰ��U��d�>H��.j���Ёn���X�a��V����A\����w� �݊���Kc��\����͂�O�n���{�_��0xtH����H4��e���z�$Zga�Ϣ����ķ��!�Z �Buf7{��i�#�A.)u�"u������d%�B���l���O�Qo��ڇ��h��˄Ԝ-Y�s#�"[�Zճ�����T&��m��g:g���ap^L�]��%K���q�P<�0D o�Q�_��|me�������lJd����3 �-�cǐVd[�R��\VW�p�K�X�b!�I��v�8y*'i<��HX������p��a�w�����:H-�*�5�8�Ŷǿ.�[�V孺l�o4�v���� �?un��n}-�]o
�:O13��y�����}S�����4��+����,u+���w%�=����aIs���m;O�4��?�t��P|^��L� ��_�3��X�X�#{��'.;"�_cn��h�o�]q�lkB�N5��2��8��<�T_�\ħ���������&��djP��/6ݰ7)�y�Y�^��|5�um^�_�Q����#�t�
m13%�e�]U���`�c�[?� � m�|8��W9�����"�Z�VOn��(�����fb��%p0LcB����x�Fﳗ���܃!rx1��Z"�X�o��9�] �"��}�����\䞱�p<l��~Џ��B�S��Z:��!%��Uxi>i�d����� V�I���Jw|˿�ߑe(a�m�.���:��On��c���ܶ���V^�	S���	8�wiђ���8,����=�R�G�p~�!�p|%<Φ�Ƈ�%Lա�	�8�;]�<�b�A�{�bd��9�P`��#Y�-�R�U���s��>*˨��@k��3LM(������k��'���O��{u-�����< �=e���"�NIU�Ks'�XL�1��z+�KW=a���mϭ��;&��B�ۖ)����[o����H����I��꾣<SuJ,���jʌ�1ɩM���;�a�A������TE��E=���b�rR��FD�=J~\�A�KS�������nkW�ʤ��<���`ΛD�W!�E���+�p�*���k<��h��B@���,v�*!���K
]KK����M�4_%o���A+�.��(~+H���i�V��9
FNQE���l�����p���ܲ��Kz/_u������m0,�j^�[��u2�F}����E��W�6�C*�������V����W�<.&�vR6�`hv����q�]Mz:��/q��?ɲ,=����Yx�/�\'i��c�Q���ٿu(����ho��}Zle���\��Q��(�U�@n��#��q��Th}uY�T�K�͹�x���v}��j��\,#�?�w.ɚ~�z�:{`�o��k���_Kv*~�J�����=�qp~w )���;͈s�.(��6�8/��8��VL~�߀ݜ�?����^� }����HOv˧���;K�a:@ E_�y�S���ń���+HᜑE�z�p��B�|������O,����T=�	^�}&��,�:�d����g	(2+vp�jk�*;�N��R_���=��0ɖ�%��EX�9ex5#^l^1����ڢc?�w� !�E� ��HIz��^7��ks��1r�Gw���__��n�gaD`Q�5[��d8	^Ӈj��]�^��c�j�� �r�����P%�-�4%�c��-��#,�W��F�w�ߩ��-�P�^�ĉ���kXh{#b���j�z�-�=�Έ\V���~�_�:�넃q���� �*��Z���`صaP�lD�Gz���K��41���_e�)^�Ɩ�K���,��ό3xE���?��(��3CAq�E񋿨�
wff���ƭ"Wo%��'�l��8IHM8�����53*�҆�5����UZ�]�s��KX��O�HRٖ�(�r���h��z-�gEQ⭭}G���0�g)#���nd9#�ȳ��N�P��a �H���&w��.����
'������I&���)�����E���:�9r�U|��h�1k�(4�0[t���0�*�N M)�n�Q�G#k2��S)�dt����ڽ�SC���� y��z*�e>i#.�8��ߖ�1P*��5�8��Y~I���ߣBޡ<>9T�2�2����&hOx�7��{b�(�q��N��i~4����-���]Cs1����P�ό?K��.������*:��0���@ؤ�D~`
�n7�>�􁢧��z��~�_E���6��t@U�S�:��}E�N�HXl���,;�nxNm��g�X�07�\��e'vU�,�a[���z�E���6��I�&�`�R�K=_�����:U���|��1(�Иc�`�X�Lu���C��Y&�TE��f��l$��X��c�:��娙����%/U}zl����FɳTuހA��3������Z�z�!�ഋ>M�j��>⫗F-n�@(cM�%����A��$�H>�7���1�p��S��s%ǧ��#x6��&�N�]�3w$�	(?��\][�9khB٘5�
_���+�4�uҤ%X$y\�B��c���nK��Y'�t���=X��� r�.۰���x�BhV��� ���C�Cn\ݠ�4����u�(�e*
K��!X���>|���f���y ��ߠ[m���&�$�y?� ��C!>^
U#4���F��x�򳫆�9Pp�f��i�!��aR���9�6�{��Hjuj+rX�_�{�_�}���t-x���]�D��,l�b�P��2.��cRv{ʃ3�\�c�б����x�3"+v���8��@��-�b�8�
�k�`m<�Et	��ֹ@GY��H��'�|�s`�nK��&�vz�w�q^���������t@i���)A��؞-JcY��Q����T���ӮZg�8%C��2WtW�� �+�kW�>�^�hY�w��e��x'Dj>�D}w�z��'K�S��Mֈ�����7�?ӄ{��gs������Jg��$��-|[J��Q�-�*ȬV&��2�WZ^�Pv����*�}?c�i�*BN�4�w[����D��2��I7��rn�ؐąY�y+�L�Lү��>x�����������W�Vٻ/�͜�����o������Ё���a@~��q}[=tX�DE��Ő�1�OiV�e74�']ϧ%#xS-d�����W �;��T�8h���2��r�*K*�$�Ƴ�e���;�޺��EU����~�U3��kb;�coK�O�x	����y���'Z��KMN$22�H\O����ʛ�QL67۸=�`�+�IFG�KzӐ�C[��1(��|���0�0߼:`��<��~��	IS[�%)�9ˌ�S�	I���PQ,�x	B��K�j)���6`
�lz�%>��R��N��^�]�v9�*�>	�0����c`�T0��B![���x{[�!>���� �m$�T�C(�ٝ��c07{�WC��s���ؔ!�7� ���ܩ(��"�-��Z�Tz�4��ǿ���w�{�E����T$.����Ma�T	� �Ӻ+��t~NS����&U���m j&G��W����!NwM�\�QM4b���0�9v��JU;����_� �����A���ǔ�S���=Uʎ��aGN.���,�U�z��EH=�s�x%�b��{�w|��2n_Mڟ���vihp���I�C����VP�ʈ�f͇;�X� �Bp�V^�^�i$��g��՛"�+��=Uxȴ�3������篟t ���E���HN�L�:�<�|��-�%��>I��w-R�a�6><��%f�
:�G[�<�� ���j, m�5��Խ�(f^�]�&Ŭ	�P��uɔ��g0s��.�͚��r�&6i;�i@vm�ID�����"�ځ���ҧ+כ@�|�Ob����������'�{�T���,:a'u�4����.]H��B:8-��!c*��Y�� �A�$h��}����Q7�2��n�ˡJ΋�*yi�#��t��(�6�'�LF�m0Y-�P�V%G�a��+�QX�7pG��bx�ڈ[B2N�$�T��a� 9x�����G���&%Y?h�J��q�!���(qǃ~K��z�o��������x;���m�!�^�]�O�,277<��,��E��@���	�D;\D*�Ge���s{��Q�5�ClDs�g@u
<B�c����q{r_N��l������ň�~ TU�*�X��d�}�d����W��Ե���
�e�� n?��� ��ҢV�&�DL�{I�]�L)̿�-�e� ��h:�YtDʪ�d}�o.�M	��[Mr^��D��2W��-�	\�k5���ρ?����.m<����|���.w!;��|��,i[����^�I� �2l��0�{;m�o!+z���5 &W�|H5ڑ�4{���7S�� Z�q��l�����c��-M�;����=9�ѽ	����)F ��T!�#�o�	*�<�7O'$֜��^�]z��[�� ւ̦�-*t�r�0�T"M&����c5Ԓ���9*w-��4X�X|£�9|��h�U��,ơ��_h��̸�W��k�3�N��ү�Dti������(:}"w�T��/&6�8��H���\�j5�FD�1��2�v-ǳY��ͼ��T�cpFɭS�F����|��;�����1���}-ǽ\U���DPPΞ�1oIg��w�!e{Jt؎��;�'�������%�i��-�7���r!���Y�׽.�VԀ��w��V5���l �Ϸ�~т��ӭ�c<S�d58�9˹�g����gk�#��Iv���8�}j��xq����!0����[�]�-��ls˹���k�x�'������-q1��
&_�t�~��>��Ï�J���U3��I���0����뗺��F�3���n!qItZ��B���8��<3̝��|V� �g2d�Q��)UB��q�e/�����k5�gu.���v���⃻��J[z?����V ���g����v�����l�0viA��^�Dm(>d^�(Gxۘ�Mr�:�
rb/���inC�C54}/Zr|&��?
gt����:�ty���b!���o ��u�z��wT�2�i>ޣ
��F�)Z8��ʙ�G´����G��ew�����]X��q���ɸ��>���|�5�]���}1cF����d~|�p��M����'�׏�u�E�c[�a��hG�j�_�;�����J���D.n��S�[���l�a$��n+����z��w�p������JV���B47����-��p�2ѽw�S\�XhVƫ~\>�v*v�#�'ȁЄ�i�_�C�}ԥ��ف;IYa�~{�f�g�� �����`��e�ꃅ�%�/�������"�
��w�͐y�5fE��ˏ���:�qb��m88sܝ_�P�D��&��l�%�p���
۝*�/��/_i��.��`�.�U�N�Cl�{P�D�Π�-Kf�����l҆�J�!�Xa7Î^\�n��ئ.���5��
�UL�f=���qw� W]�|兙w�4�����+u׽�gd����M��*%�o�RDEՊF74J�i#P�����c�zY�y���{ �2��Tܥ�C��v�.��U�q��:N*7*z�u��UĂ�+���+nL�;��Opn��HA��\�VW��4yYs�F
��'�^=�v��P���+[����̔YV~M�tN(���>� ��A����*n*Ag�7u�Eʈ���Rߕ]`�ŭ1�K7�\|����
�in��,�?���K<(�a��3=�Az�"�6Jay�����|�:4M9�Y��@�K(�4��YC部V�+HV��T�hrϟ�� 1�e��ù�5��f�4O܂�4����b욛@���F��֜o8t����#i̯���D �}��c�H�1���bS���d��f�\��[8�z��+�(~�< 7��W=�B�G��Yp�P�`L�8p��G3 F1�c��ק(g�E�x�Qސ���s~6�-��g�'Cn�O,��֚8\M+�G(9��@�De��j(x����̳_&Q!�&G�-H �t�t���ߙ�奧LJ�N�l�b7&\"Сd�Mv�B����O:y��ff2�yai�Rѽt)�.��j���ٽ�pO݊����K��1�,�V�*��e
��fh�ĺ�=���iwH,���p�;)i�^1pC)��T������Gq���w�(���z?~jo��<��������Βth�	!��`Z)�R
y<�@��{�P�|#�"Q� �O�5}z�~x��!��u�����2��q����E��mۏ��o*H�@��P˗�Ք���J�I&��7�� �%_��y)Nw�h�{{��@ЅJ����;\S��
�q,ܵ��B�mj1�:������H?m�R{��^ϩ���B�@B�=9��V	=$B:*��a^��B�U �{A�S�%.q�06P�ּ}����_❜Xs(��ۮ�]��
i����n�Cbř0O�� �g�m,N�J����rj�Q!�j��gY�ێ��
k����V!�����Y&�٨���`YBr����I;&㇨ M�u����憵�w_z	�����U��B�ix�BW=���;������M.�%��:��J]���b!W���ԟ,����>��J���	�e�YK>~��-<�b�p�>^�����y�u�B�WN��w&���n�.9g�����m�]9Q��,�?�u��h���X0�J����wo��#�C�X"��������qs���%�܃ջ�rw�7Ɖ>��'_���7t::�"��4%��_�s �F|�D�?������oĴ���ٹy\�b4-���>�E�U8'Z��1����Z�D��"1��Ϻg#ǡcwr������z�����b �؜�q9�ˑ�',�]�0$́N�$�!Lfk���ٵ��n��=)hF���-J4��:��:��*��I���}�,��[`¸�.��
�r[�V�� �N�|���-&v2���\�x�?Kr�m��te�ST�F�Lp�\ѵ�>���t�d��Q��Ā�(�'��Z���Iȳk��\���A�pRm����]Q,�i2m]<�&Q��2��pl&ypg	W�*������G�WuYMMk׮:5_mV��0c�,I�7��$�[��~h�wPh������1���XVG�*%�t��5�/A��>�X�t!��>t��o��˓4\��l����U#�Ca������7Fqe��핶��9�݈���n�,����W��~�b��>������[,@�:�	���a�����k�R�#�wtۇX9��-8����X���7�E����.ߌu��8��Ы"[0{�Ώ��� �Ȳ�e�FHJ}���6��oR�	��e�h \�Ԏ�ȹu�Ʈ��
�`a��b�K����|���ﬃp��ļ��!]z4� �Q�#������_ϼ��QD��p�I{�77)am��!������m�y�Zh����JJ�קm'I�bg�J����Q����ޢ$\���s"q� Ҏ��h;f�E�?*fb��W>1�4"Eȉ��]8�=/�m \*�=�Q�&q�A$C��>�=�?��R~ht-�2�G0E�ֈ#z؜�`l�S��6����G-�Q�¿'����I�0S�� .bJ��e!�PLg�f�,��b��[�h��Z��Mb�Р����՝�x6� 4O|2md��Ow���B��v#�ȣ���a��X��B�ٗ��a�}�@	���b��M�0G#��Q"�+�Ck*]T��:��zR��%�Q%���3*�.�n0�}彻�q�mCF����D�>�&t�T�䒤�s��i��I�+&Μ�S�Ǻ��3e�=����{�3�^�ɤ�*h�5B�ڄ��*g����d9���/���q|�x�T���2��T��4z�}��!Ef���tӀ~��T�8�+��asۍ��ZE��,��gS]|'WvǄA�X���7Ɂ� ���$�������a���w��l����Fn�&����J�k�uq��~��E$�	<XfyZb�+���r�d�;|�	n�hH�{�L\�嬳���F�=ǖ��%�� ^��VP�Ю�=y��60�����y�ަ�ͦ�[��Z����YO���� %��r�su�(ܒ��w6G�0�<g��ha�uV�2�� y�E_��j�o��'_?��f�!�𽯇j5�������l�»,�P��txp_���'�&Y�`�C�L��XX�(�w0��W�����3oKx�~����l�ъ*.��5z\����h��ӛ��'QK���b�	~�GSW��Z(W��9��7J����V�/y䂰h��w�ϓT1=T�F@.��$b�2�`+�%�e��_�p��F�֚�>S�nC��e������iJ�.y��kU�V�T�
����j��
���gJ��G��?t���n�P(�Ve<�9n��~t��.5�_&6�����tkϩ;��J�@˥E}8!�j[O�U!Qb����<I�\�:��
�� I�9ҿU����(�l4��[���|���j̑�����K�F� U^����_>�J�����Iz��62.�ᘎ�i�f_m�I�C�j��3�Ėb|��gP6�D	.Hv�ځ�����[l��G�7���_�� G�}^�b>>3C'LG(�ofX���Ɍ�v�o�2ܾp�ް�p	�A��~i'����\���>2��j��.�L�A�lY*-� W�R��?�)�6��\�G퇿0�z��T�5�QE*zI�R�	�y]�Y��e���_��5�fa"���e���6-D��x����"x\�Cr�R�|�d�����D2S�j�m��\aըH��LRC�6��@f)sU�����5uc�R�x�21V��bf�� :�e)Ly����2��&G����52�d�R+���4��@N�\�(���f60��Δ4G�UbLF�i�k���<�5��ڍ�A�Y6���o����N~Á��֯��J�~�}
�yu{a��"�Q{`�P����_�[+���ږ�8�9��A�W�<�!-1���3����B�1�j���'�7�jL�4�>��P��&(�m@��D�����Ob4Q>�p7v�I�F�O���q҃�r�;6���D�Oޔ7��xF�
#����e�<�J(KM����������z�:��:ߪ5��KYq(��^�[µR��	- ��y���X`>�a֔����DE�)�|�}��7�$}Y�8Z��w��V
w4s��2����e�B�&��d��i"7�^ˊ�b�]A��ެvVr�:�:��f��͡'��q��]�ߑ��k��I(1@IOQ��s�x��.}	�u�E�/���ie]n�2Jv�*e��5\)1]mo��?<��Ï8�J=;LT�J�+��V�����U��e�x�2�ܙP�A������a�)��տ��8�i��k�0��{#���f��{�C���ϲF+
4P�چ�BVqGAi�/ʙ�.k��P�./"�!FF���$fn��6��Hq)��i��&�s�����yh��n�0i����T���-R��[�'�01�ef�!~���O���{�@x�g��2�%
�b3�J�-K�RT$�hG��z.�̯���M}9���$�;���<� �.���_���Ok̭r˜Y�X�ݬB��>�˛�'Ճ��z�ڮ`}��nܛ�T�"K����Y%�\S������LM�V.� >�=Ȕx��b.�����33ѫ���!��蔱+Ya�������@#�j�g��m�|�)�[��!��>��s�*;>�#k�4ӓ,)�wP��'��"%�iCC�����.x�ߜE�M���d�3+����u,������EJ�0�#�|���ߐ�]qz"ߏm���,a��%,hJ���'�`{8�ZIh�Z��&hR�	oP2G��v�����2��|g4��������� �?�l���<)��~m?���
>� �6i�<sG��p�m:^�=zM���x�������ov=>�
5%]�j���F���֚�NwO��&h]������H��>�*X"O�EW�]���l�9Z4�\:Wúd6�44�'G��5B�KS��.�.�.>��w �*땶�͢������f2�E���`z7�5��U3���Ev�(r����ж�y*%7�&>\TUT3w�-~�'c�ypw��c�;g_���^�"z�9��sdj#'6�y���\�#���\>��vE&IE���=��>�U8����3yo[�fcVh���ϽH( �4zXc���͡�h���Y��V�4��db!�C}s�a H��B,�|®O�ЖQ7z�g���s��6>�w~��=2���o��:��p6p,�s�<�Q�K��8�w ���O+��O� ���Qz�Ys�hC �RH��^��۵��q�����-\6S�f;1�(dO�u4��1b�f+g˯io3��/B�%�WCwCx��@�"��H���-N���� [梼�
�5pk��e����3���s�|����}	�՝ȼD(��?��)� ����|�3<���%�1��eׅ��]]A��D2It�+��*��O[�����}��� ����p�/;Z��Ƌ8%|�<�-0�!D*��X@�,ߔ��.'Q������Bk«�<z��@�3cQޥ`�g�魣j�����[���Eə��hv�(Ȗ.e�Q����+F��[gYsǸ-���޷��$�x9^��;w�'!i�g����E�q�ۣi߽h��+8|�2�a�7h�ǘ��	��.P|EU�V�"/����T�"Bq���XR_�v�_d �V���so��I��������?q^�T`���6ଖQ��j���d�G�b�`��D�p�=,������U*x��n��T8cQ��Ŧ���b�P��@�Ox��oB9����wؐ?I!�Ȯ�dX���vx��xc��2j���7�����|k/��TP?�+�����ó�����������N�Jp���˾�Lv����MkW*���'/؋X�
�O#״n0���� y��5��4��Ωt�cH4��_�	��ФMԦ���&����kXޔKv�*D��l(���ڋr��s����H��pBSK�1���^`�6���H9����9�� eKҡ	0eEy��wYA�p-�l�E�����d�2�ɲ	0�U��d�s�L����,yޒ�F�2\Sԣ�+T�G�~_��'H�Aօ��!]�5̍�
=�����^�C�lcȝ��6IǊ��$_oLƱgi�9v�j뷵u]�T}}i�E�n�&�#F�>�ReӍ�Iir_�Dl[�Yf�p�>-�<��S�D}��kv��j�-p��4˛/c�b�;�x����jJRNb屜_HšS�b��b���� 1)��M�8��Td�@i����+���O�}!͝_q�-���m��'�z��3��[Eo�ԡc{h(u)�2Hk`rL'�j�=<&"1��0m\"�3����D��U\��-s���t��9g�Ft�>��єp��}x��t%DC_�?(�j�����,:��BWlkeȖ���lMMᙲav EKþ�A.,,�΂�|wZ�O�㷎�E�iu�a�
�t��C��y��=4��o��a$s?�jOT�'.��H�`�NHD�0�I�V�C1�Q$��[F�r�"m��|hS�H+�3袇IK6��?>��L&+c��S�X3�o�P��D܄���s��/�Y٪{(vC"�f���pZ���J���d����G$Xa�~w�sq�PP]��8����т2�y)��7�N�/���!
�'m����nf�CPOs�ج����l2���>GwK4����]W��ۦ�Y�������c�0���_�۞0̚����ZB���7�Vq�8�^��iT[dc���N���0U��?
�CF�l��G��d�o�\f}ld��U�#\��sVBf�nQ;[jm��
#Z���{��V��s�����m{�|H�A9�~]�2�a�|7�T%_�M_���f>M��x��@�6�>���DA��ޥ�`Y�_M�v��5���T:sd���<���c�6�ht(ЋZ��e�	_I@g�fM��ǭs�.��4�qB��{b�.�e����/z{N�'Vf�^*w<�p�Ϯ����usJ��֣#Y���X"K�������ҙg;r�N=�7��eB5-�������6uQ �p!���_��!�ƵTzv�Ef�}���gX8#t�O��^��A �B�vsg<Ln�=u(�{x�J:���6$�q"4��i*�^Zi6��´�u��Fp�Tb��ٽ�]�`�,�/9�1��-��&���Aѵ7X*>��%�6���p9�8S{�;E�;D�~ĥ�r��ZZ,i҄Ԏkx��YDҊ�ؿ
9��ڥD-���, r|O���c��úMM��M=��֥]u	�J�|a�"���͆�I��0oJ8�x�7qv�����"����vh�����f/f4�hc/6��Sy�S�n�_]��
4�1ϫk&w�R}��&������Ӫ�	���$!�����ZJx���e.���G ���`����� &UXCԺ(W��L����I�Cr �t�xm99��h/k��ų�����@�R�5f+�K��-^6WKi���Sp�`����~LS˧'n@�(M+�0�=Q�8�$J�czg��_D�j�X��\��e9��/�y?]��\R�_?b���1�G9}�h��$$Ql�C:gk����⩻uu�aF�1ǖ�D*/狈6��(��w��oT+;X�5|R\����XQ2���)}��ɂ��#	�l�B X���Ӯ|�TOG)J	�i����y�ۮ�";瑏M�"���U�IUT�T�����'�PU*�#F�y,zV�^�'��M���6�FOG�0�";�qE}�V�:���^_�P�t�ꆈ�
�kʃ�"��;��!�T�r�O%@ܼ��Q^.s[_e��B�g䴴�k���	wP���������	�^��&��s}����f�/F ��&�d�}�(�o�7tE�m�kȫ�6@§_��ϒ!�0F/��j+e~"~c|2.�;ՃygAn�82z|9sW��-�7+R�f�+T�����f��l��M=�.͏��:\�������������`��+�s�߳��P[�
O!hP�	E'w1�n���7C��j�k�O)]�[u�չ��x;�;����l��nYȢx�J��3\E=�I����M��Gq����Y���J׿�K��]��A+U%��C�t����@PTAa}�.b�6��Z��p�0>m|BPT3��é�8 }��A�(4�Gl��B�ӌ�؞���+
�GV6Dnʮ�/d� ��yJ�v�l������D��ac��O�҃��$�լ�6�Ǭ�ɓ�Y�p����@�ւU-#�! �����H�N#�hGf��8a��s�]�N,B�; y�w��	�@��
Ⓑ�E����=����D�����|)��0~b��hd)�}c�h�j;RL?4�yۋ�����a3���44�`���=c��]��b�/�䤸���!{��Z�X���? 7gV�Qs�Ot��)\���ʊ��~�{	X7�����~��T���<����2#�>�J�_���3��~�[M�H}#�����5��������;�u/��r��r�+���i��C�G���̨�Mx�Cĝlcz�[�c�j�y���=��%��E��Liό�xW�۞�V�Z?���ҹliE����U�A/ݞ2���$�oD�\���2�⼠���J�r?���	}ڙX�;;�F�r���0��%*�Bl>��^��)O����n��z�=��"I����<�_s8Z�n�Q�v�K3�x�W�!B���9���:x���
W{����t�xէ��̿~1�7�]����`Ʒ��������Q�ᆣr�ߖO[n%���{*	Ї�.�3�5�2�Ċ���3���.��vۉfŽ{��T���2G=����R��%�.t�9�+L��l�Z��c+³u��Iר͇<����j3�KG��I�7���趚���W�(��i���o�J��T�Y'� �*����uw��QX�޸������G��b�:R�(�oR�b��X���ߜ	"��sz�-�a���K:�<�)�?N�/a�1
�2Ztoϔ�WMd�H�5 ��ɓ�މ�,����_k�^�^���[�JH�4��@:�Xq8�&f� e!���4�~N�8��N hQY�ǴZ	��o�2�1	/~,��
e���lfbU�wPn~��꒸��y�q���sɟ/~��w<�qh�jF��o�D3ğM|�x�$Mi�t�o]>�a�I��Q5��ƸEpx?#��;���4���x΁�ڍ���8��P�����r�q����]fM?���8�o��f����-����I+=�6�|@Gw}IO�-���bH�B⬟�{��2��رG�� �o{��qv_n̘�ۺ��
Z,����?x����F�z$��.@9�������W�˱�ڀ �G��=�q���a>�%�����2�B�y7j�����̤�=�B	���~~Ӳ����h�x�r��%]q*�P/L��ȹ��'ف�8���%�}%�C�irg�b��mN2�C�����my4�[Hx-���ƼRݷ�gm�=퀋�ЛiOe0���=�E;��]�;���Gr	���s`�������˖�s�4��E��]o�sb�(fu�-��Y}�.�E�ED��p��+���C[����x���o+��_��H?z�o\ M�%�6��?S��;"r�T�>ݮ�/Td�}��+��K��F����-t���K��~��SQ���Oa���	�ō��T�ʛ�!��g�{� �/d�����/Ch��*|֝W��am����'����$��X.�B��|w����1Z0uc6RͫF����f�q0��s7��
�cy)��\y��oo�+�4N�*��X�~�����ePŎ��'$���Y�1h_�\mT�_��h:?Ѽr?m��E��k��kοZ#P9��ۉv���`�{���_Սvw��LH5L 1�Ke��?B`���o�!�U����;ʄq��E
��Ԁ�s�9��ٓ'�9q��_g�#ºA�KA�^Ϥ���������V�j,V�y-�y= �-����9)p �S>D�*Q�I^;�] �_�,�G����l�<�~iI�T��R��cVٻuN]��|�d��=��EA_#D�x���	���XIJ	0}&/A���$/�2Ȁ��=2�f��V~~龃����a�UIe&�̏�19�|�D"Gw�Cí@!��\_��"�J������ʇ��of�7��ܹ���H���<�[EE��4����Qm����\�b|㐗�3$5?�5S�1 ���z}<���
���8��Aԗ,��M��xwރ�K��!Uâ.V�j��xz��&)	�ƙ��[�#[Mj�u���ʣi���H��K�%�j��qu�Kc�����Of�q�����`���5�y�ӒU|k� ��D0�S���@�ɬBԍ&A�!o� �ڀv7�
�(5k������5��W�H���7������:�5�6��y������/�n��K����]�)�$�@
y��XC�δ$��usu�`WbH���֎	���!߆��`�����s}H��w�[�Cso�-kN���z>bJ̆l���oݲAfތC�,��� �I�uK�y1.�.��u�P<�2�u�Q,�����|��$*c�'�{��3O�.,���@��"�&'��P?P���1����ኦ>2ra�]��FC!̠Kq��Q�㤹�c��]��D>t1%q��:4>��I���'��hx�@^"ɋ]�E�]�|;:Y��c�����M̫�vip��F�#�%R��1�a�2�g���0�sEβ�L���z��H_����\�$�ꆵs���D��/x:)�&�0�~��cu/��M��k�yڊ��:g����&%E�����S蜢�81Լ� �2:�M.��a��]�Q�͓�+/����Z#��l���X�¶;F��?�8Ĺ
k.?򡫿A ���Os����R[�4쐊"�"9�M���3����b�\�T�4 m^P %��d������[�C���]�������~�'�1�~r��&/���[�����+�'ox�uf��s2�����!Cm�CL�gp	|��@���zr�D�3ÿ�zG6F����/�+?��k����4T6$�9�Sr��b(Pn9��gH@��V�0Z�`1�L ���x�J ��c�梬�S�Qc�C"���R#a����k{���-���x}$5�3�3����& ���Ò������ȣn�'f\u��4��ZCF#��s(Cc��2��D�@M�(�GBp���e�s�����T)W)0)j��_P�)%>��
�T�>���!��E�_?"�B�^y��!W_f��u��f�����i_[̬�rB��7��B��N������-�zc����H���O�[x�_�z�]>��Yt?#$z��qex��0���^��3�Ʈ����z�]u��#,8 !
��͇�69C�/tA&B�)0L;`F�PFNRP����K���G#���]�I'�G�So����Q������E%/�����.�3e����v��Jz��U��6~�f����O����_�!|�<���2�XT�}��I з����ӟMt�bE�[f�E0�m�,�L:��k�8���u��21ڌ�;�Ø����'Ak��2�M�"s�)cR�6j��m��	��ҙMH�7�C�����B�.�@�ݨ���l�@��ݎ�ġ�q�A�+�щ Jg�;_��)%8/�1*�nú��q��m��Mr�Kٰ��pbM�}~��cQ�`�)���zćL^�Έ~]��[�Ld�N�@��=ja�(�%?\��)�;��29c;O>��
�ׇ,�����8e�583K	nn�TYw�� Uҏ�U�7�8�Ҭ�n��$�kY1[%ggkH}���q,��l�D�y�*�>p��Z�`��#0�8�����ލ���!��z"��h"ֻ�y����Ym�/��E߻��W��v_��ƈu��_��/c�!R4��Nq=��F�Z�-1�=��%��?�J}���;�]�FH�	̶��f�׮Ԇj�f���쿍�]	Ksxϑ�|�(=��M5!��\��{����\�� �Vs��0v��bX�h�<�L�kkl�l�(:J|sz��3)z��-��&�ց;iY���;��̻\فr֒X�eg0��U:�H绡�!q�=�囈c��go�y�F�s=�N��6�PM7r2���G���X���Ҩ�M�{R%歅a��?���M��c�׈D��{kk��`û�*�["k�Vmm��մ5Z��422���D(=W�x|��곱�.�@7�QM���@�����!k!��vU~	ME��z�k�\�J����q����3��	��<c����o��Zח�S����O-�`޵���l+̥�rw�oܛx����g�R�ǽ�T#���3c�Lu�;��V�Ę[O�
�'�\�M��(y{�K���-č��o�!�jK���Mq!6���5	���cHſ�tJ�:#2��3hp6g�P`��
BS:�끥+ӭ��m���dP�����3�U���'���3�w�Z%��.�@-x��>�n�v�Qi(**w��۵NE#�i��_/ZL�aKi�Zo�Q �IY�@�Uq��BM���E\����	f���%F]roR���6�Grv��O+���!�f_�$k<�@�|k��+�P�7�`���gu�ˋ!�U�cG�P�(���!�~ݡ��gK¡�lPd�W<�l��T��ߔ��YS�3��Q��-x����w�u�L��i�&J��V��\��N�!
ҳd�p��Q�MAI7����q�ߙ�}�{i��S�-�c]bo���hJ��PhiJ(&��o0�y��m��j����vJO���j�U�	���z�-���qހ���I{iJ/>PTm��	ZI�E�"��qC�9��E����d`�894t3�J
�R_U��pd
d���AV���jb�=�&7���8VB`j[y�A�P���+�����(o���E�T�u1�O�x��ß�����y�]��(�����a�5� �z�2���$~'��h�(��-�G���av�����KQ8���HRNRs���6 1t��t�U�����ΐZ�6��	���
ʧN<w�����S{f/��{x�V:�Uʹ��Wu�
5=�����H$���g#0+��NX���f)DNwu>x8a�%6
�+�%�W)��<'o[�p�`�H��㚭���w�/6&�,�e�x����a���-��$�F��x�TQ�M�D��8��� �4�f0�%;���#^ហ,E�Bմp��ԽX���a.0�O[����G ՞�W�iHr��񌝛@��u��nq�1����$=Hw��[���ޝ��.�m��$I֒��Z*���Ǩ�E	���O"�uɢI�~��n��g��~�8�3K��Ժ��/�;�˵h������R���}��*����4]��Δ.�Z!<�� �rEsލ��S%,uT�Y���r��!�:ͤ"��%D���<�G�sW��j���%��S�u�<��Y�����0Ua��GW�i4���u&4e��#�'��Ϋ����m�j)F��;�.��bY�c����(���y������̠���9ZfB����j"� eI�ک
���:ʉ/A��gq}���
�.- �_S:C��_�P�d�R!Y�I0B�	ё����:��:��V�mLG��[�������z�i��v��&��$�LӋ�=LƇ
����V.5�"�V����$��y6Fsm?��7�o�f.2� ���h�UNV���4`?�����D�"�|�)�ݘ�ڝOI��&���ei@��{�xݟ���ܺ@��⮜��(��7f�V�f5)���|_��z�Ե�݉�p;����jU�/���%�x�f`_=R�v�s�-s:�Ɍ���o/ӟ?C��$���ª��\���d)��Q��/9���wp��*��u9/�KO�t;�Y�_��P����'Vʪ�$��Q��j�ǋ���z4g�c�SR�t�6*��/Zլ��urx��S�CW|%��,��w�_7�L�sʼ�sgr��r�ڋ�b�?xJ�jǷ���ϓ(�R�� ��𖯓�j9��Me`c���c��?�	��N�w��î�	%y{�#ߛ��a��7�@f�w��!W���Ƚ_/��+A��B�P>
(��"�����:�i]�)E��dz�r?9x��?D8���iYь3H�W�^B�]z�u��f��G�A�s�)� ���K,
�F�YShh�}�%�z���tp�P:���S��m�f������ĩ삘�<Jd:"�ӣ���^D�;iS?<O1ťWӜ�G#��V֤.�;4�����W�=(yV��Wٸ+h���jDa"M�@z��	��%]Z�� kP4��S��T7lU�s����2`
̸��>��g���-��[��VJ����M�����tt��@-7_A�������s��D�lj��x�o-��D��\�,
����.h��ܼ�vwyc�Kmc�c����Ah9*,hK�[.L/+�z~l�h罣cǨݴ�J0�~X��h�U���b%�)iVJ!q�pZqf��҈A��SCV�j�]~K�"uS� (�p���x�Ay�vhq^�-�Ֆ�?4<-���ʡ������%�G�k�4�R�S؄b*D�,�G���c!Ȟ�/P���([\�S�t�m��3���F=["m�(ξ�5��5H��n��� ��V+�d+���|0���i��<ya����s��*��>��g�3���N0w�T̤��׭�+�-
��vQn�����f��I�t(�� Tg��@��k�[x��hH,�x	�0ע&����ۡ�;�i�J�{�k�x�iV��A��e�'Ǫ�kc�A��xe!��EB�DJ�~��^/���fwW��Ӡ��k�>%��)���	�u�|urpv	��W4$ފ��R��J��������FC2rD��jPk���3���\k��ǌQ�r;^�6�BH�~)3����S�n�����$��W.��j����0�V���GZ�ƻ�#z��b	�9�m
��>�4U�$��I�=ꛪ�:_�HP�nA�%�h|���*;ÀS[�T�ҕm��}�5�OA�!�H�[%;^���2��JL��a�YE�>.��fzk�N��a��+��<@���v�a�R[���EB�O���E[Ui����9�F�-�p�q�uN����r߳��J� �@<�*�Y����lCO����*� _|k���S�!=3�������<�j��I킟{�#��5M�/�$;Qb�͛V
�$-!����L�f#��	b��Yч��~Zz0=|~2��U_w������b�,KqŇ�w����cW��z��Q��c� �����\T!��\W�#�Q���HS-6�봨�-
�=e�E@��W#�]��:�q>+d�&6�\�=�h���!ۅcQ/j��� �XM`�W���wR·�����6�D/ч�(@ <�j՝2�8H���e�,��s���xki�ŹB��3�4Hd	��=�t�,��F'�ԕ��,��xu�`�6H��4/��m�a��C� Ǎ�wYc	3��&��pJ��y=��8�T��~����ts��Čo���Z�r��?����:��]��֛,g����/��:� �����Qv�����Y��i���1�̍��5��iL)`_����{�/2�#�QC%�D��LY0�q�K�2���ń�2�-��s@k�U� i�"��)�<���9[ V����}́����FݺR�5�y�+��֏�s���<�������wF�A��I8�?�2Ax�)%k&WH�8����ˍ�n�z$�b�a�@��|#�]����w?���/���f�C�E��G�\�><��G���k&�U���xA�-j�8�4�a�U� ��s�NT�˺.�D��8T��m���0x��vz�eXAޯ~;�|gQ B���CE'!�r��@��2�?3�1��n��uu��e4�y��ʿ�N�'�Y�t(�nzcF.�h���e+��>�2�$���ϧ����~�6u�J�\ڔ1�a��\��	�Q�j�-X�_��H�ʯ,�����d���/9MG�g�	t����P����-Z&<�J�B�����ףo$�s� ��c�>A�:;G�޷zvd��3	$���p<.-De�N��6�Q�x���" _�bCN-WùCak�k�v��J��W�r���w[d��8s��S2�<�u�}�2���E� ���ۊ{M��j�1k�z�{\����	W�=O���H��½_�D�&)�n:Ԕch����3Y_��.x��7Q���Cd�+�F;z`���X�K�����5�F�8�D�i���N� ��h�T��EWP|d�dyV������� �#E@|�)(]
B�Bu�i4��u-�|=��d��jAt)ړ#ﶋ��ڙ-��.86�>QRP�i�l,y��$�4�@�.���ϒlYBt�q�M'Vٵ�AV��ry�g��ܑ9Ql�\/@���=I�@etZ8B���0p7Bޯ!`]�%����;m�\�,}	@�'�5���9���������qV��"�n ��h�Բ����!q�p?}�!�wg6�= ���ݤ��g�IC}�}q�s�����l��-� ~���`<�oN��r}���X�fU�H{VƼb��́B�2cQWFْ�����'������ye�y��=�a!���:u�cm��9���>�Y��%eU�a����ڗ���2|�Tx�գ�#�������$�����3!;1(���1s�o��d�����YC�N3�M��,��t�)���%�{^'}�ƺ�=�Lq Ѓ��<(
�*5D$�Uh����ybݣ_�� ���d�f&�+u`��p}
]B�nͷxB�6���H|�Fm�����E,S{z����9v�}٣,�������&J��2)����ϩ�!�:f� 5s�f?����W����V����h�*u�f����ݕڻ�L2��f]еBY�xCwM�b��/(rF��˒��;����d�ఊ����%�+�q�7�F�;+�'⊽��X�bGj=a�\�~�YJ�����e-U ���e���Jް`�.��2�wv���1Zg��D1��
���qJ{��O�O�w�g�h�2�l�����L�B���わ�O������.,v϶���G
���nR]F�Έ����2뒁`lPu��$�B^M���ʲ�&���We8c�?�uf"x"3�S6�ѱx�= HD�E{G��7���&���䣶�~�����+��Hޙ�d���sq��1���z1�I��:�TC�=|\��:�k� d{
� kz�!��,1�*뱯N��ӥw���h�d*��I�x�
c���A�6"���X�5���J�>��+S0bW��^Ф��5;�W
,�B�̮\�2 �Ӎ��E �K�}g/�4��������U*��CK�y�uF��ԗ���߁������R���H�����٘�"rM��鵑go* :����y�����qv�@q��o~Ҷ^���s�f����t��>Ca2�a����ƚ�C�U���}tF�Ky˒q��oC#@Di�r�p���C��),붂=�
qIx�1���<_xuM��WH��Q���(n�E��_t}�����Hō)v�і�ޟ���<ϴ�Hf$���ll�&	��`�����13xsTX����⋫�\�����D�}�2�/ƻ�y��;���Q�j�ZrGQ�m<Rm��*e�$m�E(��,�=8&�^H�N6��=y�M2�̾�?Un�_���d�8���)���Z|R=��b���b4�3�ӷ̍����ɶ]w��t$�2��!MOHU��P�2A`�kf�Q�}?>bȰ���c���m�0�_�BPu.�[�(2;YE��,T�1���?{�+Ņ���$W�mc��a��N	2�'S�G�$�O�j�-�/@�R��ۀ65l�V~��M6=o�ʣ�N9����ŒS��L��>�g��љ/}\�f��G��)�3�b�5L'Ԗ1����k����!7�C�b��
�����/�Nd����s�{c���gQ�}�<#M[��p�f%܊�I��	ke������-�Zϙ�7�h�5��{�o-��]e��w�)-8�k?ɵ�&o�e��l��TX�]W�qD �u'7�D��{EH������G�dz��%�E�u�\�{�:���r��Z����@7��3�Η��,�t�R;���'�,��v9\&h!]���8{�T
����
9�4H]�����r�^���S�5��Ǭ�#�?�oq�GH�@���Ԯ��p�L���q��%/u:��
�"��-��ǹ���N�r��� ��$��ǼD�p����{Й��[؍������F��.��XdW���b~�(����N���0-wƶ�J�_�� _��f?�Ղ�� 3"�ozܵI�w8��4*a��:g��<�'|=A�WLuf�T��x�WӬ�n���Ѕ^����Hk<���˥��Y<�e̺�Q��=�"_U�7^�P�`�}��z`���C���x�jw���F�RV��px�'�o��UZ�j�t)��_Ռ���R�^��3}���I�@��V�t�S���A���J=�Ͷ.8{K6~1�a'��Ô�G����~Ic �2��Ԩ�U�[+[X�/k��	����'w��Yg�)���YST�fn-��Of�7��������h
N[���пr ����`]'ąs��T���љs,*�
/�p��ϻ@v��J]
s�� ��e�UbV�*_Z�ÍW���arg�u����P:F�� }��Ef�����%%���<k
5��3�)��͇�z)V8JA/T�2�S��!
��G0�N�#A1����X�ax�3su4���������Kq"��#�G��w3dOذ�����g�cg��DbJw��\��bG�����ͩ�X�yx����͡ܫ�)-�NX�F�Y�%0Z�(U|�W�Z���?YiW�r����s,ğwD5�5Vu��*<p�2L��s����?z����Vw���Q�&D{�5���Za�z���7=���s8���B�vfg.	��u9���70�{dkQù��|!֊�"�l� wJA�\�
�v��;���?��nF2�=������v��˫��@r���C����>*f���+�S9D�TW��$��#+Gu��>!VY�o��{6�X��:>Oj�U;0!�w����lR�J��J箹D.��(f�&t�&�k�UV�fO���/碹S������<6G4��_�{/c�~��z��pw���������۪�0���WĠu��Q`��mD��u�^��&rM�F*A��4+����8����)�]x7���]��u�q��]���0P""�>j��y���wn��B���7�㋲�-������6��A���#'�7{*�x����) �sZ�≞f�}�m*��f��
y��R����_\�6��{7W�p�m�3%���=�w��֔�Ԧ(�Z�Gl��)�6�2�$4Mo�)or&Ofz
�ja�(~�&rݾyNS��w��k��Gy%ϩI>H5� �q��y~`-��>⛔�^Bk|&4�gȩ��
_,A"Ҹ�nA���� D̓���OC,��bY��_+�\�a��1j�8���m�M�`��D��O���E?������X�$�ӺvЧ��=z��	�bEퟻ9=������maON'� �I���+��L.bE�.�V�NG�	�yqk�0�%[1Xc�k���ۦn��>����Mq�/tmDb0��X�Y��Nֺ�yW��oD�Lj��E�H~���AUr����a2;��2�,�'<����5v�g�|*W��ʦ���(�F�~����1��/M��w�.o�����2>�P*��<��׳���kFmhV�X7���������GUсǮ�A7��[e��=�)���
�8�s
ô,���:�?����EU�`P].����w����*@�.��sС6r�73�GP����朿W6������
5f|}~J�[��� ��=�N�|*�89���	�l��+^XF�U#On��E�4�\�֍�s��!�.�5������n�j���� P�i*~�	��u']����*~٪���́�������>�� ��@�� ����z��B�t����N��A�����m�~P�1\e{�qǮ�~���y�T��ӟ=�盻ؙ,�^��5��=n�2�C�%�֦]����$�w�!CH�7�k���ZՏr�C��E�[�V�lu�st��E�N��ӗ��v�E>��qW�]B��m�ݔ�t��D�ɉ'�C�
���y��z�a��B�A氫me7M�ֹ�3�{S�?<����(���΅9�zC����x�/Lva)5��K�T�_"���s�'*Q.6/2L�i���������������^p��>w��gf��5$����Cri�ɳ��$�WH�7�5lP�Qf�q��*��N��gz��6�*Q�cӖ���6��$��n�h���ڢ�^b���3b髸��V4jī�Az�P�j��Y��\�ݲ)Q(���K��������:1e��J���K_�[2Wt��u�3i|��_����|����SXt@KꟀ*��w��	?�������-����WX6Ơ:�V��S�y+9g"�,��$A��D�>Q�$����N�g��ri����a� ��3��&��d�Z��0>���3� i"n�-��\�H#P6n��1��� �W��L�I�?K���1vx5����
 WRu��%�����\�gw���G���r�>��v�8>K���r��6�sn7����<�e=��7�r���)Y�S�e�X�K��}v��T�m���dD�Z�(���.�����V���	�[��ǁzW�4	;�$�����f����A���h� {�M��x��υ�y��럛K�Ǔ�EBK��<4_��cx��_A�aֳK0��1�J�%�|lݧ�	[>PE����Y%펈������cM�?���B���JA�i0����p��WaX;NS���q���]g;*�k�ysLv�h}4K1��|����� ��&eX/`��Pm���ܾ�����衘O��=-��Q��'��b���?�����!Ph� 2|�H�u�	&���o9}l:0�B����>��/�B�C���"���zo���\E�OvZ�&�Kx\B���1&l��\X�u!)����i��[���UQ{�z�V������FY��6{Z��n�����yr��^�/.���z����	0�d�d[�8��u��1�޴���3�����T�!Fn������X����|��"��C���:^�Ƭ0��n!�Ut;ڐ�O�S,v,�����:�qc�P��N���e�J����LgrС�ڒ֪3#B�Սj�y���]������]�Kw��sD��pL�o��'m�J���ךmoU�����$z;��,p����I ��"+R������ׯ�䬌 rӒ@(����3�Fpͤ