��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\���V�fnvx��ÍG_;�ȅe�~�>���9�>��Y;�0G���O��������Z����]�%��������#ҺZ�#t����כ^�$���6��	��|�2�#l=b���/t]����cy4wd�%N�|�u�!�Pq���v+����_a�K��5�c�+�%_Y@�g�����2>�7T��߯bNq��
һΑ�s}�\�
GS���xN��X�����H��Z��Y�,C�tdI"��E������E�����i�q���0ubJ�{M�rWiGa}�4o��O�����>֦�ton="�K ����j��X���r�,s��ȳ�|��楪�Qt��s���3�Fս���=H��a]����w��6m�� ����"�[�t�>��y���@p��(�8�O��!���3�N�{w��?0���}�s���!͇���=P!,��.|ܹ-�EJU���6d���Gϗ�c���u�h�"m��e�e�3&�ڡpgIr~���_�S�w��f�`�����<!(
;���J�z�c���M�XCJ�6I�+�1Ol�t���f�$l,Jy �p� ��U1��^�C#0Y܅(��.Ͷyd��`W�7a;Ƥ?pc+��=�2�h����}FiRl���Mu���KA��1�������ć����?�0�����e�����5�Vi��p���-��g�׺��T�:�!1q�W:��-wju��Pg�O��̾g~�.m%�����y�_4O5��6K���m��H.�����L~5x�8��m�P�kRvwl�6��Yi�aC9V�K��Sc���"�e��5�-$��?�Ebb#�!d�U�
�ݡ4���<��_i��IW���Ns�<t������}pt����auxW��o)��3��P��[+<K�Y����#\�H��n��w<C�*���`Q�g�$?��ɟ�2b���ّ�j���ç��������+,��)�э_,����3�*gc���]E��z�9P��×E8&�e�D���8Յ\��B��$�g�.�qi���Ì ��&}�R��MLP�XM�����$��Uly�&����aX�wJ#��r�g)-��P�ۉ��s'�o�Y�lj����Q��ܭy��*Z��5�����p���y:�� :�=���C$�a@�����?��ɖu���T�Q��h�;��G[�_2��V�AlBE�χMē#b1�5�kIg�����C��+���0�e+T�j�O��_�7������-}�u��>�`��2=ԓ�'?����70xrx���͔�ek=J�� ��VM�m�Ɇ�;]�k҃3��������~����_g[ ���r�ofNO��FA΃O'P	N�1�s����������Ώ����6A�fx���IF���
�����E�OP���"��qwA Ƚ��]tG�Z�fR��;����v���&��jh�x�ZPN���,�J�w��q JX��z!���qTg7X��L78/K5X��W�p��
�ޫ_�;�c�㋓Ɉ��a�kE%t��;'>I!8�*S��Y�uD��`İ����h���n��B�����	 ��tZ%.�)c���EӘ�ӥ����X�.(R�����9+!X�y[��W��CX���?�7+���w>za3R����x����	�?�i�Qk��u�i�%%�4��R@�X�ο�;���r�1��Wh�6﯐GצdՀi������=_3�&w���Y���h�+#	m'JP��{�`�F�&��0��KVq�cA��E�CB��~5��쮊Y��S4��)i��ϴw�Y�#;�P�-���������%2O�W�[|�>�����Rʔ�;��s*tT��������v�ԳB��*�CGѧM��=���+/�y"�� c��#A~������R5�9`I�=�A���O��܃C]���a4���\c��ќ�;�[�qf%hǒ��)c��	�{�0��s�G'����L�_�o�f�wNǻ��f`!���D���ٌ/%��t�,���q�#0��>ɂ#�,1!!a�8_�>
M��B�eR誖<��V��eAZ����W�~p	-���P����� �9��Q��aq�Y;w50�In
l�!qa�"Us��_:��o�G��ʑZe65a�tOn;L���[�;즪��ό���>��n��:��ܽ�uV�� �e�"%G�+U��]��L��.�l�Z(�~�X�M�����h��� b�����)Rj�+P�\{�ݽY��_wҷ.̇��%�����0�\�˳����)�!$�U{&s>&`!ߒ2ԥ�j#��64���������[c`�?b��?��Q�3YsM�*I�j`]gg{ը�|\*����D4=�B�,(�F���w |P�5��,\z�b�~|��ȭdy��zy��ƿ��1ۡx����-�[��c�}��K\Q�#lJ�`��Z-P����(���ٲ����L#n.�H`ʓ�v_g4ZB���^Vp�Ν݁{���Gc̝ܱ&�
b�NF�톽�f_�<���T�@�Y�fs��1��;s�烙���4c@*ʉ:4
�ZNz`��{�S��^������&�e�swq	[��\b-���u�����+�^�xeذWվ�p?�4�4�Ũ��)�Q�
!3I�D�2�8��w�R����5X��{���N�2e��&��|�	���p��5�H"�`s	�^�0�fcY]��0
 "D������_�%S�T�����-�D��+���.c�r����ɶ�@��� �F$���HP\ ������Y�P��j���9�
Ӥ����鎰Sf_O��J7�|�Yx)�&��"=���nImA���B�5Q0q2qx�ՔlMϰ�k��n|���c{\���}vL>�[�c鈵^jg�"2��
��͈i	9�go��P%:x"����J"=ܘ�Vy1��옖�w,ih�0�.Ж
�x�������4��P��A��gTR��:tk]խ�l�\����-�mk ����cᲙ��&ŷ~ `b=*9�Q>x�<H�>�|r��0�㛟[�%+�
��&�1{y!���kE�j����V�*7Uo�A��۱ܪ�Wo���$�4��:ᓪ�6G��s��Tǀ���z�*lc}�����f�X�Y��`�V���>r2rO�W��ƃ?j���1�Qp�V��_��޿�8Z|��j�J$����NW>�Ā8���PvtN�ވ�;��vT��K'���J3h9��|����ɱ"(o�FS�r:��7g�(�z���"�Ö���@d�-X�V��4��<�{ݍtN{�
r�f��q�7�v,�߿�ueմ���G�?M���i��b��Z�U��C$)pf�vͧ�~�4���`�>�pR6�2�X2�|�Š���m6&���qx�;�/�i<6-�S�v�V\B�7p.ڇ�����Ϋ�`�(��H�+b�pd[�D+j��Ϝo2�[US'_�=O{j'��|$��/�U���#z# ;��Uk���t�ǊbE"� ��pT[�tK���C�ќ\(��0
>z�����kݔx������%��N�L \?�n�B�{3� 4/��g-"$���za��ډd
G?s����s�a�Gְt���H�O��j-a�2� 5�, �]s���_Rc���{�t��V
�@�k�ne��x4���6�y�H�,U2�\e1̈r1Y����	�8hiVR�}�J7"�l�?ɯ�h��<~�h���1�USzu�&��.oIf�YC�t��z�r�?�+����"�gL���a�?ԃh���2�����ěU��*�w Һ�y��QA4�ij�w`�ݼBc�W쏲�Q?�D� �����Ƴ�f�&5�}��
��L#�܊l���*�I{�.p�s�ٓ	�}Y��·Z;���D��[��R����όHW-�~Z�1��aq��ͽ��������zm�D��+BV�����'��}ģ"�o�g��iwx� �
}cG��m�V q�&�E�}�\��Z�>)q�Q�}ӱ���L6�O��x�Gc�����V�\���ӳ-s��ݪ3oѮR��s�)L��b:]J�]�xa.�o���)�&��V"";���f�I?�%G.��~ů#��q�ms���߂*�(U��^�zV���6Xml1~���x�9߿�w�r�����}\��EYO0`v�E�J�N�����֤�9�o��]��=�r��81Q��bIu�o��Q~�)�G�H���tw����E��M�w(�{����H�� V�o��(�����۩��`#{�����ʜ9D��m�]"�T�m2;�7��{,Ah�"lF�q;75�^��8�?����r�LV�i������U�j��%b��9N�Z�PB�R�& �'ɜ)R�]l�t:��:n�j	1tH���S/�9������$F�'��0�lߜ�y�oz��l3�1 U�K��W�Ϳ���G����� eZX��N2!�֧����+��K�N�褑��m�=#��숺��b���;jt�
��i�U]��Z�ީY�7LM܋�..�@�N+�J̕O�v-�Ys?܂���8�5L�+e��t;M�楀-�l����w�<���ɦ%Gvi����o���5���hr� ��&˸���w�]���N;˚��.��~�DeNj=�j�T�`%�
.@��7���4�2y���7���b;��q�����H�Un�"