��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\���V�fnvx��ÍG_;�ȅe�~�>���9�>��Y;�0Gfz����+d�hE9=��Ys�����~�F��Ke�e9&�#;�4J̱���v�Ga�NS��(���\������������dk���TX��n��X%���G���8];Na�ҵ��TO��؁�$�[��kE�~C̺yG��1gM��Ǩ��|��(R�/|���Ƕu����XR3�7��T�r�qބx�)�f����I��F\>�y��@(�K��B@@�h"�Vsts���"��eN,��o�}�����W��V��{��]��(�7H�H�EYa�	�;�G-��mݺ�*#��d�I�P�r��H�A�h4��õ7E��G`��B�*=޷���:�$�Oj����W���9C�I�1ф�WܽcED4�0E����f�xAoiQ@W�<�8��?Q�D���B�.�4�ǡ��{��D������V4`�"��`DX�~�;�9=���o!��} 髅�=�w;=��	�֪ȕlw�Q�.�@�]�oy���w/s� O��3�k+�v�S��CSz�_����W8W��AQ	b�	}o%�|:D0 �����v���R|��i�ȕ�m۵�}�%7��X�%f���\��:��t��E��O��@�r�(��0f�9@�S8&���bƤ4���d��Y��[�������R����c/Dz7�g����;�k� s����̍&T��,4�S�.�5�<q�z��o�}y��a�w���R��;�@�{x��5��{R������ʹ��j+D����<�EK�v���� ,."5i:��Cu�eb�,�O�I��xW��sTW�f��$������bkڷ������p�R�<�ʏim��B'�ڶw����>~��ڿ��R�ɏQ:��V��)�,>}�
�L1�p��<������X[4 *x���;RK�Hg��l�c�̵�ߘ�ĂeӀ��j�}e�'y�wh�Ptԡk���%5Ί|��e_F�@�I�s�'\��M��L�<7�fɨ H�pE��m�y�b������y� j��z.�"B��/?*��H�dјI;9�[����B[���^��Ъڨ����~��q��	�?Ư�y�_�E�9�i��y�k�>��k�sԒ� ��*�"[��0��h��4��r���К���Cc�R�����|�>�o)���=t��O�_�su |诞I�)߰E�W�{k���:���B���z�t�.�z+.��!V���-R"VE_�>Q68*�Z���t�V;Y���R��'��#|C�*7�M{���#�f�_���w��5e>�^$f�K�n�tl��x���̽�z0���o�K}_Z������lk�.u��4ĖQ���y�)z�@���P�;�GMѲ��������tw mdc��?t�����"����B�a㖃��߲Q���y��?�qH_���AiA�qM� �a@�r��:��R�D�=�E����uoM�&НQ��6r�n�E��Kwk��z��D����`�7������vv���}Ԛ����c���-�U�a����]�Eξ��"�UՏ�I6���_A�`�'�ߩO^�L1�Fw��t����D�(�C].\̉���i���
[T��}ץ����>���t>��[�1�t�[-8���/�W�$�4%&����r3�s{|'@|B���~L1��^
*K���?�ֲioJ�/�3��ηG��f�}�~�ϊ�U~IF��*��ϐ���
T���k�4�
z�M�l�u��	����Ӻ�9�H"]�����
��	��9��U�d��ٟ��(��D����]�D[����~�)0�C74<NQ�@}F�khQ�oJ�p,\V=�L���� ���IQI�i��ŏ�aÊ�V�����qB�}PY�+�@��m�hx�W��~�t�ҟ�I��u�03 C��B�d�xG��Z��UsGK��!��3
m�� *@��@����S!�����k�V��B6��}
 �%�nٷ&�ͨC[��~{�2�Y��JɍD���v4 2~0Q��E�0�Ƽ�������x�+_M M{�C�������JlL0&���xd�vj=��;����꼿���Q�?��=0|	ĵ7fs�C�e�{��g�_�7�S�/��y;<٦
�.rm^A�f����t��/�������e�bn/.����;��9��x��6�>��?r��1���v9�,oY�hc��#��� �>�m�_BR��_0��5�Q�u+H� �20�׶(AϾZ�x�f���q���X�����85fp[+I��j�%�>����"�66�P��8�i�@�>+`�9o 8v��3t5���dϏ|m#F���e����������r�ǽ��[��hb� C��������B���H����HhDG{���o��l3��%,ؾF��~f�XX�ߜm�)�t>�����.�(,��v�D��|ş����L���s�Lp��q�6�Pn3�]�Gᣨ��]C��G�er=����s�O�j�W^ʁ<������@��U�"���L2hb�,�:ˈr��o]�0[�7嶮��T��d7�#�:��Ⱦ�R�o��(�$�2n:y4���C��K:�p���g�x��>�R�u�L8��A��.j�<�S�v}ZA_%7Ժ�R �i�5Vl��l�v0˝��]V�:)k� ��F�x���W�*��R�[��z茲.FfaI&oy��P�
ԉ��/\����Ow��H���F�EV��c�R���a��;���7�X�l2n�� XЊ�T;��L��	�jR{+�t�Gh#G9���wEB�*-ح_Sn0[r �#���$:����JǩzH�I��3xU4a]��a�!;X�M�X$,#���5�B$��c�*�W�ZƳ��I�%��Ym�
^�ZϘG�Ed0�4C����I����C���-w���ÃI�iN��Zc>�3�h1�V��0M�9��|z�y�cP�ѻ���5c�Lbfpjb���3�#�6����mZ%�O���G���?z)�:�%É��t�E�lڄ?`���ȇ�3���
���U{�[��B��oc�ڐƈ%N�a��ZW'/F #e�H���`
��[O�=�ܰ�~e}����I/��#4��y�Ɣp�υCr��"Z��USЖJ�a)�8�;f�"O�A!L�g�N�'_�XbЙ�<��&���/���F�}\M�����R�bp�`47��_�X^�hoh7�?A����85&��X��a�O�+��$�+.���c��f��JhV����� � ϡ?#���\4 ���wL:?=#�&�g��?&��&ݳ#L��R�(��hc�ߴ=	�Y� �3�n�KK<�c3�Yl��w����K0;z�/��c��f�����7�����Q�:�#B*�
������b\'�ū>��ӌ ��ن�p��O��hK�� �/D�/�*H)_S�DM�o,
�+v�VF4|��Fd��MF	��#j�U���&�9w������F�N{�3j�N��h	X�~�'1��(�)�!�s��g���� H��%ǛEe�zTi�H�u�C�
2H��*a���6 ����`{�����������I툷N�%��v�Y�#�'+�6
��]/��x�� ���2������rCu�?�o]2�L�'3d�:��֘����Eab���k���,��,}��Do㸶������1�ߝ�/U�}/�v��8V��-q�Ʌ�RC�8��L�U :U�u�c�����ox��C��߸��W�F"!,�R����{��Os̏�>"�x%xk�9��������;��~�A��HkЂ�wT�4xr	Dq��k���%f���f6�߅]���#PG@�u<�pSbln������C�	N�C�X����o�Na�A������n��Ȃ�>��8v��T@�ikg	]��A�d�		�%��aR��^: B�<9�/@(��C[��uK� �������������濕C5n�g��}�iq1N�wz+#ʇ�}�dȨ)�����K��c`b<�����:P��q򇾫0]���MS���[�@ Z�Am�Ԃ��+C/�υ� @��"i�G>��ˬ2�-Q�)^��n�$� �w��_*��0u��ű"����+�$���>�����~t׷���L�V��Q�1���:�$^v��.����T�ivm0v�ٚ�ٻ fIq9��B�3 >C�H�/l�4�-
��8�v�d|�+WH6�mp	�3MT��.������T��S�0����N�V��2���I��	{l�n�" A��qw%�)�z��3��-��e���R}�bF���O�ǭe�~e_u��!}��'�/��Yh�B�Hc�(�y&-�ٽ���I�9�p �c���"z7��LE�ɵ-�O1����2�{P���}��R{<c��S��
�	�}kCI�G��]��=����};m�wA4$�0(�G+�F}� �S1"N�f`Q�������jS�v���Jv��b�s�R
ҽ��������N�آ��wN��y	���Z��Yӂ�g�j��K����K���������S4P_js�I��H��*������B+�s?S�4Wk�v,�p	p[PJ]5�H^ǚ+����l�";q/j�}���-��>�K���ܶ�|p[H	ۙ�#2�JLXӱ^Ȳ�����vT� B{�,(�=���։�k�r ��a�������SEP��f'�v3\�d�%��93R�1:�2�=�C��W����d�=�j+��Sl*�4��?Z?`]�:Þ<�Mg�=g����W�Q^�PL��m�^�6�|gg�Y�e�d�Vy��T���K_��դ�fu@|OZzt"��[�;#��-�D��5����{OP�Z{�.a���J��C��T���̢s�JhF��t7&�?�5�,_����[=Mء�qSg]_�Z�Z$�����40]3����rROV�ֺ����<K�-�2�8Ϸ�1ozn��P1�t��gzM���}�3p_��qI�F�����HO�8����5��'��##)��R �f6�%6�h7�1@�����RN��ݑ
�<�ŵ��Y�W�f+���j��k�s�JO#&�.m� �fl�G���G
&�1dN���m�s�:�t��8k'��I��=LU��%꽘(�u��%Epp�)���Q�F�4�	��95�:��H��@�#Y������Z^�ߒ,�����l̔sNt�1����9-�лr��[��N��w*�U�gZ�;c�}�uw���a���)b���	ӣ�vt�jX�z�U���c�M�����sos������P���!���(ʹ��`\J��hF,z�p���s�6h�],�D�ӊ�W��6Z�>3�IM�B`�ԯfk��@�Z���&w�Ϥ7�������x��?`��OaF�u4�Y�ߥ�'~�o�F���J?.�w�Ĳ*���D�W�e��� e! �mL���%�3Y	FC���b3�&5ٿ6�5��@���k���r�.NKМ-�C���cyu�:� �u����OE��8£`�ǀ~e\�ץ3�U��pw�l��? y�`I����D_��5����C��[>��cS���Ԕ�*�3�hy\���3�D�$c!3�����<mғ���h�)m�F
��W�Ц~�Z��*��+�7�ұW���M}z�t��w��:Y��Baü9,�j@�2�:�κ�=��̋��G��5��8�9E�����yycY��P�/�'<Q��U�Is�A�=� �0�8�4��h�U�s(ևz�}ua���kK��>@=e�+�+~�	�o��!�L��}��Ӟ� :�s~ho��&�����=B:��[,ӳB���?�;[�,���YA��28	5+��6�Sð��"�Ɓ���9�j�O���LF��j��&۴�+�
��{pz�坓�)k�b�V�������|03��>��ۀ|���g�7*G"��{$�� ��[rq�l�뎏� �lsr��<��Am��Q��ߑv!Cs�{6�n^�0��j�����T��Y�-���>U<J|�������{O�O�%���X�ш�S�M�l�:����!;�Ϥ���ȧl��e�@�<�ǜ�̧g�5��S
���,�ֆs������.�]5��^ ��{�}O�nx�w�o�eX���2p�6�����ZI�nge��wB:+5��"��fN.�����>�s�*T`q��.�����H���t^0����W��"qC���s��Q`�ֳ�,��1�G
- �%���:�b��ɥ"	������+�³\���_h�vQcL3�+|��UI&ց-�-�� ÆB�ԝ�0ɕ��wB^�H��n��I|P,��r����ά��?��+��Dp秠h�3�#ԛvMsL���[Э�[������T+���>~T�	�z�f��׶��9��=�5t��_�\�`�S�^ДYMq����o}���H@xQާ��v~��'��:��q�s�*f�*��R�������B<M2�áo�y�&�=��W5�q�:��J������[��}���@�;���yB��h�`��į%�����/5���0WXKk��&7��������8��pmah���^R�H!�M��5����&�O 	}R��ݙ#ղ�L��2�Z����b�p�6Plw��9HxO��'�h|k�ެШp�8�=�� �"��HZ �:���h��� �i(�@K�!x�K���R���&�&{��ơ�ˋw��av��o��?��ŠX��x� ��ju]��I��FU6}PK�B��
��Df�.l,�N�~�����`+����,񝖁�M���*՗��}_��c���4g���	�i�Z>�>4���|���+�j��%�����`=�y�p��-���i �K8&�R���4K�L��]6�I矣 D�<���H��t�����M�\��}�u?��j�r[j���NU��K{�E�'q	��@�����h��®�����?��p�8�����@�5셒� 	pH|���g�s
|7��Be�g����yj�2�C�a<�-�����/�;��@pn��p�=+5=
�!o'n��3$w�[uߓ�ݵ2��+��36yņ�G����]��WRaf�3����zs��&�<6���~�P����Y��O�˜��TC���h���D�Y3d�1gT�3#�@:�^�G���B��/3��3R�u��
֘�
���'oݍ$P:�kv,F�尪{�+�V�o�>#���3�7?U�	{�\O������?����~�=j0)PY%>�2>�.�iz`Z���ѽ�8�4k(PXC�oj2��)�xXj�^ot��Nvn�w1���D�{ǩ)����7!�Kϗ���ҘL�ͪ�[��6�?��L�zd�E{A(T��� ��w�B�nnI�){F�GO��m� �vM�����p���
u)3�6�3v�Kd�U��3��Ej� a0S	��/Ro<�rW�Z�P�
�㐕��^M�CICJ�k)Ͷ�7�ad����n֩Kۄ����۱�e�'��hFc�dbd,G�Ү�?��C>��� ~es���1D�$h[����/��*�d���������zk�v��F6B���:�w禿T}6��	E����3���ͧ�i�� B`N�THQ�a�D
��3g�Ŕ�ߝ��y��n�s��3�B_6�\.��9s�`D��2@׏��MS]	�G&��A@��m:6�6�I!x��ɮD���`���G�4�b'c7����R��pb�c��ѰB������ U�!���l�,�$��=��
���ʞ�S����k�WFA(���u���E�w$9��}��-&�����NF��H���B�Im�Ia�����]]`A9�t3�T|	�!a �v)�x�bP���Ox�o�/n��9��gݏ�Lu' ��%7��7^�:�����8��z��4�i��
U���f0��}B�>׬6�'��"'�������oGWM�z!=G]�nǆ��MT�q��0�VH`�__�eB'���`�$^���~�	�Κ-VV`�[Iy$�`��ܔ?����J�&�d�'��G��(���ז+��ӣ6�'τ7W�ɭ}�Qo���+�f��1*ʥKd��%aLA��sԴ9U���B!�Fh�J���v��4�amب O�"���zha��{�L�,}�l��u]����(�����p�֔�&�`�����ߟj*j�T�@�D�Xg|�����9,F~߀��tH܏X�@ ܶ�#�ֺv6?��z�EGv%�}|H�����b�SP�n�2��A��L��p�U��)X ���q�6��&������5�#��K�S�hJ�;ԺC|�Y�Q'[�ls(���z~Kwt������hM [�/�>�b�9��^��奄��[��a��q]��kmX	t 7;�5�Gμ��e6������BBO�;J |�-�x��fN�-�tP^�~K�j��<3�B[[����E�V~,yd	V�ŭUB4�P���^�|MêV*&�W7��V�{��j���/��v�o�0P��|������{�M����:GՇI��g3T����\�:&�ە[��y�[�����!JfTl8et�9f���'�ȅ����7�Y/5�g����@��J���(�@�&O���C��E���/�I'ɠ��`-��:YG-8�RȏM�����M���:�*�2��>�+E��$� 9k�|�4	��l�/P�����Q>= �������u�����mاQ��G�q�}��`�pd�p�qm"�^�I$��CA�kg]ӱU�H��Z㌊�9x7�yfƞOum�p��&?�A�c�D�R���V�'������I\��&��-����������.�}=f
���k�>e��k��n'a����p+k���6��I_}�� �Cݧ�A�=��P��L$���.aqp��Bu6�[�NvGɏ~��X�dV���/�י�P)}G�^��5~*z8����:f����RIv!�K�e�Bj�
�.�7ZvX��.��ԜG00 �� �- �(��<�#H�-l9
�S��N��A<���<K�i���
M�O+�k��3ԓ�\^�G$���-?�l�hZ���⪰���9y����zp�G���/`}AxDP�g�@ٜ�12�F�|�D1=�wf'9�[/w�<6mK�&�S*�6����{gp��Ur��	B ���ʉ�/� �"�~�m�7�B�9?'�|d������
�*��������z��L�Ѯ~,3��ث�ӗz�ߏ\���Z�<��Qk�Ρ�Q���ƍ��D�"n]Ŗ��M7b@b�t���3���w�ƫZ>`l�5v`�~���}��i���^�:Gp&�F_9&Ґ�yvŇ�$�z�o'd�.-��5P!!�O��	�ė���$����j��J_�S��s}DF"��/�K��妝������.����f���!�����F~����,t�x�T,�m��/]�<u�VMPe�,8�����T��$��Hg��WM�<^���}藱2�w�n�42�@W�%�݅��ԧ���ѧ�����=$D�����.�c�-��L�0M*W�'.G-C#�PJ2B��m����G�b�3[�[o4�}�ݏ�:%�+8���K�1b�q�rI!����8d�d/h�h��r � -w�{�/m.����R�[;�݌G��HW��>�K�	��%���g��ď
q����R`�obQ8��"�����O>p�t���!�k�j�@S<�\�̎�����4;}9k1Snj���=���a5����j1�yN�:��Lx/iW�<#n�BD1����=2�|���Ű�D7�:(;̼�|Ђ�8�?Z\���Qu�S�IV�qe���⎤^P�.@����G`�(w��3	?́:F\���<�"��-��i&�!�-�Q��Y-
n���P?0�#}�[��W����Cת��3�?��D��j��Ý�NN��i�X(���E�K�DE>���� ���>:ۭ��7J`��x��Թ�4�	'D�����Cͺmy���zԖ�Ԅd�g�t�.B��gi��ˁ� S��~�^I�b�!q����v�H��w"���57��&v2��5?����#�8�]e���e��3x%M)��80p��Y��r��K-���v|��.E3\'��h�gj��'#l��F�'��b���O��9�\a��B~[�/1҄4�&*n�F{'~z�E3�5���Z��ٌ���,qƱ)H*�3�rҒ=�"�p���ڨF�����_g1��?�p�3CX�_�c{�8,�к����m�.t�j��`5�N�j/O-~��S�(�LzRdֳ�ޘ`��N��+���a�#��w�t����X9�������������T*Wh��;�$*9n�Pq8D�ϒm�lG�( ����R�����o�i^�ba�M�wt��)�r��$��j0"u����� {S��\w�Lt�_��1�geBݞ��Ө�2��@D�7��kWFP�zKB3׃�@�ws�g��5)��0����H����߀�����7�K�M��e;�r}�h�L��Ve��{M"�~�d���%d`���tMѰ�嵬�Dy������[�L(q۩(�{��_�;^K�#��Y.h�a�
�E�������4Ȗ�.��xX;d�#(Sc����^�0�!yK�c���z�kB��~���n`�x#�A��'����.U��C��H���Q�}���!2�,1_��{N��D�������X�q����1�5���`?�QK��n:��(��V0����/ ?yQ�'��F�X7�m�'�~<Da�Nq&���Q��چ�������A~��P��� ��<���sV5F{uB�.�s�N�'�c��r�DO�/�,/94V�T�=`��OW^����g��둰�{T���"�@˒�[Y��q0tf�DPL]�Jg�D����g�5�y��.��Lg��IM�܍��,Z
 =����[�B��Z���m�����
�������/�Mm\�h>�ۍ�#��h��}q++~����X��>m�=&t�aZ4�`:��q|���~�r�n�
�d���}��O���1���K& ���}�#E��U�b��jh��̧��s����7�5�/騂�ʾ�2V�i��"�٪\�/�W�,0�[��L�CwT%�Y��W��<��8G��},�,��^�q�z��.�z�ȭf�:��*�|���#��#�-v���l���k�䢬,a���G�_!k��Y�P����`(k(��}������E�)� 0���B����߹�B�ڴ����ò$����D���ʫ.�i&�Dh!ηK��I_��64�d�#WYM�c����� ����q	�f�R�{�uo9R��Q�,A��MP1�4�Z��o�!����,�aăS�(P��������LO�Eq&w@�1�n���ɥv�Ɓ�B�@dk��?!vqx�(�rq:�J���˝h�f�y�xXp��y�IQ��#흱���X����Ь"+��<s9��-��
�ذ<;�o3���1��=�X�=��xJ��?!#�xt�-9f�"��z��6����&�w'ەJ�3ݠ����v#4G�����g�|G#��)_dat��z9�qnP��˳r�T� (�c�
A�ꟑ;��޿?Q�D����8�BZZ9�*�h�ĥM��*�6�6�F+*M�t}1&a�V#Q�m��Ξ�Ys՜���v!^��'d\�m\�"�ıΞױ��9�5^�D��
>u���~PY��V}�f=�c�Y���Ic�~I��}���H�2HI�w�ԙeKj��D��u��,����I�ѭ�#�bmD����4.=������d��=-��4נ>xK�����4���" �`�x��[ĨFQ�:H�'ŝ��c��0��|T�I�ٺ�+��Ƭ�@��e����p�8�{�ue����*-�,�V����}��J�r�%���78{r����5��8�=Nj!��x�]�]F�����g��׸���m��[���'7���+-���s�bE�|h�����RF�d��_q�����-�sԥ��p��\����k���<�ɖ�����>�ܪd�w���6�f3�_��-\�x�Rm��»���l{A]M��tP�'qe�:����`��UX���{�d'�z	��;a������j�2�Uxx�s�t����E�R2Iz�r{'��i��~/�tS�>� }6��2�XS}�cQc����\��L��MgTNo�C�]F��X�H�R�6��k�l�c���qճ-[?�ΐBe�����JΙ�8�ӫ@B�M���_�>B�T��nA��p��&��'�J'
*���ߡ8�r����T�!-��셗� ��T]��7H��lz���M������8���˞r�p?�C���jE 	-q���?���Y�1�*H���u]=�b)$!�IZo����.C��\�F�����=����'Y5��;��X'�y"X�/Y:`�*�V�n�$P=��*��܍��xVj-�%�~������������.��KP	UA��$އ��`��Ơ��ay�oL��Z�:��β1�j���1$G]�r�쮳���T�"���l�����
�
"���(�����X�/O
�iP�q�k}�	.1����5gC���f�X/��.s�F(َ����ߣ��c~���8�a�$��H��~�H2�{_���On}��K��|�Z�}B� .N�k��,XO{L��M���W��O�k��N�����"��I��א��[�Q���R��$6_���/}������HR�8���p���:ȍ��?y�ui=do�^F�1�!���ʀ�KZ�?z�bx� �L���.S�QV�+��.,�\�yj���*�q1O��j�G]����Tc+0�]"{K�à�6�ZpTWQ�ۦ�{\��X~���aS��"��=����|/6�`�_0��HN���	���;�pr�M
xW3�����ZS{Th�������QM�_�O!#��@G�DRs��M��f��bY2���:W���P��.�#b ;u9]X}����$����������Tx�/�aEܡ�+�1uM�*�ɳP��B1�!�8AV�<ND�l��U�&"�-�4�%�A�=��N�#��%{��&Ե�98Q�RP�[�P+�S��������H!xG�H|��ښ��^~z2� ����Tq�|�T���p�R�z��G�Mk-��SM|y�,^�����I���b�r	���'Ns&��YWQ��1���<����MM�,�-L/�
&C@h�h���@����Ã��?ϒٟVrq�}uae,��[
��_v�����&˼E���a�L$t��x�z��U�S*E$�k�srwDqg!�Ǥ�Ϸ"���;��ש��j����+(�>����q;_LT�I!ծ�� ���T��1��^����L�e,��M>N��!���E�!�]U�EQ<��[��	%C-�U*�%�9���]�>��c@:���Hd�˾0'�o����fx?3��TY��N/pޭ�|;ڙ�]!�����M�B���	*�0�׋_�.�����x�Yh+[_�!wwKF����lG�&�B�?aJ|��ovp�k�ĕN:��|Sl��Y��(�?Y��=6!z��Q�� �kL���#}�ŀ J�� yT#��n��E��(�1?����U��Gٌq����=)z�ˇ�;z�t,=�ɛƻ|p(�:��<�� ����y�>�$C	P����S�=��ˏ�Q�dx�G$�+j3��'&�#[+�K
5�c�R�����"�UF�uY k�濹&�C����(̟�H�(���[0��2���N��!ȘH_%k�M�d���͡c���o�!�&�:O�UE����P�>�߂��U�ilz��I�r1�� J�wCe0�wlw/���N" {f��x�#�(�ʈ���6���^�Z�Kw�'���4�����D��PG'�tS@��k���N90��EvM���F ��L�lIM��*�/2"ǵ�� ����a�f�bnf�ks��Z�k�ڤ/Bˀ��t<�N$<��&��[�2~%XV��bO���߽�����?���⭕+��.^���[�8>�R%��;X�!��QrcU��Q)�P��}I�mB�n55So?�+�Q^!���v���-�/}L\O)�g�o>U"35�n�c.m<@������hXYr.p��������l�Ux��8P7>�A�O��J�A+���Q&э؉l�Wn}F"�é�ѫ���a�m���U�Ye��~�ىB_(�pyծ�����n������mZƺ���j\D�g�r����&��gB����@C��l�>Χ��@�cg�+Ҧ'�O�?\���w��}��-(9���3z����5�Tt0��Vk,���w�y��'�A:�XW'��/��P��	7u����=��#b����x>|QwBb�R�c7t{]��N�8�}xܝ�w�����E|�x�H��6q7Oe���	��C��� ʢʝ�?����HJV[�+$��:X���4|{�Y�[���B�w�s�Ϗ�ϳ��1:"�� �.d�1�5�6��Es��FY�&���C�e��{^��\.���Imq����ݧ��O�q1q2�#��Wu)�!��U�+يQ��P�[�.���7]֡�Y�ť?�8��_R(�s/��zܛn��c�f9
�_�����97����B�F\ Xq2�T0،�ٳ�[Ș������׊q�!(��i�Q@_)/��8�([<H�n�FB�_m|#QN����ѝ9�p������d��V�w��}����5�,�e�ޓ3��P0Z#&��e�F��T��������y4�l5ܝ�V�b�27]��v��c~��*�)��Y�G��v.ޗ�N�������e���^�u��ܮj��/}c�(0������)�)��?S��=u�j#�C��F2|H�4v�d�<\�9W�j�[ޫ�ђ+��?J�/u���\��;Z����]�z�����ק��>��#���W��?� a{s�/��A��|��24���$m?m*����b5�d��D���spa\�� �mZ�˗g��Sj&->r���3Y]��
r4C��da�v0E����k��=���-�$윑0F �V�t����G��z'[ϛ����b�m��44 ��.ɛ��\��8qه���}����<�Q�Rt��Y����i+����6��b���M+�?�V���P?KHm����*(w�Yc${�S��/�k�� ߊ�\�q��q�˜�kH����m�@|L���V t�J��>*gMyi�Z{�%��(��2FGw�q�v�|F��+�?WpS��?��UJ	)�*xZ�?7�dZ��'�r)�v�A�p� GB鿗�p�R�}��Ȟ��o����hC0$o���g#;_�u�'o�ۉD#1�WN�& i������[����v�Xp/��t%Y��kXO�
r�
�E�D�E{Yn
Lw�R>�\��d�w
ɶ�2')�mZ篧�C`%:n5꧓�TWg!��C]��̞1��8{�ۆ�C�Hɹ�� d�[G��F��M��q8�_��Iп��k�r����?3�?���wTqn&��5qKӤk��,@<��x�sP '/q��qX�"�'d�j�3��}�&q�_"��S�j�X�0����ͽHT˖������N����`� 8�9@pʬ؉TD!NK=ƌLr���ʙ!h1�i!@��@�ۨ��L6=q��u�������'�"�p$%ϊ���	>b��[v������PپX-`��E�0�VF�b��Qk2���"��+r/�,�O����J�/��t8hd_Z���= ?�T�\Ԫ�C�߸?Q��߭��
������'����w1���h�:�I�r�ȫ��q�inñ&��ڝ�1�3�.�1��O���PKg<9�������vVlC� �4Bs�cHߛ����8*ŻN8�>�\�	�c����5�e`fϢä[��	-%�d%�B�hD��VeHȇ���bdM��5��/J�R��|ϣݽGVa?��c���.�R����g��"%�����鐙�#�hh�����k���_Q��X̶=��9K�9�9�c��%�	����a�VO��_9^^��6��|Dj���!�E�tjOxL�������a];.��h���B��Y*"&{�ۼ��~~���ߊ�?y�3	u���aHaG�P���=+�įWn�o&�M��Ë3!�7,9N���㨥�w�/u�N���Â�����I��2�-��.f��Wk���b���$(©�� c���C&/*"Zh	h��!֕�lGbp�vE~�_�����2��LY~dD�E���^A^�JD�����˹�kN���\Ck���c��FbbBo �ֵϋ/�3�;�$�=R�_%)�p���~J,Hm�T��.)�h��ӗ�P��j�,j�j�Z�1�\r���<�n?mL�MH�r�[:��&A��r&���\�
`���q\�/�YsXh���_ $��"�?�N��P�/V�xM��YpA��DCכ���i���a���*7�)���F����7�|c[���p�BxR��~U�&��'t��6��У	B�F�DC��&3ȇ�ңTl�p��'���E��?��t{%3�r����{�y}�zx0��?�c�˽6���_�� �����gT���rQu���@G�_�ϵ�=�/3=`+_�6B�l�60�t8iT�w
Y9l�B�J�
ˢ�
� t��T�)yZ<�:�j�1�No���W�4�oI	c#8�
tVȣ�˴�	��e}YziP�8;�r^����2_ը����m\�1�F�N��IXC]�B���m��}���q7�T��'o�����S��r/҂ed&`������4�%��ňN��Z��|��P���7��.b��(�����������0�Rc�wh A�۲�-���)ɮ�Q��x ��l�������b����ݛ
;��x� y	m�ٝV���	BH��Mh��I�.چq�ta#=������d�|��e��\�o���i��J��t�]K.����x't�8�T3��[�>��m�~#�L�����ү0�j؁;|J������d�Wr���?Mht�M4I�lt��A�c�˥+�um�=>�?G��陔(�{dW��@M�K��*���A�,.�zgHP����l�E_���oB�v�~<����:)����<�=x(�p�W���W���e�?@�A�E�U9 �j�#I����	�U��WX'���w3^�$�`�/Y�A�iC%�����m�3������j\a�I��v xvf���(�ޝXPՈh�2K�����ؔٽ$�y�K��!!�:��?�Ӆ�XMg�Y��*W��O�ia ��pyk߫ᅊ�����5��9|+�:�˛��G �X�A��"���:��.a�G�2��gᨳ6�E#6��/�}
�O��l�M'O�@j�b�ф4M��@ vfD�_��M|1��<!�x���o5��ңɎ�(�	�&#׭������[�X��8+a��PSB9.��1��-���qƗ�5�i�}�LyKВ
��9�q���SJ�Yz�+�P�K�0A��(^}��6�QY�܊*cdS�G��K
��)64�Z+s(���se��=��_�|������^1�-_0��	��r��yjY��l�.	��W��_��N�(���`��,*�Up��㬙��F��i����S5LY���~�k-����Wu�R6/;2�^8�|n�'!��bݘ�`��X^��\pX�ш�{K@:v��[
^g���M���)&+��⩶Â<yI@��TлN~,�J���r`�B�g������|�&E�S��l�!`^L3<%lCֹ�\Y8o~���r��#	�ҋg3bJ������_e����;�SGag$ϡ'���C�|���h�F�)ĝ�75c�[�����O��^�涠�1��4��D��~@a����"ы�♲�>J{����r�[�X�/pUBb������*N����F6'f��vm-oD�$)aEz̝h"A9T{_������~0����cv�j����_��d���9Z=~�rO�<����w�u����c������%r�Py/
�XN�ƣ�g�] �2�/�]C�)J�B��"v�OT��Ņ���"q�H�Y��u��T��{C,S���ө����:�sDP�.ci�����������]��1[�ޓ&�W7�	���@F��;�kgY�g?x]�k�"�^v��q����d,�sG�`�uJy�����5а=��e�R�s�� �ѻ�Db7~G�5�
{D������s�p��D�Y<�JZ0R�h����G��ڱ�y��Gz/��P9_�+�%�yw�3_�^��D���t9Y���a�8�G�4�5Z�����/z�}%�!E]rPтj߼��t�u��lBT�͙/�"~y���Qg�-
ľ)�i%�5����͡)*�42��Xx4�z� �؄�+	���iu0�� \~S��\�LA��7��7I�u4����ӛȕNt?|�� <(��	#!o��,~o�e#Rvߓ�5a���i��F�p��L�x[~��j�0sK������ȓgy2���E��W	�
�՞v�O
��c}ņ���x�d���6�̳M���T�1�;��Ǟ,�>~k>Ѥ�Bf_ᧁ�dq7r�+I=�0r�6�'�(��g�rTo��T�q����7W'E��]t=��2Z��|f���f�E�}0>�,Ց�>+�'�����QNʏ�p��*J��N�zX���(���Z���y��d���u)T�t�_��OT�ūY�����'��˸���� �l�_�����K9���d���]}twxσ�G�#sv��E%Û���%'>=��"C����G��9����5�Q%!�o�h���w^ݿ�� ��[x�5�XH�d?��̓�n��w��ƅ����[�g%~d��胡���:�筙L�������ʣf�=�i��P�;�:���w~����rq��t?<��z�Q���	��@֧#��-�f����`�X�*��E6~�����(�6����9q��-�0l�]]� ���J��������bb�� !��濔 m��`�����0s�ֿ�Q��EY_t��aXŮeEW�\�Ӭ7G�P+�|u���A��S$t����$hDk-�c�9zڱ��2ط����'��[4�ܬ��<�a0��"��]f��:�\`9&�wpNh����T��\Y�c����D��;FHԡ��@�؃��*��IZn���d枔%���F<6�3U�AuL)l�� :
�F6���]v~���Bt��"��Љ{�	�s��Np��*tn*:#c5��u�h�Bb���u
�5呖G5b�����&����t���A��R(�S؀7�������YVN�Xў�벘"�@Z��	��������V^��QD�bg�R`��T����è���N��s�C�������+W�)Vw<	|��s�D&�XGl7�v�Y��N�y.��ІK�~tV��i�>eK��P�Ƣ��G�]��$���&�E���5>��	dD;���Qfc��oă�lפ������| �4���]W���0������4�c��R�A���}Q�a�*t���B�ܲ����]�+����`̳;��+F1*��%�����ξ�������uh�]�{�W2������S:�̠Fi�BV'l�6��R��Z�H<`d�S6�;�����k�?m/5�R��D̿�Sޞy"�!�\Q�_�ǜ93j���4C��n����vqb ؅���|�[�U����#�2~�.�� �ˁ�SI���Ma���f�$`��)\�"��l���`X�<P�?��^���.���e�C�]}�y[#���>H���7�x�����qF�F�*pg���M�k�x�<_�k�2n4��%�%$jc��
�+	��C���*^om�h�EI�y	Vѻ9Z[x�W���}�6l��*�68�P��g�Y�!�!���	��Xve�%�	�BU| �ǭ�lx"��t��{Ka �S���{%��n*�

P�(,�8��G<\�LX���t
&�J�p��"��77�q�@sg��gF|��t��􏣙e��c<y�pH��dH��]^5�'��mÎ�<%o�p�H��4r�7m�Ǧ{�n�w*a¥PQ9k�7��l����J�GLT 
����M	�mq��&����@��Ys�Rݳ��{5��V���#�v�ڧ^I��FPK�ڜ��I��E�α�aK�7����W �����2fT��$*���?�y��5�h*f�}�R����@f�"1`�vۺ�\ ���:�M3�@ס�]��D�"~Z��#�̕mY��7����ù�[�/ �"���ם�*d"��ӗ�Ӑ���@��9��j��k �"�������q�}�` �t< �'���x[�j�G�bLˬ�;o.�}�'~}}�@�:�)b�^Ê�W�[݃�w��s��,���ޮ�"��>U���Ϛ��d0R���^-�.��"���蒵�<�:8^��?��
�:��v��C�o�5��0s	vW�H)ra"[T����y����:U��?�&m��b}[g�]8�v,ԯ��\!�����aA�QJ1u�q��5�q�[�k�6��D��r�|�����/�gGv�֡��z�usC��z,�t���)߻Pܢ�|u���?\��z�OK{m"`�?2�A��ƹ�ǁ�Lk	����f2�R���5��i1���In,�*-�Y������3S��\�K���賊j/c��;b�W��1�l�%"4����t�🿢�F�V���X���r�ₜ�)M�BЌҍ�8$�!�B��K��/��/kϔs�-�7&M^�����bV&Yi��=!#[��-�g�fM���O���� �f5$��*�������4Թm��Ɂ��AZn��o�l�|�֢4`���R��K� �H!g(��O�@(��L��KN=�����3f�Mi��E���)�d�e�esZo��R���.�J&:��a$R�1���i�,� @��5qE/7f�y�� 5c<s��LFZ\h�^�Z��,��$Ɩ(����TXv�ʜm�����r�]���8�9|ƀ�GKߐ���y2,r�t�5p����w�Z�2N��|�p���U�H�Y�a�T!�Pԏ�ܤ�;���"g��3i��5#[�գ@+�����٦�Aχ��E��������iT��FD�A���Ot�)SL)H>���u�]��X�^���� =�9�e�����z�ݏ�Z���Tʺ��������P2O�z���'����4MK�p<��Tq0�����*dm���z �?zK�S5��a<h;'��Rd\���u�;�K���n���:,ێ�=��BEi�+H�Tw�Ŭ�ɾ��e���hc��)\q��Nd���
d�\3� t���'3��,���:ɴ�+��ȣ4wG��0 �d�!L��|�wE��4"-�|k�;W�<�.�^�c]pF��<!Z�/~(��k[�2�٨��ڀ#���nt/�K[�P$D�O���
�0!!���Qm�����p�>#���Z|��Q���x�퍮@��� m�G L,,˖w�7��b�����xҾU���};6b��U�!�p~	}g`���7lw7��ڮ��\��=�!��*�yƚ�B��]X�yF��u!䱚�"O��'�
�	MR�{�$�&�(��}�����Q8:#����$��l2�jz�|��;Z�qv�lwy$X�{���`�	�HgQ1���+��`oE��el�e,�nj�LoI�
$�rw)0�U���b�1��[	t���șRB�~
G7_��9���W�6klV�T�|�n�_�S���Y�mc�!�E�.�:DrMU�ݠ�:oq�|R �A�g�Q��h$J��_�ۙ��� �����#y}�+j~N|c�����},8e7�kO�^F��Zv�t7y� {�7/���l�Xe�������fP�eX�}�]<���H���J�=��Z�]�����01�2�����1�p����u�D~Ѳ�2�rOQ����'�I>9X��K�i�7p��,�|IP�:�CwxQ��}�i7�g�<+H2o��ϳE�E,ʺ�7eD��F����-ѩOM��%��l��R��[�0�6�MDX��r۬���
�tZ4^݊��4D�C� �����r(�P7���_��}�xmf$Ȭ���*g�{+mQ'�'B  Xa���woK;��W�V�(_�Y칹�L`[\��|yT�H�I7��%gzbí�]k�	�Z1���t��0^�V�M�����tm�9C6?1Z�8�ŌE�6��i�w9�G�ޏ�Ɖk���x-\�*�C��;Fg�`�1�G�@�%�A����N-�t�7e]�.׃k�v$��;�-F�-�5�%e ���3�p�ˈ��������6�F���,���>`qSm��|�ƿ�=+z�'���PQ�y���^�d�+�bmd�z�{��q�<ń�����8:�P�6�{	��֫���ơ슏\��k�A���?��D'��3���޺�۪��֥�?�n����βvA���̑$�)��e|˄ٜP�v���$��l�l/z��@�R�Y�wIH^K^���� � ����HA7�����p�@ ~�b�~T� � H��uf�_�!����V0��BS��E���O�,)�jR��YH��7 x
��	��P���\SL$��?�5�I�4������aDP�N�"S	��������Z*�x������$�M/�[]V���xv��� �3)<02d�� �##�"P�Q�p���S&�3ߜ��o#M�R"�m{7���ؙM��é�t���>�������:��5��?\�s'�wE�8����� �6 W
�iON^u�/t9���Z��=(y��A>0�[)�$§)�����%6TX�Wڏ<��1k
�y8k5���pb�� �Fh�Č�I���?��)=nuPD�غPm7�1!�V��~��]J����N����X�GD�1#�a��.-���V��+����F3�E�T��vU(S�jE��0��5�2KjJڪLw�!ֹ? �Z��ډFsM���0Ŀ�$!���{`���>Q*IV���{V�<����K�do��Yr�V�����]�W:ԛ���	��Qb#�v�`�z�2�a�Z�<1��aZއ�V�V���q�qQAAJ�7�k��ʋ��k���c�L�ي��֪���E�v18�8�n%yT)Q]ܴg�"�^���ǘ����i����~f2	dN�� )H<�8�P�J�ގGH�>��(U�wl"�t5k����<��Nc�/��V��	���.�:P����2��Vo|Q!%�yx��D"f��xa�i���;�x��s��2�DƘ-�;�0���_�S��D��X��|B����O�Y��+�4/,��:��AY�#< �����z��~�9 �#{8�N��XV9�& �]��:�k���ل�.���efP���*> E(Nf*W�i��>rp�@�G����V���+��'+� ����Z�H�A�OtX<�|R`X�+�Sdoi���vc� ���-`��@���E}�O��}S\	BU��:?�I_Yx��:Y���`u5P$�i���n�`$��5��\�sU ��啖�+��K(	���L�8G�:	Ώ؜;�6�14Io$��ȼ�F�p�u�v��T.�����_���'�Poʞ@��51��73�i�RH��6T��)̌z�g�Ǯ������K'}R�1s�O4�Bb��I��\<i�<�����R�h+ZsX�h�Ry�y����l� |��c�1��.&C���MBz�#�ղ�{�6.ui�Z����q�:QaOd4�Sucu�-��lz�/��.�1B��+�W�p�H����ӹ�ۡ�a����G@�3���T-��R>�� /�L�+r����Q�v$%��9�7�Q��=.1�)$|pV|�R-)�Ha~K؆�����c�:M��P���@df�#�(�|�+�Q�lK��ߩ�m�Y�;�7K�Zr~��m�=���,�9�����[�O�5z6����S����3/f���23<�Ar⵼9��Pl p��r%"g�����i��H|�J�U�nl�h��v�
��S��]@��6���2�x�'��V}Þ)P�,�x�g�8t��!2��[�4
��.��Z7�|XPO�����kӠ�]�
X<U���]����c����j�o	��RV�U��;���nX߀h��!l1𒮛�˵J���9�\4G(fI$��&w�RP�6*q�5}�˲^���h���쑪�ǜ=�~�ab�;��-�k�2,�7�e
H�4�_�6��>?�w��7�
�X�č�g7!�,�g���s�L���`p&]���p�exƜ��]|�I��l���!bb`M���5!����bP�\il���%�
���M�N����}���
;R����j�Ns����`�>g��1�؀@_�73|����6o���{)��<���o��4i!�]OȜ�[��]���tl�����l>̦����H�h 6#�
�>�N�l)i��x3�T�"�Zƅ3T
K|��زY�ۀ"�+�d�=�!/��%�;��U������*`.Gi
�L�V}Ξe���wz���	�3[tri�( ^�}=�t��
I��E�X���\t>Y�A(]�;���,��-$ť�f�,�Z{�*��b,rm�w�]UIl�wIw�y�6�� ��GX{<J�
'_^G"�n��IA�B���Ŭ��(M��2��Ȫ��uO*u�)��),�����y�rQ8b�B�*Zeg�}6c��.-$����֧�`g׸���%<��FǇ�[I���t�dL�*j�B��GykW�\n��o@G|3~]�K�VL����|�MbnM��MXa�S:�M���0�A�:�3��!�Y.���jU�/>�_�k�늶�iğ�	���rq7����v�be-/�tnbCP�2p��?7�D������w?��B6�׎�t�eҷ���i�<o.�O�36���MbNg0}ѱ
�&�gU��pO��z��9wf����"{�O���� �/�F�1.�-�4��&d������g]�d��������c�ޭ%j�,>�,C�������H?.�X��w����Ʈ���l1�FfA���9��N�:�)�@�9Q'��4tp�s�ʘf(
˥q��_�TxA+c)����%	�H_�	�����,��G�p�%pi�x7��Z`-��^	������/�:����{�8�yy�@ƶ� ��9�����V�o��B���WBL�mp��9���
H����Y�ێw��M'�[��0�.vy[����.Z헗�[�t�O�5JE�a�c��t���W�3���2�ȥ-%�¡i�g�ϫ��Sd��
��l��V�{;u��̗��>��!ю�8O�3�d�g����t��'���Iuȭ������Ʈ����ZS踑�B��M�2ύ�����>y]b:遙�Щ�p���LG�t݄��m�R�; ��w&�p}&m`��{�[��A�D��e�Cx�Ņj$��H��ҁޭ�)�U�]ïX�HU�qd�}�V�d�֮)�Uؑ)8��I!�Ve�{Y�T�����?�)�d3	���\�=�E��9߭Z�z��::`��]�n�6ܗT�&ky{�o���4���`!�ZJd�ʑ�NS)�v�?<>,]�)�g�K�v�Ũ+�hG[���q{(� ���17�,��&�WjL��/��<%�%�<��4���),��]� agFa_�Bd��D��E�C{RRvdZ�7�ؤՔ��ĝ�⒌�C���s`�(�Ú�b�a���l�.���F�����f%1�D#gm� �mJw�
��#PtY��j�@�jm @��砑�3J/g_6Z�w!א�=�~�/��9K�z=_)ϥ����M��1�&f��;(��,��vԔ¬�m��=�lբ�S�F�?�=
 o�ɛw[	���K��
`K0�U9y�����o��(��4�󜬐���&����� ��M���	޿H>g�L���~ƿݹ�|�B"O?y���x�Kt{��7���3.�����A��-hY�hz������ZՓ��9и���z�/��88%%S�	�;<�-���.�8�-x�1Ia�����|RNwۖ�u�B"�Y;h����L��"��;�f�ZaJ���M+^��Ď�w���O�rl뵧�z��0�5���$�� wX�c�:n Cף�b��f+@ X:��  Î&�O�V��&żNi�s
n�t�iF���.�i�C'e�È>,��j���Xpx���}�L4.Ǳ�ũ%I2=�2��pal��8o�@5�z��NS��3��E*�Ax/��=ˣ�d��8G�3�C5��K�����	h�8���:���]��wQhW$ċw�7����G5���ʁ���n�!�rT�>[��E*�����=^?���}.q�.��e��O��B˖m�_[�!)!o�+�,K8H	J5��pJ�:���KR����6k))|�������g�T�@�>�+Y$�c��aq|Zb�s���=)t��	��|�l��'R9y��	U�w�/6+�ƹ���ǚ�r��=�;���Ȗk�f[�<b7�[��*��՛������y�H�4A�q/��X�,bS}y� gַ�/�L��xTm|��ue��R��w�A�߸�x�� �XwP��|���=E�&����r�.L��E�Ym���P����9 �gC�B�'���8�L)�,�[D�@1U�+�
�EH������1�'�N7��"b쇳��!@��y��)
-	荖el֔���F����{�~��@D/8�- �;�
��gH�iI@�@f��&���}n�ƞ����C|q0}�D]�&� p�Vp�������̬܏z4Z���Y��4/U6�`�7p���<PilJˬG���E�7q �C��F�SHjU�g扮}���֕ux4��	�C"����.�)��d�!�)�����A��d���pCG�[��Z�0�٦�c���a�;�݀G�D��g8�A`_9��2�'���$��]v䕅�Y����ow�7Zz�O�	6�kS{�HU�4�RX�ğ@��G�FD"�����̅,=п��'^͢�����D�vi N�'w�ȴ�kzc�*��~RoMS���z�W��p[;�fL�DN��D]�Ǌ=ݲ ����5�b(��7ल���/~O�Ti�"!����LQ�r���7ZE�j&S����\y���	:�=���A�y�R�M��, B�S�K�`���Dԁ�%���d��c�:3�5�P��>��7�����j�x��`�ݡCٽzϨ'F5d��k۬�,�Wz�;�YwA�/�,lV�{b��^hM��,�X�$��\NH}}nCHEٻ���"�?
�11��e���Jk���Y���R�z��5>��y�*䏜4r�����X��s�Qs0��k�T��!��BS�A�1����`F������8_��X
8�Ν"c���3�7{X���	�K�|��@HӁ^J,zmG����XTj=����}*
@�����4�KK������`y�b	m���93D�o�LT�������J+��Η�-�i7���""B�eu A�L,"�;؇�k��DBq� h��9�3���6���=��Ͱ��G Z����U�g�;�}n�����}ǻ�*;r��EV���F0��cF���0ԋ����@xV�&A�V7��nw�}�Pq�q�0�1�b�WO�}Y�P�1I%S&�@���J��g�EK�na4պ���nڽʟ@��G��v����Tz#,��SY���v��T��Aל��p�4���1�{X���F=�w=���rJ��� 2Af�>ʍ���2'�n�<����{5򖷁~HcC��U��5_T�O��L=M��s�ÜBz17k�~�3y��4<���NsZZAt�jLRa��+W_I�΂SR�r(6]t��U;!j9����K��>�j,� [r;����՝�i�%d�V�����1C����[�f���H"|���ִ��hl7��'�^�'��$f�؃�g�*����H�,�Ⱦw2K�~��h�a⚎BY�� ۝-�[�����M��B$�f�N�UL"n��5�!*d*G�i�;G�Id4����X������$�[���R��ꞤYpއ����-_{������8}�4Ts������MS�R �P ��ᖣH���w��||\���NA�b�Mz rY�tA�a潷����s���8P�V*�����.����ﻶU��z���ӡǠ00
g���=�YA���㲄ƫ'��GuEGw�¥���Ж�|t$���1�G����n!%
��Q�|���jpF3?:~���m�Pu�X��Ȫg���wԺ��Y�+td���
���R����o�s��FL l�bV��Ңo,1��X�v*�r�_�8_���y����}���z� $�5A���7��%
������{&m`��)�UG=�(a�b�H ~,���f�g���K�_��6�3��HcK�M�(6��1JiQ�멝6���j~�Ǚ9������.�B����[bi]�a���b%^�u�����^���{~���2��]w5\^tibفk����R�a/:ȸf�UcO���Ř�@��R���u���w���: u(.�,��.ϝh�C�H�G�?��\j�bG:ʕ.,��rGg�fib�>Kbm!�b�������4�J�λt�I
��)����7z���=�߸W[3����Q_��U�F�"=Ŕq��2�xu_L��������n�~ ��3iW����'�7��;���FU��N����C�"���{I���e6�E�v�"���J�Y�����S>#ϑ,�1�qE[�31��v�#�m��7���)�|�D ������V��� \���u1G�pbY΋�	m���8�}�s�i'���[��c��N��rF{������d�����#�0��ĵnJ�o�Z�$�P�����Վ{��/�y5�[���a!k�3b\[���ȓ���@{sS�T������¥���.C&����7&l���N�g�nvդw/�\�f��,]�t�¤�]�0��~�.9 ,
#��f�罄L��X@��R�W�o/̹������gj�)̄<��vI���ȃ^����8��ک,
��FC�ɘ�t���2�=�ɋa �`�\ ��R�����E�3H,l>�q��E��K�U9�i�L&N�e���n�ڑu���oP
r햵���N4B�C
�MV��"�4����e"�`�/|�sqVF^P|`E�&"LW����;yq�9�$9�:��Bv�ʭ��	 �
��۱�����˔JG=��xwG%�ʷ:�6� �=+�OT��"��0�#�E���kMQY_-��*�&��*Õ����|�t��9hpJ�A�O/�*g \�M	���r7�-��"OD|A?�Z?�ӊ�D�L���Uȇi�k�
8U��_�F�ƟCh_������I�v��dO����MݑP?�&��{���,`�^���S�)�Ӫ��P��sNlO�^��@�|/�dnLjQ�m�y3��P&�0�[��`eH8e-R���H�`1Kk�� <lF�R	%��
���h��Y�S�.y�ܡ�?>�����·��lv�G��)cK��E�VDOo�4a�͌�^ py@��VM�>��خLT�ǆRʑ: �W�S�}[T"�(B�V<2�%6�<������t�D�׌�
t$3��'�*`���u�)��*�<OX|�=���Ԗ`��៼�ܫ9ڙ��<~[K��.e�Q�Ƴ�΂W,�]f�-�V��$���o��a/�6#e�.���C�T˟��B2�m��9�oN�="��:4[���/�-���ϥ�*�q��B͛��r�ߒi�O$�>	a�]®��4F��Sy8�	1�F����ڂͪ�n>|�>�a��l��T���:�\pyF@��l|g��G�Rmx�� jk�Ǘ��w2��⺧s���[��nb�@�\�C�ʨt�6��qq~�5�ȅJ�. b�|�X%Y���;�S�I���11>�pG��%����B�x�}o=�7�`&]�\m꠹�G~��������CE���O��~���<�D��j!�L����b<�r�H�� �"��
9��(�+?9:��S9_T�4���O�Y�������נ݌I<Z�1�W�jm�����ѧW:���L��8�a�,eh�ŖqZ�z���'����ס�>����,vb�9��J�@��=�+ǿr��g��1�T�S�DN2*Q�7��p�<71O��K@nj�.D�qS
���Y��`�HN���C��'�W��uI��p�D�Hۄ�U�����0�<�3U>t15���.g*E�o�~^]f��k8�hBr�qAĬ�x�5�b��n�� �l��Q���?<Z]���〙@�˹y��s\^�N_2�0�C�V0O|�~��|2�6kldnF�I�I��U��-���@�k﵉ �^�y�LI}�
kl����*���^�.����z]A��/�O=XZrI�՟؎;_�	���+�@Q������:UN��C�a���N,���	c^���$���,T������F齧1%��ʹKU�?��@`�4�qI��|��c��Ұ&�mS�U@ww..ڛ�՘���f����t���xzO��a3�B)��`��c@C��ձGY�5��z�r{^��륩ii�6̒_�h5@�(��E�z��J�7 ���v#8s���g�ki�v��#`�����?k��<�,U�99��q���qC0�Yʂ-=�Pj�G҉w4TNȖ:�]���G��M�(kRC^{�v֨A�~�J�����C�f�h�,��B�@=V��J�$������^���V ��jd��!Y���E�>\D����Tб��aH�]s}��g_����.��v}c�}#n�u�=c��v����LN��N^����>���E����!/Ss��ư��Y*K�Vݣ���o�����;�k�wE�TPĘkX����t���FU�ًU6�(�m���҅l�[��x�N[TϞ뙟�2R�� �A��������H+&�,�/7����J�&@3�����^1r<����z0+�Ρ�1@|�>��[!*8�;�9�,��D�{��z%��?���H)�ء�D'�������%E��T�N��-��u�ᔮ��t��M�@���zR�rxm8�:U�[��8l� 8������`���<n�T�,P���a��wa���O�(�|8{F~5?ܻ��%�A����Kˢ%1��_ُ����Z±��!��!�6�	��"��IG	6n�J%��ރv9)�sv���^�[j�O�'O���D���ng�����K���A�����A��� !����!_��R`����h�ef�Kȷu�Y�t<��\���Q��֬�SF��	�ؠ�G@?y:�PY�Z�@=�hͩ	(�1	�r4*�F�&��,��v�
�����W}f�f�A�ۊ/K��:(�<40��Ү՞ۀ~J��,�ţӟg&�!�EZ���h�������3��eF���?T#m����a�EO=I��(�(���CA��]P�V�����1�% \��K�\�i$ut��i�M['7�,c�9F.�6��A����;K��r������\� �S&؂w?�˷�wg�<�di²T�����G�M��j�$PҘ/l�r:��A�L#��E�cH��.�۳U�7���Y&�wR;[�=��fEʾ�G�\#7�B�&�oT*����3��G݁�sS��n��!����88"�8�!hr��|���y�Ǜ^��^��g)�R�
X\r�[��%#ݿ0��ents2�I�Ӎ|.�Gݜ����,���
��l t���'���)� �p	`D	Vc�%�B����i��K؟
o�A���
n��B
��n0�q��d���_F	�G4L
�c�g��-�6~F�"�fZ=�W1C�=��΋��jdP޶��v��e�z����p�D���g��5U���>�&��3�Z��b��Q�쓿]C�M9!�ַKHT	�x�*]`Eq|�Q��7�G��'�S�7���|Ne�?DƁ����&D�33���Ugz�E��圼���6GY�s�d=Ԅ�����[f�
��h�=�_���o拫k��G�K2�s{H�s����a������3��w�V'�?���$����Ȓ� ����������,/�F/��,�[����ڡ ~s����\���!Ó���an}[p>`���rB��]�k	�H(d���^���i��mL�a��l���P^ֈ�ꂦdw�L��/�l�ވq8>9��	k%����Q��_�=y*g��L�ghM[35��Mv�`w��GN>�2�Ϡ�8d��|k8i	>�
��alh�v�
kL�#M���&F��P&vkja�d�$[a~\ Y���X\�n�;��68���ל�10.R�p�l�1K��� rOP8*s�,��|�#������?k��7?���G1GNn��)�YdU�^���/��d���Q��K��F�:`���aP(j��Y�9�_1�\`��λ�u�AO�Àb!g���@��{��&%��ˤ��	�َ0"L��⋎T�B��_�sP�!S���2� �BЀ7-�|�
����S,��M�הe,�OU�W��!�yE/��+H���A8��&�R��ʹ�x��9:��*٣t�����s������b��v �(U�����Np@{�:�O������~:�+C�.J� ]3����x�K�m�V�͖Y���/�%*���!jvP)�`*+u��Jq��<j�X_�^��*��M��]�U9O��s�$v@D���.w��eہ�ݯ�6فP�QZ�_۞�X��1э|My�M��rj����)yF+n�Bٕl
rP ���a���]���F��x0E�o����v���74�eB^��"V���ݻ�D���(6˭m����1X�j�uyÃ�.�^~����/�~�j�?`:{��hY��	?���r�ҒcS'��LX��@�pczNÖ� �wk�	�c��g���䤒q�39|k>���)�[u̇��W�MG�vz��p�S7��)���K6H�����Q�5`;��d�/Jl���D�We)3�>�?������ ����V>��4�[}&n;��.��i�ϗo����[��/���H�%�Q��a��^0�,㵳^��֏�"~���۲�$�0�D�e�9*��w����ܓ���\j�+�hy,@�ip
?��%vȢ�c�\�������f**N��p��S�����wM��W��Ȭ�A�	6������eWI4D2C۳�:+ZF�|Vе��`��S8�_�|ng��h8�M� +NӒ{�[jJ�����t�Q�;y��P���	׃4���j�e���4�n-���_�����5�eet��!G0��@/�2L�+�P��ϸ�LP6h�0�*ĩ�=0{�M��a��2E��N,zPSg����s?.Y}Xl�Ϗ6�-�@�-�u���P0Z��T�JE�/�{��oȠ�' ���f����ݐ���X�}�`�jί�5V-G[y�Q�uO�g��J1����~{j[���tp��Aw{�U�>���N�T
��W�mC�B�֤ޮX�����߻����J2�v�Z�'͆���|H�w��)�j�JO�t�<`͞Ӑ	�u�}7Y8��r���D��~��Ť���5/4$ġ^B-�����"�n����:�d�$��=��my�ৡ��"����n�&7v�n_@P۔|��o��i��Ρ�αc�݊M;����L����-V>���ZaKk��U}�dq+8�
�-���T�׾u3^� �i{�9�����N(B�y�WU���3��N >c��*cf��o����]�]HrTզ�}DzD`e�1� qprRLƾ�\�h��B^q;*�0Uª��t�$G��!��P��r9xސ)�9$�g��q�4��I����2X��<�ɱܤ;TN������Cb�>�a�8�@�e�DI�C�I��ʬi'�SQ�X�NM�\󧁆�#G��p<��w[A{m�
a���?<�i 0���%�ԓ~�LW��[{�<릆��5�b�!����R���2Z*<l1�A��褯Y_�>O��Ѫ�@���n"�%���<%V�Y�m����P!��a0���B��#?��Қ�>:� 
�%�!pyg�"�,��}�1����S�ǎ9�@:�L����~��ىQpA����\��j4�9�^Y��j�@(�T�aU���R��g�)���i��#ݮɒ�_����`G̚rgWk��]께�~wɁ�uu8���0pvP�5B :v���/*�����?���4͋��D
L�8c',�d�K���V�㐁mL�:���Ϋ.���m*]�Cj��d�Gk�@���8+���_��5���n�����ޡྪ�Z�/��L]����+w\jH������D�1���Z��nHuF��\�U=��bCz�6�@8:EI$���S|CJa%����@R��;�wy�7��B���}o9�rea#����� ؖ�Fe�ܟ�,�y$�u�5�a�I'| ���� ����4
*���/�������[��v�g�{zo�#<h���8d~$%E���k}�|��Ͳ���db�����.-����apdt�r�`������q����h��Ȃ�7���Q��j?64K�G���mý~�k�H�	��1�#_1��6��,3I�Cn)̳��ۍ#��m��h,���˅4���K&ۋP�Dt�U��q��E�|�B0Ć˿�^���Hw��k�9��$!Vm�ڷ�P�`�	Is~�r(�`%h\����m�)Q�JPZ��j����I1��4�]�%�E������{�0*�k�f�D�t�d�CsOP!�l�oY����Ơ���_�e����g��o�c��ӷB"�e��D�=y�n� eT��&9���D��8���b�Tb��8)v�xs
�~{`��#CU������A��,��M�u�+��\���#�, W��P��ڶ�?�t�k��Z���dYi�߲��s�¥C6���hŧY�8�������l�D��("�h��Oߤ�R����>�HYf�� �����&rO�fqy�@�a,ՍW���Bu����E�� q���1�b��X�+'Kȸ�f�����A��2��L8Gr���N�A��/6�h2~�Z0	m�3t}I6_8�6�.R�Z��U�\G���2��=&26�B�d�7��KR�B��xtc�>|*=�{`%���4�������.x�Do���aPq��e�}����ب��mu����x2؈��}m��%Z�u����h]Q�[K�L��\V���c�l/��>��b�����n1NxPþ��T)_���P�܂�!���(�t8^x�r�'C��{om��k�����sc�H�eB��}�D B��*�{�������=���a��ίQ�Tt?�h���=,T�w_48ZH� ����R���}Q�}ΪK�e�xpu���oyW:�qIԝ)t�jzDXB�j�M /����Һ]�x�8}����ȸ�3y�Ȧ3��=����.�~��~��
���Zw<��(4��Jp��)�ɳAl�24��q��T^��
�/��՗�3[��A*�Q��8�G���b��4���Y���h�q��|��6��8����N�~88��F� �c���������a&X?���r|Z�b�Y_������h�՝��0��)A�[N�������J{+����$�c)1&���*��<#�@�o��3G���'kX��8:K�Ns���eU��cޜ5r6S$�� -�Y��7P��q_�x�按Q�$��%��7��Y�`k1=��ل ����vG.��v�d���s�.����p�� ��20��Ӏ�q(_4�������E��rZ��� @4��[\r{�9,b�~`tR�~�@Yd�Y+e���3�)^��/r�@m}��T�5������ e��/"�2���/�at��3%�Pd�%cTW�4,��[�N� 5��C��h�ٟUƢ
�.�l%5+�,�����oq@���K��=!]��`�a�Z��
�m"A�T�x���+ TY�����T�{��A	<�2�y��
����a�~�����Y���O�J-ހ�~��g<�8�lЌ��I����涄��K&/�W/�ֱq$�!�\�1�d>����G���}@zN)�O��f�o�MT*cS�x����$�{La �������8�_�ʵM��>5ڔs|�~
�6��]{�S`������r��*z�F�L�D����U	t�n�����pQT7�EWvNjXЭ�'�Q�"�6l�y/�w��Պ몷Ă�5�;�@�ʧ�@�B�.up�[���k�@�0c��!��͎ �^#�0��g�Y�£�9p~����сq�(�`B�We1K{�~�Ĩ�=o#Rظ��h¦��Lwk��7��@B���,__�1����ǡ�&&����b�d�����z#ڕ�Ÿ���t�ĸ�O�?��SJ|�,�D��~rI}��7�u�Q�H�`����|\���4%������+�J66�G03˸m�%%�/����=�ߓ~(܌P%r���WN�Qτ�u�d
�0��� �̹,�����jH[ԅy��H+������ee9�[4Z��Cm�k�bo|U�6H�+�
9K������N�e�~;ډ�=f4̕�w#�n6?�&G�+R���27�廷
���G��D�x���}�ؠ5I�����4��.]�=����[�F������
���`7S@��p����Li�c2iƲMi����U�#�����l�&n�ݖ,�A������մqO�P,,�:�����<f7��M�$�ߧ��+>��Jȓȣ>��]�DJ�ol�ʞwMY�Ѝx���h�j�qy�^���:�K��¢U��m}Kg^����6��}�:�ZkA�uj6��/+�G���h�8�p�@���!}�2��+��<&�u9
��)K��[�f�T+���C���k<����$Gm�W=�>�.��$Њ&A���6/�Ʀ˕~��80��5�1��te��J����(]}��y�����z�me��=A��7�����k�<9�^�e�'�5%t��,Jðp���p�hK��Q�m�?�-�b��)"5y��Bq�b�W9���9D-��t�٤��1��d��@Q&��-Ki:)V#�V��8{
��hp_���aWcs��M��U��lr:��h�����E�G�I[`���i�'b,u|��1`����Q������d�o�S4	�-�Vi� ii��p֖��#�Z�\��9}ĝ`�N�����ʍ)��as	о�Z]��=�\��w!ZLvͼ��r	4Q?��),M�hC�e��D&�̿��\�)�~_^��`~�"F��U�nuJ�h��C�Z�
WEY}H����}�ב���F�>��Ç,�u)3Xt��%,M�P��,>b^���"GIkg,/�v�p��8cZf���+��6|F\�]�<�hYo�R�m9�tZ�@7���^3��]�&�g��_MmG�Zr��&�V��,� �c]��9��eŐ�Rȟo �ٹ���;��~�Q-�;�jd���2�0\t
��Ȣ���n�;^�� o�1$w����O��ki����m��=Ҩ	G�]���[�Â��[�u�m���sN�O�R�wU3�:^�0P,̒�D`�nT�#�z۩Htt��������*����a�9�U�0����*�[?�:{L�_��v
n!!N��G�m����[���Ӈm\{�?`�����n��If�h�"d��"�D�u6S.*���3�(؄��&� ��'��t��@X��_P�V��EiS�s,�rq�(�������p9\���� �+	cI����?�~N�Y��;\#�Ԅ_��R�_��;����	`�"�����K��c^U���H#�m����th!Eb
�  l�g�t�}̽��y�'�]1���[�\]�'��{������	Km���L(͏����PTP���0f��2��i��]�#�ǾQ r��y�-}���!^���K�O��'Kޱ���?L���Uθu�/�xҠ��o��Z~'��Dd�T#u'.id:�Xt6_��#��D�v������M�=�2Q�Cbdf�V�/_��KD����k����;��=��z�����6���f
��oE	�\�Q��[r9��
*)��"�RR$?8��("��c%ʟa���a�U6�Q*rPs��GR�Y5'��/���o��Y����͉B�"�����rS�����w��&	�����<�D;O(�u�a0����Dd�)r9��쁬2/>��'��jp�o�����%�|5�9?�� �r&���)xW�#uD�(X�a�ͤ���-fd�Z1�ݐ�
3���K�e��[��r�Z��`��/Άl/�v�VP�Q�����6h~��dw����)��񅁞��Ɣ�7\S�2�J_~�����ՠ��=��»pA������zs�ū
}S˝����V�rj� Mh2)3�I%d�gO�a*�%���;�#�Uþ�Suo�>���e&�T_�P�:<u����lEp��c��;�F��WA� ��ŅV��F~'�BE��J ��5=�����{�#���Hq[T409ZU�u�Upx����VA ����#��&���"�V��&�9M�j�9	��� �u/�
=�ˁV�1�:�9-�6�N�g�?pl!YG�$�1���&%(�3Ԛ�hH(��'-!�˧<�d��햾ҹ#6�<XNs?�t��c�~X���@��S����3$ު
�y"�`s��x;�	Գ2��3���������Ċ�o�',�qV���ñ��nNA�ҭVg�ܔ��?�Ѣ�V �\Უ�!�~��[x�A�k�R��Ȏ.��FN�U�[��#�-�Ӵ�-h�Ӌ���K���l-�^�E�~�����ɤV�+�_2oo*�*ă�G	(���	������r�=T�1����Rқ���^�]��ÉP���X�ñ�9o5U��P��2�s�`�ىqm�-����!��}?3O��?��>�����.�7>,�w��X�.�zY�d�;�$X|MX��%�+�+.��Sz.��9���>�}�,�(x�����bg. �W�[�𵑺7ze�"����F+��{[�g����<IݗQ8$[-�W]�^�" ��0BsU�)��D��Wl{��ܯ�B<�+G_��8�nh?ڍ�o��b�<��èE����S@�@��zt��$.Y�B��Q 
��Ҟ�ϓ]�Ǡ��S+��p%
�������nƋ6��h���כU
�h���_�K%�L�
���������Oo�t�u��D��]��s/�.�f��i��GG�l�-�|)�V�L��,oHʯ�F7����b�ny�9�����n�']$�������������t��eM��#�B��P�%R�Ǵ)a���9���%`����	R�!`��Fk�fΑ�-9���)��r���%+���g��q�ie/v��I��(���Y���	�Ec������$q����!�	7����T3٨H�M�շ�������cSL��'�FHE.E(F���~�xF��'R�r���٠n�դ�S�����������:����o뭃��y5�{�m�ې�UXd�^�C�� =g.��٢��G$joj"U���{�W��r�)�S�d�Ə�"tV��PX�8�&9��b-l(�lU"���k:6Ca͉^�@X��L���?�lt�w��yK$��lc-�-�����̇eU�2�l�x�\� �MJ�˕��VH��x��9��-���R �F��%TI��cM*�ccG�Y�[8��3��w �p��1�i���[=C��X^��g��"FA���"���w}-�%x�I�_��|��5���%0�e.Zj��ҙ�����R�Mޏi�a{?�������; ���5�P�+�W}�btF�n��b��HCyP�7�1]����埽\�1�~�`p� �������n��F��mR@�ɵnI� �Ц�ZQԐc!�\��?U����9�HK-7Sx0�WS����"<FL2'�}�[�|��$ �(��7��b�)�7�Y�1���(��������>��^:F��,r�����_W�O��*s`<*;�a��=�O���љ(��z6�?�t����g��XƜ!����wI�N�q*E�%��~>�'�YeOZ�E���6��X�>}���+�M�^EQ�߇�NM�k��KӇ5��m������Pa�vfF9�׎�~bP��g'��:�I�ܤ�Hs|�%�crT"���ז��VQ�V��!�!�2�r4fbt����]	�l����at��&�䄱m'�|�ZT|m1Pv���
i/�i$�㠇�*q�t9ظ������_ �gu��̞=ة��H"*>"D�݉�#ư�@|%���Rk`���+�Mv�}u-��5���KO_rn5��������t���h1������\��X�|�C�֚���ogk�����ԱjŌ�"�zPf�"��(I���GŚt���3}ވ �o���D3�32�����ޖO3|�� n�s�y:5>�17Ձk/,ۣ<���lA0 �V<��iq����k�8�eBh��|�1�76y�!j�<�R)��*1C��^����og��|6J#����.>���*���i���B]����=��t
2��%(���c�P� k�|O
 ��(a���3���pk+���0���&�J�{�cOhUa�\��1��t���r�tc:�faI�J.��E�I�7���S�4͎�8Z2?���Δ�E���^?Pt��'%g2��X��8I�~��:��t��.�Jָ�`��j����t���m�k$��G�� �rj.t!e-�z��u6�� RY�ґ��zÊ���=��]bӮ�8�%��Y�u(�������E���-��Tn���:6ʙ���D]-;�Ǎ�"���ğb���]�)��w`�s0��b�Q}�s�(��5|�K]E��q�|��Nc�򮝰.#G�IS��1{�`~
�����S�1�_��vE�a�pi.�:�x�f�fa��1�g�&.J#�_B �����X't�-��d׸���#�F�� [��E���)c�Vo����D�b���e��ăې^�9� �̋>N�Va�^���'�Uj�f��� @�{��/��j��0`,7o�v�k�y���{,=�������I���]��$w�Xz&P6�5Q��Q��0/�p=3,���K3l���tc��r���ΡeT�g�+Hp�DƤg�񰾮�-�_Ljg�[q���KG�GE]��Ɲ�@��Q��L�РiI�t��.7>����2�t����?��[.��YU�����Gv�eM(L�N+*��X^��҃F>�鼅1+�] ������֑�_�[po,~zX�E?}/��
%Zw1�J��#��)��`+��E~k���0D)z|�D�a�y|Q+�Z25�͵����U]A��I_1(x�'��ZR��3:y��H�t�p���)B�[�Qq�_o&���Fb��Ud��J��(x�e�k�Ά^�h�9��TY$�YOy�xQ/�/kN<��߆�;�>h��T���=]cr�T:���v��C�1�'���{�,ɀ�h�;�ڱΟs��M�JyI�#��B����C�)�������~��������O$�~6�����|I�&e�t��s�Y������<��0u��P���l%TȳD�QG6ox#�׋e���M5��o�~|lU�O*�����5C���m���\"46J�$TO��)yF���8�O},�M������'����?k�G0bC����|*\�%4Mo�o���jg�Y�0�<��R<�h��
A8I���g�\�4�	Z����Q�/E�!����������6��n�q�e�9��h�j/�01�,�ؓgs�rJ�`�"V��p���v�[[�.���;3���U��j$��ϻ��S ���q�̪:ј�\��w�^���,C�gFO�.�I�fӬ� ZH
��v"m�M���H+Þ��Z�;��G���1{�8�'�` p��v
�g������GaƁ�,�OIO\��m�w�e�a8����-�a&�"�2�Fe�'t����1���J�&�?	��ٰq��,_�-��I�*WJؤ���I�ܕ��0�)�^&� ��y烤���G`��*W�n�������5���xOP-t��}�bs#��j��$.�N;��KN{��+qY���n��QI�F8�5 ��0�Ɠ����^�(�E��N�ƣ�������u�B_/�$���y��9o��� ��;�"g}�PQ��ջM�m+a�%#�5���g?�DRJJfD]iuK�LH�_#����ϐ%��)���ggw�	��M�}%p�U#�i;�i	����_��hM�:���e��vE�_8�[d�,?xr&�����K6������hIp��"��xۚ�j���S�+_*�(<����̔�̝v�׎�~,'�'�Ե��5�Dу�S�N=�G���J�Ps���8���7�J�c�(~�ρc��ݹM��e����v��S�٢��)=	������G��O������B�n+�~š�`e�I�R���/04�A?d������~)}Q
VW��P�[�ȋ������Ȱ�ԃ��}�T����2��4�9�����m���y���B�2V��@"���c���:���1�5��U�!^�E�d��(i�H�^2�T��b�Q�En��U���m�~�%2޷��t�\KZR�'Z0��PW��P�U
�m[UL\ӞzZu��{4�+ܹ&"9@��b?/3��o&���܇! �g�g�-���K:�	���k��{H�&,����єF��6�����-@f�,��9m���Ep�j{�י��{�dCFj��c'���4E�Et��a�(�m��@0�n���kFF�$(A<������L˒P���#���k��k��a5g��[މ6&�4�5{��`��"��U��,!�X,f���^��>��nQ
4wM��B�}YFB����I�̨
�1n�HJ>������z~>sf�����}�;�ǃ`�-ғ�]��5����� O�*t��N�6�n8#�G����%s�^�r��P2��V,�ܴ)|xb��|T}ї���#9xQ���E@�X_�ifq]�O���W�o�*�a�%����u8�E�u����^:��}�tO�&w�`i ��k�vls~/3��N�[s��Y�j0)�z;в��^�=H:�ؔU��K�� �h�/��\z�>	� ��Z�%EWWO��v�֣$�^y�$;�-H��H���U��܃wKd`�x�=ޑ�"�8�hW��0XQ�r!������i��Z+}i	U��δ|b;�i�3ZlJ�V-c:���Y�i��j�.��b�K�7Vb���b{xT��Kb%6��1g�Z Bq �'�a���3ʫ%�db����F� A\r���>��N 3��B�c����*.Ƀ������寊�U��M��с u3�-�OXmO���>i�K�C̹��-�������>�}O˦q	n���N��[����z�,�U�`�����P�4� �XL�%/<SY��eD[CA^0��B�?�����4 r^��"�Ͱ?�/�:X�[1�t±�ƤО��I~�y(�Nv�POO��솖&1_GH,�ƫ�st��u+��� J��)*y���a"���a#��	|�Ab��� ��ԅW���G��Z�j>�K�[S(��=� �8x�|��5X��ȧ`S����!�\ܲ+@�=�80��gzS�-}7�5�^�H�p���sn�9�5�/k��ސ�0��:2'w$v�=�����{�;^.��Ȍv����9��$5�O��毰��x�X6��F�Si�S'��/g6�@+ �h��f��C)��8��Ν���Z�K,K�2k�����XO������M�(*ELt����)`qd>�v��D��SȥԱr���e��D��S��ɀv��?6���-�:nU��`V�A����~�!�����I�w�T�eڮň|�#eJgq�UU�}����gn��Z%#�.�F�;��j#����S��������d�*[���\�6y���$�r6����t��5*Am����=9i�e��\����9rS��M���;����m��-��"�_�	,?�u��|-[1n�:��*��3��k��)����4}���V/@��\~o�G�I�sa�����Wt���L�/�E�&��w-��h�vW	��[.B�:b�ݚ?4~�N+���_|L�D���
C�)�s����̰$9
�\� ���l9K��_�v�yɶ������މ6��V83�?~=�!U`6$kb�a�>����B�� �=!�6�������^v�� ��o��2Q�ft����_�L���G�鴘�*Z���YB��}����찹��U|,.>���'�yC�B� ���=.'����D�A�F��=�C�"�Ϡ��&=�;q�M�jb���F�n0�'d#]��$e��.v�({�P�`Kі��G�h�$s,��w�ĥ�#���KV)=�UvȐv�9�j_-�ᄆ<�X�tyg%"�hg�j��|�N}h����ĩW0q�hom�sREy���a��"��í�I�fLz�cW��v|}��������l��7��nuĠ��:(F�<֌�,���0�/3/ۯ0��໩Ǵ�&��P؎�Q=ҦT�n����?e��6w|�/`E����'iM�}���"E"w�?�;���i�o|���BE�a'�}/��9��H^�*A��W=	q�g�ҥ����u)l)"��dB7�� ��1��e�W��H��i����m�)�p H�Nf���~�h�~�/��-ߜӆ{.�j�"B��?����=�K�]N^�i�DI�`F�:ߡu#�q��<0��G�Nb	��K��gJ8�NtZ�c�S�ѭ�c�-�m� �(*���6��7�⿛��j��(e}��h�x���t����򌎎����!e�)����0�����Z;\_����@�y�쎳#?����MD�~4?�\_���|U�P?֕�t��f�����Oׄp�s~��,�/'��\v>QZ�Fփ)��)@p|ߠ4�
�WY��f�I�_>6��uy���@P�-؉J��B��僌���ᴢi
	�a<�#�$뵒qPi�͐�0Xڞ���-j��TA��	�ym�)N���2�s�O� �9[�����`�
��N��3������u��d���U��G�Z�/�{��'y/��+s娹N2G(��S#�~?I�Pfr���H�G [��/�/j�`�2�����,n
���&�%�盖r�{P2����q�}#B:ܲ�\��eW|��qK��T�A�C���7g)-�т�c�{Qm#�"f���S��t��N�ΏKҋ{
��
���a.����IH����gu�aQ��<�5��$l{}z;��j��B����T���E�ҝ��Q?r�@�b�d�R9�2������eɳ	'��G5o�o�9��}��"��he��� �����~w�9ۓn1m�������;���C,F�%�߹b��2{�3P�<����Mg�j�q��~$cd �C�M���2�=��S��~��q��f�3�Ⱦj��qYq�7�X@P"=!~Z�"��Q8h��s��A]RH�9m�3�cQ.��[:���jtj��ed�)�"{K�S(")Lx�O ˋ�Q���;0����,��o�c>;��:=9�������W�X��|zyIv�ve�R���mC�.M�������:�yw狃�m��5e��S^�n�d��8ܝ�-]��o�<1�?8�,�����l�P�{��nTZ�=�� dR� �E^}ʖ���0���k5���{w�IV�����#��o��o[�UF�lr���~�O��H�e;hJ��!�����Ы3T�P���A�\f�&W!c��=��i\�����9���"�V�!�5kW0x]C���ODZ��m6��y*��.����xH�sg1�*
�2Nj�|1�í,���Q�Ul82��&�w�e���̉���婠�mS��o�s("z�q����\�����R�+������z����� A�w��^&���e�_�G�C�vz�i5�8��r�tÌ���e���1�vk��}���T��Y�c�oтíK�+���+H��,w�V�Q��#�^��ëv z���4���f�ܪ �P�,����"X���P��rU-VD�`:�� A^ĸ�c=ۛ���Þ'U!8?'��	��1�>Bѣ��6u�e��Vr�"���7N KL�%�/"��q���Co�i���0T�}2E�t����uč�f�5O�[?�@�;oj^'*앫��R_�m��tB�,f���z���բ��BS��#Wj�@��vy�S��3���}�^����0�S}�5�����y��(�@��Ţ(�<�����5�C�@��yTi~�/�]�BM�:�����1����v�BJR��b��f�����UA��{�8�H��;pP�go�3P�r�M����&�0�,\��N����M ��I#�����J4����z㊹*����������ƕ�������N��,���e��'��j����h*���R��9EHk �������F�D��� +v�W����8]K���t�x���vl77b���.1�>�|Q��z@��ɡُX�Kr1���"�F���^�46��:�~��4��ɞ���M��.���L�6m��\��V;]	�Y"��%	�/��<�1l#a�wD�
%��Us�)��%�q����ւ��U��Y<�ϲ������m;DSMxd��-�Xw���<���|<]q���'�ʞH/�H���D���W�?X/�5°�����t1��7�bjĝ�f'c���ڹY��ϓ~7����t4l���k��b}�C:�@��3�:��:��1r^~[�m��!��:7O1��(���+��`ir�
9OtΙ�B�6\7@�=ʺ�p�|zS�L�R���_�J@�"	���or6�=j��bQ��m�P��꫔~B�S:�N(X���퉖��>X��+���^�R�<���޽l��M`�]R2jM���)V�����آ Zɞ#��g��'S�q(�L��PIX���G_��+z����s!r1?��l�L|g̨���2��kL����V�I�9��,|�|���,��R�[+E��f���U�I�MPq^-~H݋kE�w�)�Mm��Ջ!7�7�?,n�g�	��>$��@�a�N�+ee@�>�Sdo�$V��2���0�� �MGZ?�b���:�-���
8�	!�[� �v-$A]\�(��E����[���ϭ�����ż_��3���٣�,9o�qK�j�tut�������Yu�@ZF����i����{3>P��H��d}A��6�1-�ڃ.���7*��'�j%Ur��
n���zu�k�K�B������B��,C���h�R-�	���|a�/jto�%�׊���ٝd*�Ve��j�ސ�$�+r��C]8�N8Q�	���U�tQ-7\�Ji/�����LU4k��VT�`�T�-�!+�
�@�����*+�C���'"�P���&�hI}������*Y�6\�a�uK��;�GU���j�I��k5��+.�8�90�@�A��G|������ ���Z��j]�NY�mو$GBI�ү���E|P��Mk 13���e��()w������5<K�Ǜ�@m�s�ڱ��-*�A:�{��2&M�"oPv��œ�<���� ܥ�Iv2�s��n�3%z�;�W�><���%��t</�1�oW�[�{Y?�-*t���M�Yf�j��) ��]B�^��"�z�Ȑ�)،n���;Qf�i�2�,R,[t_�挙Zv�k��O�:�p|j��p���0EN���q��p�ia�ۃ�5)e��0ę�u�p��N
9�w�#}ߘb�ze�Viʴ��Tvs��[B���c�Ԗ�?w$	 Y9g����;����J����{��G�s@U�G\�/D��S���?��_���0�?��h�R�рO�Y���;i`�"j�Ǥ�%�:h{����X�	A�)�ď��5y���L;A舖���H���77禫fM����\�<_Kw8~x,�!ȡQkm}�z�W|)�>�h���|_�D�$�S䂷}+�4SZ��[��t/{ej��>����w�������Rɹt�,&EK�5���9�<����v��,�3V@u��&��<f�S�q)��,pQ�f3�Bj��J8��l2�,�	-ܫ�8�l�V=�]���B[�����l��.e�ь��F�{	�pXpJ�v� �������i�A-�9!���'�P�,HǾ�4�E�Y0��-�B������O�.>�g��
���؉���^#��� �]Pfȿ��b�c>m3c}݇�M���m��̛�q�����7����;g�B�NHn�t���_��<�[q&��|��8�)֛?�Ƌ����L�-zų�3`��<���JC+�ۍaJ�_=�����,�38j3qɇH�p�]v�8��qqFEP#�ւ�	d�.Ľ(�]��O�y�9$�8�/�Ra��}�I��u�(�
�.?�Ⱦ�%�֥��t}5�o����R��vg�_�Xcs�J�V_�8<���G!t�O����m��u��]�����*ʬ�΃g�l>T�-(ڹ�i�_b��H��W9�� F�/����B�b�4�g���$ �wAN��#��6��ޡ��-JaMf�/�,a��̣�xGMs9M�F�7�Z�:[�b;��L��	i�6=�����RVB|?8�ŮvK���ܪ9�ʓ��8"XuK^�ҺyS�gAg��+[	yYD�|O����~�1VݖS�����.G5�o���)�7A���l|�U�_FÜ�0�Ɖ��� ��RI��I�%�p\GE�+\�
�D]�_=q��q�,�/�_t���~e8I	���j�����9@�$��
#r�8Z��v��<l��6��*�D����^��N�	�Q�]��rh칂��]j�p{��k��^�&�9�M�I��8P�^k�m�h�����;�������dFֹ�VC�z4������v��&ẹ�o"1��t����=��[ׇ�5X�rz�Y2f� ���z�g��[^V��PbW��`n���&G�}�񰊦0mw4�Ϭ���V� g�۷�o�����n/��ʦ���4�\tV��T4��ɔǨY�`�L�$�͟d5�QA�����Wn��3'^�O�P+li�d��77~���3 ;^@Q���(DBTxq�~9�?����d�F�_E~�˧�µ�ގTj�Q>�W%X�:"x�&0� tl��YO����X��/�
����R?���*���t���4ȟ����#ˣ�#b�2e�x���=��O�_�(��&E���F@�je����R$�m�r��+�B"Y�2�������!�+�����s,]�V�v��ס���!Yޔ�?%:��O�L��Y1Z���Ã7���X>: "�">n&�'wĩ�L��r	,�ԾEjVL�L�]�v���`�j��&������m�R�o�<M�?��n�i=��C�^�PO���T��p�ۍ5&=�@�q�_� z���}�c�3���2���������g�cW�p#��{�g�7�eɤ98R�7,״��r���$�Ԝ��ә&'�A���0��kc��9{����gx�y�m����[�T1�a�����W��<3�`a��;�}̨?G\��J[ ��0����	� �����rQ�cmY�S+'�&Q�}�� 1�� ���5�T���Q�|�η���ܕ�E���w󤳯-@;u�_G�v#��1�d���1�E7��&��`j"��ln���޹=޽g�`/r���"G�����?��Λ���zX��XeF每���� �OP�L���$� ���1⋀U��s����E�E��2�6�n
^�����d�I������*�(#����vL����n�̶{K^c��o]�7�x.�#��.��V����N9�u�4<�ڎ'�-���d��Y�鿋8�����4���@(���`�RA�&49���Ա��%vr�$��`�
��*`��.KҐ�&I9; �م�̱�
�Cg��3�|0d�o��.�9&b���F�Bmq� �v������<�9�FKD+���փ	��\�1a.�o�n�4���Q�M�T���on��� �z�!� ^��9�?4�l;)�6�,�{1X�~q��I�]��1S3�����
��ґtL��"��.B�h<��+ 0�𰌇T����SO���d��C��=�W·漽��렁��$��\))%b�a���w�HKHq;�0���LJƕ��̞�Z�Q�u�pPU��w>��ӵ%�cj�Q"�1��t���LU����#��Ȋ#��zK�|M�ۭ�T���Y\�b�^L�8�W&�4�ިɪO�/�2\&X΅
��_��K�vVX�R<oYu4z�Uu-D�Tߘ�j؅򄘛U �9^��V-O.��\~��%[hU1� ���`��j�]��"h���d�i��ur�����Pjd�������uyLv<�֦�T��x���mO�~뜂m��P[i~��'�F)W���rO��~���yL��v�*�1�8�^����Wk�"�)x���k�F��͍��0n�������3o9A����.�g^��,���]!X ��4քRr�/�ـ���vg���m II�G�R�0��%���!j�jIcd,"�ڵ]����������49��I=�,c��p���<���9�J�_g�fO^��;d��+�'l�B2�(����AϪ�l=��h�W���wU�=@�#�6:j���f�b�B���$@U��6fA �]�/I3���޳T�S�\��nGKx�;Zvk8>��y%���?��B˶Ϙ�/Fu�s�v�É�9[`#P7c]�`L׫��x)BE)�y���n$0���	���f���ڢ� �l��I��Qd�M	�K�>��U����D�M��~~��s�s���y�x�xsCO���z�H�<�x�S�,�����%���\�ȈP�yR+veJ7�a4�/pW�#��B��z���̽3�i�߉�ZM�?B��	A�'|zl}Ȓ�F&7�M&��y+��<�@�n.�?�%��x��ti!7�����լ�F���A�`&sq&H�,?>���{��=JL@:r�|D�W��0�0[�ϳ 9 u:��|%���L��@�����^Lj[�i���v�6��h���@����ܬv�<�Fn�c��]�1��?2�' 5�8�薽��ȥ�	�#�˯$X��S�����NeR�ڎ�D�yAbFuTX�w^+X�S�`͟#�j�%�t�n��V�ɬ��p��?^���j�����1�"	�3�#�!�fYA���W)^S&)�4-��ą�1�����T�=����k">����Kq�k?;�7A:�;k acjM
[�Z����ŲW~�g����
���$!Z�|�P�B�T��JA+m���__9R�Z�����Ƣ��b݂X�_��4-�I���>�wʇ��p�iBާBx�-�s����q-�v����
yL}����}$����[1}��QkK�*n|����y�-l��[a�$"���4�ţ|�`���NR����V��6o�cY!�&�ԀW|�S�L$ǽk%k��ǩQn�eQ�_�n*�A�s�$E��33��J#�1�������=��|gn��ђ͕-�3�DH��	��
@��WA~��^��ba�|�3��\"C")�|���"���8�e�m~��Fݕ.��]��>�:��)��1��U��z��3�����aT>�r�c�&�RM����6�������M�K�)�)�e�h�+�Y0m����r�H���/��8���m7E��Ĳ�K�����(�ŲV���$oCf��Ӥ<@��LXq'��*����{U����fQskVbp�}<��Q�p,�����]�~��#��W&-����˱�a_j&Ǎ����T]N>�!�GX�����khQ�6W���6���?-\�6ϧ���B�A_ٍ���x9��zKs,��y��$#8��v�}�Y�	m/e��M�J�(y�R͗���*��.���VX�