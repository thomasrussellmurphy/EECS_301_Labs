��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\���V�fnvx��ÍG_;�ȅe�~�>���9�>��Y;�0G;���u_֘�Α���(�(C�nd�����Jd��T���(h�v����K,�ߪT#!�1�v�����|P?��H.�+��م/���]�%?��I���oC�\��|eoyo������\_К�X�Z�1����8�b,��)����ڏ�а�.Ԅ����ߊO(�f)(T�0����"��>U�=ȸ[$���͌���G�C'�3H����c~���'��X�L㽋��#&mZ��;��4)���c\7Tn]�Z����!z��1j9�51�0�W�c[yY�G������Y��W �MϲT������Z��Ģ�"2�Þkb!�C�?sÖ߭A��}D�q�k��̗B��p�y�[fS4ɐ���ȳ����[
��:��G��g:��@�W��f�T1�+g��/&�l�pe�[6�Cf����S��.j�מ@Q�$����F�$�#C#��m
�l�ɎX� -6��(���M�Q�\� � �'�{��PǞܡ����t1t�D4J���QδF�����`�%��-���S�v��o'a���	�xpT^b#�����o���j��e�={�4���x��f�'�Y�K\�
�q|l�ǲv�֜.\�RZ�ſ�V+s��ʖM��&���{t�y��j0�������ghM]�`0KݏN�/�K�Ź��C���{S��H-X٧��/�q��c"N��䗵�9Z��:��uөK[����>g�j����#s������Wk�:��o$��>]&�ޥ�1*;���1�z\�群�6'N��|������C�O���ߡX"��\aQ�]C#{=w� ��U�e�`�䄹��wn��N��Q�kG�؞����h���D���"��DH~�P	x6Z�2U
�q�2�v��w�ܡ+1����3�I�b��<u����?J�ǔ>���r�'yy��^��>tG3�q�?�C��v::�w�\O��`��V,��<�5 ���ì��KeA��"�����ߗ�scO���xq�>F"D��V���(z�� fɌ��JJY[l5Xp6{��0"��0���J�;&���noi���WN���{�o4��O >I�8B<\}�l/7���*c�Ζ�pݫ2��{ﶕ}E�T�/Z��X��V�����J
5
�i�{����ڟ�=	5��S�_�[Lp��4���	� ���<��+P�Ęa-�8��'1�*�M���s�*@k˹��Zͪ��C�pm�<�~���3q�:�8�&ᆋ��x��ݖ%�
�a84eFP7-5rO���j��f;JF�@�w��'������W��s�j+��_����\n��m���껦;NN��l���*�����B]_�EK�G]�zn����i9؅����u��4@Ŭ���d5�X�Ia-���iZ�Nh�Ǯ<��4��$�Ir��;�Z�G����SV\	��B5��J��t�Ԃ���9�tט���O��p�~��n�����gt2����m�z0����ZWt����+��		������g!��2P�mh�s8���+g�#�O"�T��^+�^���!��<��Z��(=����m�o��͊0Eұ�G�U��� �Ux)5�Q�j�닩p�	/���,4�A�N�bF~L�L�
p�K��M�v���PqX�k!)�u���Ah�Dy8���%Q�G�;���ߺ3f@��V�`F_��J��gO�Ҍ~���J>Sa:��w�^c4�"����oiW��T�����M�e���׷]��M�J*-ZxU~�6��k��y��|nL��*�j�{8=^͉
�:�:5 �3���q.�n�������UQg�E)J�+i��,�*lǢ����-�4��{/�3��q"�i�_�&l��f����I˥_�}����R�t+�4f��ԫN�DQ����*i&is`��.����ػ�-E0}!퓫S�������yy%t���D��ӊ�z��y/���H�����B٧��k��}������"��V��n\z���.:T��lLh&VZ�E�av��x.&F5����+�Q���i�`,[Q��iWq��o���4�G2h(��f��X(Zh��65B����*���
,���{.�˷ r��6}W�6p�h*����=x������M9�)wj�$
A��d��=_��H��Dߣ]Z�x��b�JsI�çbD[���S�c��2L![���K��������U
1�}���
� \D��׀>��J�����))&�L��1OQ�#�ʺC\)?=�pjN��aM1��'�f�{��"Ce���B�U;�����{�D���s;CM�[�����dP�<�/x(�2�N��v>�zNf��X�w��Π54�Ճ�����, ���R3�n{]�Fg��Uɑ �s_�o��v`�m;�B�p'��<�F�>*f=���5���`
�)旡����i���"�?����PAL��#�|�}��o�Mq����]�rhT�v:���\��IC��n(��Jw�;�֠�b��Ձ׆��͵a%��\��������Bm4�&�I䀓}�NY����Rl�K�ǠWz����e�ҌB84��
�����Е�Э�QIQ�H��T����e�{c���g29�6�-�Ex��(XCi+��^��Rφ����qzb/�6łW���������w�Ҷ�,��EkiD��ف���}c�����J�c�!V#�yus�
�X�����\��-��������nO� �}C~Pъ���&Wþ�7m��^L5���/��$�<�]@��jk�I`��)C6�tZu�@Xr��F���{�������������]���aq���JS�
:o�Y`��[\��Ty��ߤ?�������S������iXE9���{��J��anґ�����>\�X�3�f(��^�2,�`���lɩ��5�)��Fs�O�׻���rBF6��*<�v�	��賆��(���7;nŃT"�TYJ�6,���f�*i�ՅhP�[���&h���iO�i�c����|��R�Y���$�[�HQES�T���n� �rL���/M�E2�P~c����ՠ�h�-�>�d����E�w0G�,��܌��!\�/��������Si����\�~����XB�����
�w���	iܴ2MJԣM�c�][���S
��!?R�:cR=,��l�k�yCz��.�K����L;p@	s���yl\� ,��#=��59�&p��la���[���/O��'z�k@;W8؇��6W�'�a=1L��ȵ~�k��93ɼI�-<���b�i
f����f���ГX�Ⱗ�=Kһ`V�&�����Ak��e0p��X������ܻ����1�/5�3:D��]�-I1v��*~R�ܢ�����BU����٘؊4H$I:��6�b-���)ͷ	�56� +ߔ%�����,�S	dI���[I�t���1(?���.b����|0�Z����I@�����!>O�''��øF\\y�0%�q8�a�{��3�.�c��g��3]�y����s#��Ϊ9���+���$}��e���P�&N��(��D~Ӟ�b��W"�CA�l� ������O/�� "k��ݪ0��s��x�UiTKsO
!���=�` ���mb����_��P{��Y��:e����kҝ����WkDK��^��v��V@�{�3V��^C�t�
H�N��;$�\<�}�uJ���ܤ�]rc�O���3�E�<�K>ֈ}��̰��4j�t�R��LU�d:�9�%�Q�v4��E>J�?�[K��0�a�<]��T����D���U�8=L��dݔ��և�^ގ����á���ʫ�7��w�;7�346�;�Z�#�)$�+)��y�d�>�SD����X2���!��=���#Cޢ �n;�$������jQ?	��/��P%�#d��0f�?�r��tE��V)�ݵ{1Lݘ����SR���>����3_r8�z��d%؛ne�2�3$�.튲|0�aK*aة��0�H���ix��@UD:>2jEn�ق ��q��]�B�2Ӵ.T�hS�{�4>��0�;����'NB`�ˏ
s�=��:��k3����QK���޴N�0���MZ�ph<I��)'f�.��@׋�B������[e�.k��q�Q�9��ù����նx-����p0��Ȱ�[��0��Dv@Y��w���(���q%~����_F���$!ka���qg!�M�\k��5�c�
�4 �Y�����b`+��8�F_�^�a,$sW}r{�R�9WY�\�[�<K4<���"���x��ō �sS<�L�(\�ɝC&�H����o^�N�y�i���>3';�}�7g�n⓷K�j壬H�H4���~PÔ/PZ�*a�gn�i�"UwOٟ�g��$����7k�IV������#���{	!ɑ��Rޯ4_�eL(�K+-�é
uK��ڣ` Wq���K���n���$Ҍ �8���R��z\�%�/&k#�׼�e��&��Fz�S�\���T��1���<H�kF@�{A<�WH�c�f������-�����ɪ:�άyܛ�$nj����Z������a��u�D^>"r��TD�f�wH��(����'���/�+�f	>�hu�Ex¹�6�e�$��뚟�M�3�i�s�tT�]��(.��#��ҷh�7EI���n���}L�Y	@�9'N5�K+�5Z4H����
Q4~�Iu�2��^R'���pD�P�r}%�� �i���5�����z�G����4��V� ͝�+� �ՏbM�N$R���`&���݆�<|��9)��"6+�'�ڀ������ ��+و+f�OPR�:���Y�	3���,�:�:�����<f���̴�[+�	c �SW��>�e�&p{������O��Žsh���X�h��M.jĨ�n�q� b�5�=F��Z�"
�)���X\��k��5 R̷�Ѝ�&4d�`R��E�D�}��h9��/����ԕz<�24��CF��gj���|���9�����y�[�3۔�r�7��~���(��hU�������m��i��M�w���q���J��E1��{*�0������l�k��LR��9��|���,bquh��jV�Gun	y0�mn3�O7����{��ԔA��&��gx�q���;�r���es�{�V��+���L,�O*'�#-�$ar�:���ܦ�*�^R�IZŊI�
��t)/�Qi8���1�|��<�)��v������	ɩ�hEܔUFL�=�<� a��Pv}{�Ԡ��l�'�9�C%�6&���n�$v�tk^s��U��k�(r�g~tu��M������[V��o�~X���a�(�]���7)l4�<<���7��Z~�a��Bz�����f��E(�V/���8q�������؅]~��U�	�B�3���s`g#�@��g�I����զJ����F jz�@\���a.o[fY9�/��0����2v�>c?���?
��w�,p=wC�mK�Ê��xk��0JT����UNpN *ӓ�#ܬ�-��<�<���I�"����Ȯ��/:��'��I�ɝ����pp�A��Hz7h�<h�d�\�$�BR���u0?=��{t�h~��iK-��!������T��wI@{'�@��R=I�z���N6��:�e�E�1ь�D�W�3yڄ�� Usc��
`���$[]��fr�lq&�ejR�l�����r	�Z|��k(��ׄT�+'�]sWZuv5z���Ͳ���t8?PKn!I1.T9��1F�4)���88����Z3���1��vk�e`0��x��G�EL����4�V���H��������I9�W��K�8YUJ��>�(�{ȷS[X�{���&�� �� ��p�B�������t�B���  5�l]ޱ|��� ɑf��K�sg�Ʊ������n�T�T͐o�H���,���pݚ��B��������V�q��\u$4R_�3Dh��>&̩��@�h�����,������6���Ʃ�R<+��dDȰ>3�Zg\l`�x���G�.��,Y���P�$��Lg�#^$�����mL���28�Li��c��$�TU��p�>�����.s�v8mn�����M�HY���)�c��-�ڜ�^0�e\"�ӣ�Z:�E�0��d�1�U��f'��1-�+9�G����N�/[�GN�V��^���6&&W��t,aم�M	x����dPO�Ջ����B52�1���g�V}��\�����v�v�|���o��m��r*��A2Z�+�����F��qɱ�'�o�R{��]]� Klo�K��1*��4r����;�WC�I�b�RTΤ�4�k��!��&� �u,$�k"r�r�jlA���<�^@�F���c��r6��Z��$�Be��ü%�U0�)�Sٱ�*2����5 8�oAe���c���uW�/�"�Dff��HسN�c:4�9@%!�6�$�;;�I�|�&��t�ũ�H�	���>���\��赙��Ѵ.���D�hE6���ew�T�ɏ�P������0�o��P3��9m�'�K  �c}V��d��iy��� r𷾛��d�J拤79�LD9
sR�u������S-�#_��x��,�.p�l���1� Ý{�����e�*�ɬ��2$*��D��p����T�넄0�{��H�	�a~\1���&4 DĦU��6u��5��˹��·Y��r*V�x����^{�&)������z	(�9��3GF�Yk���FEܨ,ѡc�a�A�Ph�AQ�5y�{�n�����A*��������M�5��pՉ�}kXӯ�}�t$B?_���e�����(�hE+
D����r2�ML�9�MY�� n�\ �O��0w�8C�v�{���)�p��l���%w#�(`���Z��w�{�[f�V��?RJ��	�C|64�y7o��ת�.Es_�?���ݨW �q0x/k�'=���2��A2��<��p�����������O�*xqU��0T��,��v�[T/�����SS�@ n�i��4)8U2���f����{�*�fkU�*g/)��ݔ�>��Mde�Mo�� 6n�������.�I�DP�J"����
V����#&��4�4d߭|��Hx��)�uXq�l�Z�/��<���$�Gv��0���	e`ܫxΎ�S�t,$q�:f@�v�WX��t����EM��T��15�u��kl��)�9�j�V��Fh����F��]�7�/o��P[�Du�X��r�T�[��03��VX�\�7�w7���l��S훜����Rq�Xnҏ'�X����4_y�@����yaCɂi����)_��cy-�1�xSi����U�p��T�I�(���RcZ-�z8��U��GsB-��-��k�rF��2J<i�v{v��H'=X�%�[������;�:���S�߭�Y=@�znG�/@���#��j��<]��0٦s�Z
����DP� �C��>x�r�2�}Q|vceԺp��ҁ��,v�:��\s\��˰�P��0�cjn����}Ua�ۛ��	ܼ@�1:�I,�9���k�'?���AZ)�n4���УuN*g�)R�'5�!��I�7_w�r^KILYĜK��<�k�my_��l��Z�o�-�4�Hް炷}А�I�2\C;8"�y�G0��d�3�W�������y�
����g�AU4Lw�C����m�ɘ�ĭgPw�%��\Z�kx@ɘz��a1��_S&3X�iS��C�� mS� �&�7{n����Yz�k/��E��Q˿
�7��:ܮ���y革N
~N�Fw����FC����4�^�a�g�ʮ�(�8���kӷ�	�B;���L;_B���Q2-5i\
��3�!�]����̅ټ��o�R��c6->��ѷۜ���}U׸h)l�Į��q�|1�P�yJd����P��s��u�W��S&�%�LǓ���8�$[.Ֆ�f4����.�ֻ��G�睆
�c�hV]_>