��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\���V�fnvx��ÍG_;�ȅe�~�>���9�>��Y;�0G���>��%����q� l@r�F��X�QM��\����#C¿\�U`���d�l�|�#s&�]��{2U��\�=k�;GTbZ��~YNܟɊ�#��!�#��G,��;��*M���j_���t�S��2���UT�PcK<��ԮKk�:hCQj(w"SY;�X݃�r����R���n����!�Dתp�%h����s�����8����ɺL�BMDN*�O�C�[ j.��bΖ܂޷�G���"O�O~�$Y�d0_�N�wE���`��l�	Z���@Zp3p��Ԣ=xS��ƣ����P�Tv_a0Z<Uܯ.t
8\9�	$t�����!AI�W~�����`��t��-������ZҟO��jX�
�~�+b�3�u���xZ��!�jip	柢�`�JS����Q�L���# ۡ�}��^T�T~B�����g�(�:�T/�j=;�h&��+}��PF������7	�J'dw��D� �����٨��;+�l7�S�V@����jb|[Q�/�|�>�q|����.�tt
]=y�V��)@�����2�a���*��U�m
�<��2
�e4��Db���F����Z�!���:ز/���p�'���#��V�}��1����g0�+�O�
ɣ�`Mr�L(��P���ɹ����6�J�; )��Δo���ihm׍��q�Q��^<T�7ɓ!2	�2BJ=���T��<d��i���7�7	�e�ZY]�2-�����OW�-�s0'<�9f������̔�Kl�"4�.-$��M�NzW����pf���\�6���)�lU���ޓ�7�%v[��8����ę�ˁ���+�@ca�^�ʘ�1ȴ3-�E������H�<����Us��Y\�
�+@`(�[ V!�o�~la�E��jö(LL��-���E�>v|�Ѳ��Ғ�( �@��* W}��:s��J%K(���}o�bx�rpR���emgpܺ�)����L��gfsMn��׹O�x��@���xn��㉜�ac
�d�ݸyu�ثt=����h�Aޒ���$E�!����kN�� 兦**nіѼ٘I���)�8$�} 	-F':����~�A�����L �!2����&����yA_SպzgS9�[v�q�խ�nA����g>Z��@�ꈎ4yY�W�O����^)�E����F��(0K�r�R;��f<	�b�%;�s6��Z��7?�x�OT�"Q?��F�3#p�X�鵓���Ϲ���(C�4S�z�������BI�����ƬO�@#L�F�z��3�B`4�=G�(�`2S�~�o��?1�Q�
��ۡ�h���� њ를�^'ܗ�^ڭ�F���q28f�B0��V� $E�Ř��&�/����^6n顇�������+�ˎ�X|k��@=�ќ	;���aN�`�yU�<.@O�*K��^�=kK�3�T���zO��	��^��Z�h÷>�ćF,�u*�"���z�s&�x�Y��N�V���^XA���ߕ��>9ů$�4*���2���ب_�+�0�����MԀ>n$� �#4�������, ��_�k�#�^�8A�ù�����2ǩt�lK2��r4���&џ�C�K~��a���d�{�d ���Ʉ�W��d-M�Q�O�Uj~>�8j0aĜ��,���Iis�b��<�������O�`p�D�h�=�1���|��o��~D��'C���������pFM#��Ɠ�,�5����5�5ijj�kҼ��ݲ0��^�ل���'/�ȣ�p5�V�W�U)�/���@��ut��8a/bd$�Y2r� ��̭|/|��N��Oܦ�3�����~í�C�^����.w��� a�]�,�D�k*p*� �+m�"��ک<d7RQ�%Ec�X�֠�����n�,�e����\g ZGM砭M�� =�!]�K��YO��*����p�*��+�|��X2�s��-�,�Gl�'���H���#���-����52':��	��0��2�Vwm��
X�c�HPK���&�o� ���g6�K�_Pf3X*��IU�$��Hv{���ou��kE#3t���lD�p��	�%{ۑ�r8dd}C P�X��9�����+�/��͋�L��(�G��"z&	M�T�eP�#4�R���@�{�xתp�������P��Z�R� �_����`����bԛ$!�\bm��Z�2��b��bهC/yUR���i�@D�)գY�~[{9��NT^�TU&�F�8�3Û�Mu�O���:�}�����hk���Vk���A�~D<#��}J�;�'��8�ڠU?��%k'�-^��m����g��T	���i��Bv�h]����l<��Kk!Վ�i������>X�td��+��u��G;��Eį����b���p:)�m�I��,0���^���_D:[3UF/U��*ޛCŞs����MG��<���}[o�̅��ƯUt�l�*�.���B���Ȳ�ۧ�Y�(�`�1�}��Nv����!���2{�N�7���H�e��ڶ�io8�� ,r�e;�&>SYy�����G��7��C�sQ�c�_MGq�%�r(fr����ɛ���(���0�W���j_se��y�wk��������䟪�m�i�>���&�U�qh�Ud��L��M�%�Mhg���(�$:�,/&�C��.h�%5
�D���^���h�����=��$j���b��?D�L����qG��6љC�z��;��E[[�rL���Z�g-2C�>Me/��=�QW�I(��V��J\��){����G �U�)��L�;�����bV$I�Nu�M�C��~`r}�
l����ðCҙ6���43�r1~����/�/s-��*M�u�.���Jw��3ţ/�3�c�Wϒ���/Tz�JRR��I�2���:o��(&'L7=r���^�N�(B��걌O��i�z��u[	f+�~�
�3ݮ�ٷ�k�~hy�J ҔJ�r���9���3�R�������} ����g�o�����SNLzњ'Q��������H�v�S\�S��:R9�j!��������@I<�0ì��{����S�%f;~O�c)�DvG&RlC�
���i�^S���Ы��ۙ'�G�x�H�7�N��\�u�%��1�=-1�9�Lz6(	����9����ಱp����=HD�
�O4y�ZW3�*#�B����yc�9���zO�S��nͫ>%�(�
�Pɚa.�#��JR�*&��B'
����+C���������4��0O��+	/d��>�i�y�)z�;cCm�J����H�G'��Y�����ˣ��r�k���_F���V/�`��q��pl��6"�C���~^��+o�7liXǜ�����<�2�/ͮ�'ߩu�Q
�|6HJ�-{pTj��y_`�)V_= hb�+3_����u���|���zsc�0]9�z�,C�`j(suT�r~��>-�AV\��'; ��Omh��+>�9@Ľsp(o<��h���Ib�ړ{i:�� �|v����D���Z'��6�m����g�y:�:���7uȳ������y�� �E�Q#���|Ġ`���m��+�S4	�Y��@��������L��}�C�������{:��?ɿ�/l�a����
�)��OYfƔ3��⒚կih�Ql)�gg�ybC;11m{9o��b��=�.�KK�H��krtV�Pػ�K����L#��I[��'Ȥ����r�2�Gg
S���v�Yu���E�3@e�R�G!���&�yHad	��pԮ���������I��C���48 �-��V�[4�"/��4cћ�]�D�3�i��hI��(�	��u��Aʐ
�w����?�Wco�6��2|�����M�!0����b�j��!����_��=�<���{Hg�"*�T!ß�X��
����+���2ΰ��[1�`S�ж0�$^迖��|O�ey5ȵv�[��h����6��d�&a�b���%��9�k8<�%2�=�i��EWC�@1�z��=�n5Z��l����R�	+#4�4��L�z�����囧pK����a�D���!eJ}���Lx�JA	a�A��Wvέsp^W�O�u��uU�=���?'����}L.A�Ӌx�T�������U,u8P����>OX�\Jw��.��X��?���;|�gd��М��)�c�i��K}P���e~��Y%k"�`B|G��	u0�x	���O2�����׬Y��GA��m�����k?�I'P5�DNC��rBH8-�n���Y�[�sۈo� z��7|(�{�����a�ڄY����zO�#�X���{�a��V������ϯ>�j=��|���'q�i|�-F�w�0}]`DAGI~���?=��A�F�*�Z�n�8�A��� �{BZ]�oz���a��k�C�	�����&`j���2�r��Q��`1���<�����u�z��r��(n��9�� v���GF���bV��'I�_��g&�+P�ڪ�h�M긂h���SR�h{�m��=j�����-�3;�C��G,H�;�8k^�ꂮWu�RSC^?j�.0M�����}=@ݓD.�D,p���=�	��h����۱C�|����^/ȣ<Y��T�������(xl��F�6v򨐩Z�'��M��V���/t�����ec}2�}�_\h/�͵��z�V�������>9m1QW��?����n�̖�Q�����dq��)}$w7���c'�M������+a�\�d���0
*8����7j��Y'��j���^��W�0]�!� SݒZ׊�?�����@W��Z�4�ق*�FT�Q݃��	�����A�7�K�u��,g~1����q����.�g77GJŚh�x;�BC�U�%z�<"�УH�����짎<?�W9uP�����&��*{i��D�j��S$$�XY[v�� ��5M��cly��F _�$�Z��#�޳�!��Y��>��Uhyf��R���kc�J9������>f�B�$H͋�a��:�0rg��99ُ�����l�Sm_�<�1���'1j!���{�[+������$,-��J���ʚ$7�=��6�l]�‷���E�V���������x�_�-#���5��6�i��B�}P^z5qD�o4ձm۫����1�R�9Qe��/l�x0���
��#��K����;���
�ݥ%]��R
���v;�����Q�lB���?�M��L��أΈ D�'u��5a���4X3Dn��$������j;�/���>
D<��a ƛ�#V�j���6?U�9�w�C]���o�b�i�����󲄁�������Z>�i4���gw�a��R�Up.�C�����ч��A�P����J���.B������8[��0h�����Ul�r�y���ع����Σ~�veAQ��.�_�$xO$�������]ۍf�t� �#�6`�[�Q�Gz��O�v�a1w�����"R/�d�xTRz��w��û��2��Ǣ0U�å53`:���b�#/}V@2�yBgm	�tg?�ɮ'T'�{�����87(ŖΏ���$N:��C���E!��V��&��3_��VB�� �^��j�<���}�`Hm�"�Zg'���W�$Ϭ���k�G^n���  �e���Ӱ����V��_��]*5·9n*�����-OFĜMOp$C�0h�����/2�f�m�F"�~�-yh��+nE0��h��� �#+����b��M|�T���'��<W�.&j�7�"0�'��Rc���ۃ�窺��8�L���y�e�c�} U��!��#!���.XȺ�}��{}d�((��T%f�b}M)N�g���NԻ��]"����e�� �0�/��h@(m��o�s�{��n0B�,�b���d�/�SBG{��N�ԗ|C ���;)n�@d���{q��&�gA'(�5�T�IQt��L�T&���!if4~�:�YN�nCؤD)k�J����D��`F<D^Qy�W����n�0_|����Xpm��N��f��pKk��������fk����c��
��=Wp�uN,u�����z�g���X:��Q���o��9�D��Wm�$C���?�X�"�E��~��+~�M���mx����������qx���M+W`v~n��2�
^!��#��d�����I
}&��t�R��M5\ �x���@�d>��IP.���%�*љ<*�u"8bh���"5�`<�gƳo���8�ŏ�x�i����
��D�3	����g�6GV�d��Mx�y���P;��oҙ� ��P��:\'��?��w@�%t�KBAO�/���k.��"�� �T肌��>����~�;w�!SO��$A�gN ��#Xx�n��G����DL�&$�4�)�mљ IM\�q����+e�PmqbvHq�4Gמ�uKVs\e`���X<�u���b./���)���6���҅�ݽ-D���R8�����>������K}e�~��"?9���e�);B�*�d��4�w�uT��O��|�߼D�q��s9}B ~��,�<�kY,�Z� .HG<����ڰK��"W�C��u%�u���(՘A�X�c߲�-l�Ee�.V\�; ���X�#��-j�C�o5��|eT]�5����yM.Q��g��]��S�!K�K����>��H���^Q�ꖔ%1��-32^i'Q��;�?��Ȣ������j�Z��f���/�=!�%������V�G:��M�̛��C/>�f��cQI����e 5
�
fa��k�z��zb�5�-	��X1օ�}�,��9| Q^M�8�T$nxl�2ͧOXG��u��.[fM��FZ$�)���r�bPi���bk����ʆ�Rg��\;�o��룀����<S����	�@8�Y���oE&P0�w<��Ѽ�~A���R#���o}�>�q%�R�b"�*�;�٭t���Z�qjC���8��5�&mD8C^	O(�YQh.�#cEЀM6eJ�yGQI�F\0.��eb�D��<poL������l�zE�1���[+T؏T�k��Қ��9��X�٬��t�;���/��m��ܢ�X9�$�T7��+�N����k܃�lDK'�I9|1�iw��R���E��a�Q���+���"���Z����Q�!<oZ	��<�B>OgKF��·�#���XZO>�^\)���7Y�h���G�kF�ޙH�ɻ���k������N�(+��������Z1��9��(ԖײXw �u�	�����;�x����X�*`����Y����7�ޜC%԰���q���(�2#���̣ǲ ����"�v2բ�F���p�zDH�J%Ns�FK�Nm$�k�4D4�Ib�ͼ� �e�^�1��8���Ώ��u��o��D�>!n�sjN��r'=8��N2s2-���0H�$}W���Z�jO'��{'g^C�:�˛5;�WdўLLN��hp�Q�$�����? �!�:=G�0���f��Z��A[���x� :����}k}�v�2�l��D�c@?2m�%
m;S �r����9�Ӈ��g�ˬ���}�,�bR��oG\5���͏E��_�� B����������ߵ�%YkH�d���"}0��C^�'b2��))�17[�A�z�����a '�XT(�X�y{@�@��ڨ�z}<�*���w;[�d��G?�ff�/�K9PǙҎP�Xb(���ny�ݖ�o�b���o�(Nr��9����d*�Z2����7�%��G&�S��g�y�S��T�b
wj�'��صw�`m	W|=e[��%p�q���ŏ�Qk�'6Z���?��؅@���(�h��)�b�BH:�If�P�y@����jVp{cԯ=bS#�g%�=��F搵�!j�,���NZ"2���v��3��F�߈UWU	�տߑ�����I���1w�R���p���&oc搩H�����弙�"�T�ΏD�K���(�`_5� �P�H�j�Z�F�*�H'�ֽ�Є����U�3/��D�A�g`;H�l3؜Q��W�4x��*�џ��j��i-�;b���7\=��E�������)�;�)���	]���E-�3�US1	�����`7Կ�Q��G?�#���^x��n�Շ�"y��t�O�8���5H��nj$���+o�^��ѽ(joQ����)��D;ؙmS_�c���<1XkFp�V��?K�iS�fA��(��j���R���Ԣ8����I�Zl��L#�ose���~�Q��nf#"�K*�3Q �I�@��/�;~E�>y���	�$���2R9�{�ǘn��'\�Ep���=� 9�}�09�Y���B4,V��Ed!N�c���!r�OJKZj�
BX�=��L*��b)��{���C���b����P(:�����^T|+!J����F�k�"1��J�aUJ���]P0�ɷv����)B=k)|����~�,c7�ӊ׸O�����}m���Dbnn.]�[
&��,~�6.���w�
��l��φ˘��h��N:5��F���!�C�un6Zu�w��~��Z/�6�U��AKix�D$���+nM����Ro����5R����4N��-6Mu?��j��^�s�	GKԼ�N�U�ۺы?�^�t��/$[�ճ
R|��<:'�xl���vi[�^OCN퀮����1:� 2T�k�򑎽���A���=�W¦&�1�ٱG�o�.�{���������6�Lp��[��'C8��c�o��2�^�;���_��;��`	s�Ep!����W<�L�T!rˣ�y��[+���z� ���Y:�ј�K!p]���Ռ�d��o9%Q߫I���z�n�N�
n���M�0��Ρ@�d�R�E��:���XQ%n��iz�����,-����0!� �F���]ب3��ht����gP�̃��]��ł���c�΁/����eTe���s���{,�hހ�+�}⑸Ѵm�+���h�g�C�h�X���V�0�g�n�g��7�faT�'�qR�o����:,-�j,�M=H�xټn���E҅ۮ�{F27��\��o�׎ ~0�q�F	i)xO9��>	����C*�1��s&K�j �[���'ܲ.k8���O�����7�qDb��V���s ���HQ�؂��k����Y�T����C�mp�t�}�l���fTZ��\�E0�ږ�!7#/�2�|5�b"/7E�~q�IR+��H[ɏ�D�`;:�ǲG�]5d����w�l+�C�]Ċ�sgz�k�����&WB�UO�HM{KKJ�=t?��*�?,�s08��F7�ע���S���D�i'[+l^*��A�>����wCk���aSP	��[G�R��8����/ř�o��Svc�و<�'s�]��܅[>�+�S��Z�M�W�B�=h���$�(����C�/�����վ)�Rw�,�N�CmA[gz���IL�����M��,Qp���*�=R}ۣ�9D"<�k���$=zz�v̝��hE��@-{�����$�����M���I��4�&SD�]/e���m�JN��S�ꊉ�@�z�H�ll����{\!��4�R����fk�om�^���n���64ms9�keHz!���18��gB?���Dd;.K2Ey$�sQ����
c�%%k�χ��;#�b2���?�#�����ȍKr�n�1^D/���	.c,�"����H�&=M�Ɛ��d�#�F�B"��L���}?�%d�$��=��1Tv 
����-kfH� �
g�}�.I>�gq���|�L�TORG��7��4�+��M�����̉~��HՌ	��{���\Jz����d'��-A����G�_6��<��k1Cm	w(�J�Z�Q_�"/�>W���|˧��|�Gܦ��-)I[�@���v�4h�Z!q쪯�Z�Mȧg���Q�Q;�lcM>O,�q���q�@�@pN�o�v����l�`V�CD��T��R@S\筙+�K������9'k��W�lE�ն�s��rr�_�1�6����ȁ
��z�>� fziR����=`t��g ���m]�$����rަ�S�8D�!�����_��~��uJ�Ksڽ.Ⳳfz0M�/?R�N�+#�.�6&<c]]��ue`�JA���*LB�ě���m���>�)j0<}gg�B�X���z���@�o�X4N�Q;��t��Ӗuͥ��&�0���0�Q�4����8��b�Rz�vZ5;��D ����͖=����,��/�W�O��ñ���ͪ���m��9�����&=�ܗ�4FZ��u|�sLfMW�?e7�1�w��J�<9�04ap	�EU�wZL�0�%���9=������Y�#K��c����_���+��5�G�����R)�:1��B}^���~��)xx�y��VQ�8�Ns���"Eng
0c|]/�ӥY�?&������[sM@�Ba�� )kˎ�R�C1�=� F�x|:�8Ȏo���cq���(T蒶��w'B�n*�Jn��^R�;��酣	�ͦ8�ʳ��J�2'x~��d�0nR�Jq}����z,6U��g�(7����]J����v��%���m<�`���N��)��nd@��;��-Y�5��v^I�M�7�X�0���EcC��;>� ���w�^Թ��~ �m�����w�W�&i�- ��&j�1���s{���5�f��@fJŊ��~��6"`76��>uB*� È�u")����7�� ��b9�=�z��p�ha]���I4z��������jb�_���/��Cb���xI*+igRهs�-�&w� q��7*�L�:K��;k�|�ި��w@}D;�4~H��ѹ�����;�BB�s<���g�LdZ-����+��N�Th�.�2y՟�S18@������&�U��7h�0�	y���+�ߘS)��4�H��b.��xYI|[rN�k���F�U�v�/|k��j�P���m���z�F^��}빦� 	�w�k��,?g�8��!H��=���s~���g��x�J�f����d-��Z���KV�B��P
~s`��-[�	.��c%wڼ���ۦq_j�J�6�hX�J��v-�}5y�Y�J����A��k��ol��:����_�7�ҀA���q�5����V12������U�fs.91¸����C�1��٪:R��K�cyk�)�.�2�8S��1ɔ	�ZR4�;�+�{#y�rl��{�W�zO�Ux|���r�E)��lrv�F-�0g�����c[_z�c0�Q��h���:cCLχsJQl�g�^��A��AP���{��[����V0ԩ�tgP�2~�M-���D���P�(�����~�%T^�S�9����%�ﴱ�����4���=΍�J��*g%&(3)��z�ƶ���ÖS�:8Cq����*�t��Ҥ��;Fu]u�����0�Q|��p�1Y���"���)�cX�(����,9�y�@"In�Z�<�,��%�f�����(�?�fڔ�Bބ%�x�9�<��c����˪˟���� ׹gĐ��,J�����||�2p�;`�w�㭷Q0	t��U�0��2���l�t�|D����_��v�rW�ω!�߄K�B�4��������A���t-D_>	��i��Ye�2#^�V�ø�׊�L-�gZ�+����7=����WG�ݾ��\��(x�?��	2Y>3Gy��y�~u&d�(j�5����te{`k��uFJ�-���j��s��j�M��;�d�����/�V|������Q���B^O�T�"�)�2�s���:wz�Ev2w0[��7,
��;xl��J�1F�?��AL�3�'&�N;����/t�ۤ��[�1����x/��e��5�¬}�r��9yƀ&娄H�>b�äV�R?�MPe������!P���/�d_y�Y�'k��HxEz�㺴�X�IY��|�	;e�W��n:.!�f7'����\l2����O�'����|�pi�Sf�!�BT�VE��n�:)� ��q��В��+��Tf�j<9H�rܲ[:�?�*�UH���邳{g�$+a� ���k����!dyL�#��
���'�Hn��R�g2�t��H���E�Z�CRm����mj��e�܃����[$@�YL��3e��>��d&1������$�T;�>��i��]���_��O�I;�f�^��olۭ����q��w��â?a��r�ٵ@r���/�kW������wk%]����q��A�3�Q"Ϭ�[�V+��I$��O���c`����t�,h�-�L6
�T+{�������wJ ��\h���6|L�ѠI'��@x,�ڂ�U�(	$`��|�x��ӥpf�f����a:�(8�`�
�C��@q!�۾
�����(~ H���̖�ѱ�X.�g8א�~�RP
r䑭���y�a�b��q���8����^����V��HkG����
i?7`8���)��:��+���[y�5�A�X=���F���E��Y�5�b���ǂ��v���;|����W���}�&�%%�����	g���?tIYs�4ޔ�����#��:�)m\�/FѶ�œ�
!��R�ߤʌi��+�,�x���k�g�4�O1��eh�[��.�Q)Ʃ�2��:�S�����&���,�U��Y#�B~`�2�Ƨ�Y8��G�����8Z��>��S3<�/6O�Q�{b[��S�d�l_�o8?$����X-@-g�VS�,��Ԣ[��b�Z���O�P�i��/~3Z�Ui�l'�Z��?'��*ѶxO~O.-M�Q�]���ӝ�.{q�i��)B"�ͨ(���Y��pQ~���`#�.��6\��k��U;���Wm�A|����3�LL�x ���ǔ�*��y���B(��!��^6
�u���Cޤ�����D��	��#�&�C%�._
����
���V�R^�Di"�q �6��+u3�Y���9{虷Bp�x���(]���S�:Y�6��3������ ����4�x�O�`�E���u�6~*@0A!�
j��D}�#��R\���|.$k؏1�t�P4�x�J��Ź���ȹC�Kո�h	�xX)�iBE8v�Z�HÖ��6�G��aqU�I����@x��p:�w��| =�bS���R´n����jY���̝��*���a�$3c^F���&��ݚ��3�ZB��y�6��M�X��t���Eӥk?�7��ɢs�"K�uy��%�2#�n���f��f(KQ�0�+� �;���V�������G>����]b?��s�~d�uH��1w`t�7�Z�����}�s�iΟ�-��`:��gv�E��|����4ޫ��=��+=u����>��(�P�>��x{S"��c�t��')����	�����ա����O�tR{,�Z@�1�R4��m�L�({g.i��c)�/���^�����+a ��Kd����{Ý[���类V^gK�I�&bW����2P)�'�V�&��46�10��Μ�$�T~So�L7	����ٯ��u߬��/G�lRa
V;��Dy�Q_"Q�=&=�4SP�'&i"9�.NT����Vͩ1B&��z�>j�:A�lTCdj�߯ߞq뗬��{]�\a���|m�v�d��&�ـN~\C:u�{9���/�*��H���:0��h�1֫�F.�9ٙWR��؅��Ĩ���A��rC���kW�׮��4�6�8W`�"��1�Y�����׿2`k����\��ܳ 4b���%m`r.�P+G"�ds4�>�y05�_!�lLtG멜xAP���ET�f��ѐC��?���H��]� ��O��_�(�sY��7~����Қ-�P�E�^��v_�3�:��=E^�^�c�]C�����/2Se)|�r� |��^��.��{m�6�-�J������:�#� �]��v���R����mY.C*> �rXNK��E�Sm��l����Q�P�3 ���D~o%�����4���N=�+��֣
JX��L�#�|[s��1W|��bBt�Rh�֝�C�[6�ؠ�O�aAn��팥4![y;����L\�e�b^J󧥇�M��ʥj��~#U�q�0�Or:��!p�<���#��x�\0��R��7�4C����^F�h����_��CG���Dm6���A�X�'��i���L���U�L�	u�0�Ew[�2�v��_&Uq
4>4i���np�M,_(<��~-� |�Ӵ�4������$M�����l]
�*��V�訁�z�<M::IE�'WA�x�$�u��z&������7��|�n��5��Q���E6���XT��F�ޘ����&?�#���R��Zm�!fQ>��p�����?�lX��/���8 ��/a��}���iV09�+�|�Fw��h���7��
%�5��;� �@�7l�	5��Ei�J�;�,?ҡ�9����A�kڝ 4�MP��N��{O�'�-ʪ�6�O�ZxҶ�3y~rӏ��J���-�[4^P}z}C��\|}<�߷A��%�+e5���Z\�ïqV�L15�Ӟ57�`�w���M���[�Ep�O?��g��2�+&"�,'Jrϵ���&��!Y�75��R���Q��ѮA{�{*���_���b�l �odV��<O�L���c���]���`]bS�36�d#��H��g��*/����(Kڛxځ̓^��ЊNh3"�[�k����a��i�#�C��b)>�&|��H>���qd�T>z���6[E�tθbA�s�A�s��?�K�G �T�lQ��S]x}�%�����.��1d��m+�EGcW��P?�Yy�K`����?qm]��6�����_1&q��ca���>'E�T�5;s4q��0����~-�2�^=���j`�ۨ�� �E��/'ϙ.�t�zT��G�J�]|((/�w�~�:0��J_3oQ���5?3�������ꧦCwZ��;�ɷ=��G:��ԏ��_�Xw� ���Jѫ���{b�I�H�q\�t�:A+4�Uu4Ɍ�2�D�n$���}F�4xﲥ�;��Q����A��}j������`X�Y,�۩�궈Թb&���nv7y\�����ϚF��n�yŨ��q�4rV���$&������8�>��$��-[p6�ϳ5�*�%�O�Y��C�!5�aPX6�pj6�'�!_�E���	���C���ds�>�3� XčY#� �U+����Y&�];����o�ٷ %�q>�Pcv����X�̶h�����u�HD�LK��B����WѸ�7:B7�l���swI���ݼ�h��I۷!�p��G}�C���ҝ���u��<��8T�5*���I�5,6���!RL���k��5�&+
��f��	z���	�C��������`�ee�LAE�s�@EM��oJ�h�R�"g�F�Q�PEK�3΀�&C!�9��1z�$�i^���72�mb����Ϯ���Pl�~h��<�֙wA�B?ߋ�__[���&�U�_E��b�{Ge���`Nۓo��-�� L4M�p6pH9!�	��1E��O��.�t��M|�Ds �v2$�ǚ�h[x�g��f822ʢi�7�!9��	&��΋q��(6��$�k<	05�5�ݔ��r��_�O��\������&w׫|ڑ��^�P�*�X>�&�Y�
C?<cǝm3���C:�E�����#��UI�����\3bU���X,[?/��s�5C �fG�� ^h=T_�6���``y?��K�y
��!Vba��$���Cղ>�E�F�e�=P�c�!�劖�D�_
ʈi����9��	�X��f]�^^=�w��B�k�`��7���T$ь6�_�z{"g��5��2��f�V�HI}��xmO��m/]�O�B3L��x:g�ݎ����t{�"��ڽ�5?�[l��{�Et��͋���h������5���a�F��3�E����)1����%�?�#�S`L9����ul�`1�c��	8	���x�K�:����4I�U[$G�Μe�3p�� l�\e��*KX/K�K?�}����4�����B�DTӮ�����Zc��/Ν�4����SJ`��"^�j�l�W����إ�=��`\}L�O�;���Z�c����SP�=��[��}�i����d˟�Xi1)Ut��������[:�ח-�AB�8tY�;�����2l/P�i������9��[��u�r�$��ZU��F�4�����0�&�����x0&��3z�������΂2��F 6פN�2)E��5g~�f�Hx	E���^�����G���g���t��R���0K͈����8��ܲE�J��~������v���s�o'�����m0�+�����D#Uz�z$�����5�Ad��&|W,A�f��QK	 7��}E�oK���6|��]�	 UtTF��o��':fD�(t:�R��c�P\��`�ғ`��e���-�7?��`p#3S[����}�*KF*�$�8z�)��m��>����eh�4�@��"�K�\_�̓�Ѷ�s$� ���[�t���}{ʇ̞�������J�ֿ��H���:��7i�.���sh�Xj:��n�8��Z��#l#�
������cr5�ͺ9 
�!���w��D��D,�?ݗ-c����N�R��wk���z�"++R,��,�C�Q�L \{uڕ&vWG�(�~B�{��?R6ٿ+^ґƈ���d~v�v���"�"��,�b��N]�S��f�D`�@ڏ�����wr�s})m�P��昸��@�>��6�6%6�����_�z�3���[M�c����`ķ���6�jo5����uD"g ��+!��B�Б�}���c!.K����/7ԫٸ�N���?o�19�;'&~XRޔ����u�a,����i��\ u8�-��Axz���=	��]|轚�'�3QC�o�^X�s��/�P/(��� >�_���SrT���^���`\S]�S�i������lۗ�Q� �Nl�#��e�����L����8()i�Ia� 3.ُA��_ [�����av��/�|�E��JN��T�6����~8X�d���G��ɓ��wq�T��+½W:�}��(\�І�F:�ʚ�Y�mRm�p���w�7�)E��%����Μ+t-�(���D5ξd�ڽw��`, J\��l�ǓgݗV�i�(��>pI���߉WOxޅ�Ǭ2�Pp�$����ݙ��d�x�	M�Jp(+V(�>�{��dS2�\�
u�v���={&j��bq�n��7�y�B��M��N	�U-b��Π�q0��?q3�i?�u/Qf*��U�ٝ��uc#�����$�O [��hߺH9Vt�\��_�K�5T.Ea�P۔��չY��^��@�$��wA�+l��ۭ;ͮ��C)�zb�n�y.ɯ|��"L��_"��l�(|"�F�';9U?�ՙ��r��e)O�ċ���+�����l������ \��j!����U��@�)c��vzʃ%D�vU� f���-���^5� ����|�Ɉ�j��:�����:����%�D��ھ��@��?��ZYbR>b�胭��G�$҇������lu�U��
,;���ϱ�;w  tA�k_|�\@�I�S�"eU��d�zZ>���n��y�$�] ����`I詾�I5*y���3A[׀�a��~&zՒ�U��Qn<t��o��s=�&]\�o_��ij���g�i�oS3�\m�T}��������a����֔"���۶hLޱ��^�m�8x�@ ߘ����L���D�7I����.���R�Wɨzn���E��^.bL��z�q>���"��9��/�S�4���Lh�=�b�8	�c���3�C��C��Wq�R�Uj�����@M]���ig��j��G�}U��EP������.�UF��2�D�(-��h�ͯ��� ��T�`������Z>�1P���aZܜ��&ދ�)��0�ƕA�� %�����c�Vf+sWi�m�h��I�k\��A��F�D��G����Qq�������:��*��f��݊8��YXW�O��m"W/��\Y|�#;M�O>p0ņ�br��{�au��BfFr��3m��S��3�ً{!xd�Z��eF��E�=��s�d��V��2����Ŗ|������b&���+�#x�M�j�R��|\��O�s�T\�8��q� �E2�3~"4�%v��Aި����
��7X`��@QW7�(��&9ʑτd2��M&�p�~k���&�&N��2��W�ߠ����\k2���z���:j!]�*/�E��S�{��E`�T��eѯ������=ˑ?����4�Os�Z�+���N\\��NkAfH��JԺ�j�I�f�D�(}9��yf]�DC��7�s� Գ�]d���5�I�@�p��zW��� B�B"�t���ګ��'�D�z�È4�a�?#�R�̩�oL�.��/��ȵB��e���Fӧ[��Ÿ�:��E5V�SCGHhZ
]��9�r�M����.��10��3�w 6a�<���� ���_���h=�`1�f]�q� ��gm����3�rDv�=䓿z���j7�:/�Z��Q��N���E�-�,ғG�	�"��ï�{����7�<��s�c��@�Wh}����H�UB���?��t�$�t�r���!���/rnPV���FN� ���_�^8�Y%����7��I�ĉ��J�9� �ɕ@"c�ͣ�R�CVMmjg;2������T~�t�=yЩk�j�Eivt�������W�_N�*��F̆��xo9;H�H�A�8���o���*����%�t�::�rV�Pl�Ӽ��dg)>�E�[y²P�a�Rd2|��p���Ղ�FO:L��w[e}\?�s���r9t�7���i��S�=�������ן��a�(���[G^��J�f��F{s������4k-�zU�����t�v��]�0�<���T��ŏ�����<�Rx��JQ�@��F��O�]����V��y7��fg{�ϖ�S>ʄ�	Q���\zR#K'2Fe��F[V��);oC�y�,ƭQAJ����ǚ���H�;���*�~rM\��z�"�_:=$��^,˜хn3T�t��;NJ�xi8,r�m��9z{ah���D����
3�C~vK��K����w������e�2�����MH]��9������c��N�P��L2au�tݍт�������� �����\��ﷶ6m�,��q�WB��k=fmQZ���.�m#�F����:��i�7���uzs�SH��,~�
��}O�5ρ<V9�Dw5��R�� ��M�U*,V����p�*���j�z_�蓀+���:�l&�z���/����� JsJ�a��(�`��<Xݎ�X��'��A�z��1$�w�~��/̙|3}q\��" �p5�X�v�Yʠ���6ʴ�f�J{.��b�(���֦�7�O��bխ��E�6 ����I����a���S�w��ee��9�0ae ��2����}��&�<Fe._�uwOdC;�L��%q���۹�mk��r6��,�m���n�oݖ�q�k�d-��ZuQ�o�>p����G����f
i�p��b���!�8����˷^��E�?��B �s��Mz��r1�={7����^��O�G{�X6C���������GO�w�a�2;+_�g{��q�Y�.��Ʃ"�� �ߨ|<l`
�b6����5E;���B㒂3n�i��v�;��AW�:�S�H�\�'w�=P0�d���r۟�(�d��~o�9[�om��%8�am��gg͵�S���MԃqG�G 8L<W/9�vl�6�T�EG���oOK}=�[��6ja\z���A-�ǟ�+��q��b&�/J�S �� ���
�/�a&���>�x����,��5�ꐱQX�[gSvZ��Ƈ�؆�I��$��ݫ�6�f�t�ؠ���� z�����u�P�q0Ns�W�kŅ��8����Kv���`�? w�GL
(��C�X��+Z�c���(j͞�r+�|ÿ�x��2L)q��^`h=��8?_����P1����5%���x�k�̵�Max
1*��!�id�)�Y5�D�pr�JF*u�g�a������l+�c}U����=������31�`�"
*g[�U!TS��g$���M�{g�'�o�;���e�]��6vͼ2��$l�p]8'���F	gz��f�3h��^v�]8�/s�v�SR	�JKQ���6���Q(EG[����W�n���E\���1y/m%�V!�=�?Q�Nӕ��7U��.��$걢y�a%�a����l����N��deP�"�\���5�u��1h�����a��~��ț�.⒢q{'����?9=� ����% ��MtTq�(W�����ip�J�S��ձ_1V���m�d2謽����!v�L�G�=]�o��b�f0�Lu<�����0^S�7(�Eȥ�m�X�����ms��25S���i�8Sv�_�C`5;(E��"W#�`�Z�8e��Ī�'>���cW�����u̘V��,t�d�k��!4��ċ�vLN�"liR�H��g�I)��ӛͦ:�@�=f_�����k?[���w
ܷ,Gx����:��]Ϭ7���\9�c9��d�x@���x��v�6�CAk�S��]}��"v�VR�;x��n,�?��79ڸp�E)�a��B��4���5"�l\�����K-���8$���o�ឆ#T�3�	�.���?4y�$�ZP#R�������M��d�)�[ƴ�D�N���0�W�e�� ��a1����eF�w����6��(]�ۗj%�[`�:a)-��u���v.�:"+�1(=NO-�L�yO�y���w���n�,��K)����c�0�-��cF/	���ur�hJ�⻸]�����@J�N�RòEh)��I�Q�92�[������,��C�A>Y�$����R#ʱ��r;�ɼW7^��,��?�%a�����f"'� NS�A�˚�x`�|���R7���L���u�7��z�Ԅ�C���`^��##��e��=,��oU���k3���1��~���w�0�	-|���wW������̚��F��L.�pZ�*�_����OJ�7�G�0e����jA��:�0<�9a�%��4�\�=�Yt��Wը���a���hr�!	*>�i���4��p.bm��(d�l����������XI��X���`�ǰ�f1^!��c1Έ0��m��J"�,��_�����k��VmE@��cdtݲ��N��6���7v�4k$�Ύ�d�ӵ��p z<��YP�!r�Uw�����7�GCbxRh�@��DRm�q2��vD[L|�Yd�,$�lO�*���J��Ӂ�A��=��H��N�F��X4M���ph��E�]�9�d���$j�9|�`�4-HP��@��+�-r2�wElY���Q�yd�c�g���}eBm��gQ/%zo4x;�D+>�p�T｢2NцPŸ"���c�*���@�+��� �͝��5Js��d���a
{�XN�t�jc�<�Ss�r�D8RG���m5�^�8���lˊI��"��:{c� \ bǬ�S�|�П����@�+[o�;�Ӱڣ��:�֜l	
u��� �I%��{���I�Ѫu�+���M/�/�?/���|9��=��M�����b�̍6��^��Af��pq|,R\&��p����k��O*5A�!K�E����0������ ᱙pU�l��E>�!]S�`�;�����j-9���$�5	�忷>9@���
3��5�(+�?�������Yg���� �!��.� 	�ƉΝ�t�W���Z���}��C���4g�ܡ^��g_�[�Q�&F�����'C����#(`�^��:��r�A�l��`�;�Y��(�om�2i�;cI�������.]�c�+~�E=��]f��5:�T�y�Q��Y��Ɔ�M�K��^�#*r	����{?`�_)^����6�YȒ��1Sd�����6��4�_s"�ݗW/io(��;������Ws��u<|ﾼ��<��ŧ;/4m4�L�ڣ68K�X���9��W�Z8����i�V�;�1��%�9ʤE|
��3J�mY��t%�͐��x�_���@U�\p�ٳW*�$�tW"�c?���]��q��󚍪%b1�bZ�,��k����	�K�����@/��o�``�����1��۲���v�re(��	?��L�&�~�*T�;�B�vh�7���qU�=l��y'_{�ׄ^��v�n{�n<c�?��n��S�&V�����B���s+�T_+H�N�4lV����gӥ�h.a۾�9F����o�Jƹ�r� ,��V�CY&�bZ{E�<�[`K����v�@G�gKlIQV��.{�8M����±��L���H����U�}���?�����a���$���3 �f������0�o�_cx������Q( ������D���-�� �o�+H���/�y���k�l>��bXE�F�"Pi1�����7�_�Y`���^G�����������1l�kz�e\A�!)�c�M��P�x{{�zh�)�';�m�i	�.@���Kz�BeE�jk
1J��Նg!�8�̦��GI/X��⊨yڣl�]�%��N$e'�'N׫�,��Ì�S�в#2?\�Mbm]<�x�Y�l���gąu��6��#�}�=�]�b4�#�2��LZN�)�LI���m�M`x�H���n��I �mupR�v���o:��.y+�)�����I���8M��{��݃y�2��Q`��>Er³�e��-H$1�%Ѻ7���k>��W
þ��mg���z�	F��k4E	^�m��sj�RAJ#�������;-�1{e���E)�S��3r461[�cw�g{g6ee��4� S��į^\С$�*]#O�� �����z1Hѧl����3�#��~�ox�{��"h�������X�@�P��f�\���QZv.U�XW [��jd?�T���'
��5{���� �eO������7���x���0�q�	�ة�؎�����w���fO��aH��}�'(�<��cD2���+�w����ˌ��6�'b�ңo�d-� c�S�@_���9u���.�Ś��I�mTG�u�Au�C�>���yH*��^f��v��_�C����1���g�� k�UX�$�ĻX�=�-㿮Ѱ�:ȗ��Y���/z�f&"�Q�T�AsA]�D�	&q�a�&J8����먟Y�DOo�%��eI�H�)����E�:ޡ:=�n���JL�1`�D��E��ٛ(ic���D�;���7?�Nn�%`{&���g�wCmq5Ό(Ž@Y�0�e������ۉ���M�j슸�ASi ���?�]�|���W����y�P�k�4y?q�K�F�q����3��#I���5��2}��v�i��42Q�x��N"+=�n�~mt�0��p�(�NEGN���������3��ʰH��$�p�]���� +q;y@����z�	�Z�QtVǓ=���c��S�}z�7j����1mn���d*?�����[�����۝����	R�$V&\���z�R+��X�X�<v��� ��r\I�!�6��,?Zȃ@�gj5oJ��a�9H�i�7��%����Ԧ��`�Y����WI���p&3�}�Ԇj�\vj�?���(��:�L�1�lx���V���я�W0��@i]8��냓�G��}��k�/��<qjc�Ŏ�VV|�=f�����>+�§�	ZT�����,�а���z�=Q�ܶǧO�jΗE�gR�m(��[7Y4��.�.8m�Il��?�n	^��o&7�E��l�&����{ش��lo��N�u�[�C�c�W$�{/������*��O�S��-�2Fh���0�Ӳ#ǆ�����d��iY/�I,��k>�R�Vf���}�Q�
�,k�L��,N��{Ъ�ݴxZY:�l�Pr�5P���쵂����\���N���b�{���!҂����ᩮR�tFd��9$�9y�I���X�3<��\I���'�H�x��}]�B��$;ʨrE�?��'<i�nl
sѴ���.av�>ky�O���S���Z�E��gg����e�j�د~ �5���W�P�2�+���B5�h���|���aJ��dӷ%����o�o�8Q��"̴6|2:�e�	���.	u��G��p@lu�p{ƹS|���7�!�[��~ ���DٲE�D��zD��B���J�j���Nsj����-#��j�'*B�f[/���6!UZj�5��ѫ}l��o�בn_��`L�.Xݯ��tva�@���+(�q��3,����_����a��|�Տ���|&��Q,\Bq�y��U�sA�J����\ID�wUeb����B��l+����=/J.���)��zZV��?e�;�3���I@$H�FQi�?�)�d2N�3��O�aa�_�>g���%����č�tkl
��;e����^~��+�\��h��F$�Wң��T��˧l�\n�8C�X|ާP*Z��7贃#��A��;�3hi��\K��$��y��h��?�mؤز/ws%�~��+�� 
���ۇ�C<��%��5���W5.�G���*N!-Vc4�d[�S���Otdǽݷȧթ���Ю#�4|�eQ���2V�P��'2�É�@X`�;���`�+R�-��R9��=�����X��]�o{9$e~��?��&����d*9��*5	!�D�U3����[Ґ��q3��/�>�g}�2���n���}���Ǜ�CFZ_����^Px\��^Dm0g�@�\d/ �!y��n�}Ws$CcB��e��QO᪼Òf�՞6�O���OQ0�������e'#3��6��ɹ=�KKR��i�`ahe��G{P�h��-qܑ�����J������	B�� ���E��_/aKtu��z'�S�Kk	ϯ��M�����J�O3��XDK?���cw:�FN�C*�`\���{ynOz����.g,���3ɑ��X��[�O��p%�U;yn��I����I:�d��4I Gw��<�s���ٲ�;�D.�-��[Mi)��.���h鞧�Ƙc�gO
sM]!��6�+����܍����@�6Yk�E#)�0(�I���5ځ��Z�5}^�Ihq<H|v�EmUm�1�Ud�Tw�i��1@Ε�I|��ǹ�{{9)� N�>���Q3����УV��[��3
�r�f�앸���<oM����y����+��"����j���J���w���d��^�:���R_ޜiʔC'4�"�Smc�'�� ���+����/��Ӛ���6oMP��uW^x�b>u+�,M;��>�ca�����������2��9��k���#m�B��L�-��~-�eP�����{
	��{�<t�� �R\�&�^�=q�O���-hz�I^���4v�O��3����zq9�o?�ۦ^5���M��=��^g?Vf�!�k��)���k�߫a��P�6��(MTv�l��H��/Jޚ��$bҁWs�n��I��x�Ͻ�*D���՛jz�RIf."9�mS�� �yή�_�������/�Ϳ�����!�|���?[�]��P`َ}G�z.i\�	$0GP����}:���i���-}���x��JX�栉�i"=H���M��u���Z�����w�X]�R�d5c���FK4u$m¶~"������A"�ǅ��6T���D�fr߼�v￝>n��}�	Ta@�7)�b�!��u�!���Y��˰�݅�r]��yQ��d�A�մ����:�
�lϊ��$W����a:E/R���y��wk_�T>�}<��=OD^���p�֒�L���$�aE��Z�"�I�}��=OhAZ�2��\핂l0>�S]�5�UW.�c�IB�3o�j��#��h�&Z�v&��@�I]�&[�xi�(]�:�d��>���I��[���_�ෝpU�B�}�Du���$�?�+���:��32?��Ε	X�B�C�x��U{p��)4���xl6�����L�S��� x6X�~��cS%�F�E��÷`n5�v�F�cP?,4aVp��&�p��?P�£���r~���+p�$�w��N����d�
d~֧����ܟ6Q"��i>��+>MV��8最�W�0�q��~�s;��7F��g�ar�*�-��F~k۫ڤX�Z�ƙ���ʎ<�t��o�[�{��7�/J�f�o!��Õ@��4G���� �3l�Tːh�Vj}���9�KSs����kB(��gy�`Q������R��C�r kuaA?(��	~å����)�I�$���(0W������C)_B��6Y&Τ���ϖ:�
Ɏrm��`_��I�뜕G��0�"3��.�\s��%O�|���9U#���rR!8 W�G��1�_�����GQ���8F5����Ci�o��B���%���M���0���ؘ֦����p���2%?��龫�&�e�nIB��Ѐc�Ӵ�Fb�i:����2������:�H6��
y^�)�f��O�ֳs�Ar�RU
���Q���S��|2�Zv����M6u*z�>�v�R^=��g6��F
q4z�a�m�èT��-.M�Mjʔ��@�۪\Z��L��.3�E:��Z ��R�ל��l�C�Y�I)�U��㡄zn��gw�W�X� ��>����v+���I�9
7�r�|Ʋas����Ӻ��Y6�5�4��cͦ�^��9(�����/�=K���=}�-XOFv�U�ZD� �Ĥ=y�7̭Bf+X�*�����A�Ù�):�������6ɱ0|P]�-N�{�f崪�j�M�񊁍� ���
;��ΞL9�&O>5N�Q��W'ee!��nw����TmSn��� ]Y3�O�J��u����z;6��Vd��D�����N;�i?Q�F�����$���tt�"��J�K�m�@Q}��F�^�#����J�����V���d�GQ04���ǓGM�jЖ�?й���jj/�JR�.�oI�����6�Rt��1M ��n������%�k������UQ�̲�>�?��t�7�������@W*bԼ7�vd����%؄0�L�E����A_>��v�
.aGO�f����q���9̅�����0N_��R��L��.Ǒe6���dd���͔�p�tZJOGs����luvڟ��Gu�A����A.lO�ߓН;�.(�Y�"�I�_�����g����ᇧ[1�3]�����`��l�sE��]#ڷ�&������Iz9<#:oI����g� ̄����`m��F3�/�q�fR|�`���L�q;G�)�c�[�	��z�zڱ� �E�`��H���(��!I�e������o�am6K�a;$	_���a���SDu�;ʸ=/6 �/Ti=y�	X��'�皨^�'�s)=~�r{:kJh��`/�I< �b�% A�\c40�u���n��j=�2�!���)?z~lr1T�����%� n�3�m_�/�ǷjA�S%|��i�<��7���8�E�����/�	����w���2�Vcǟ-�p��xrlᠠ�+w�5��t��58���q]�w��O~�\�ǐ ,��ת9j�ĺw�.˭A+�A��U')Ȁ�nWf�EN�*�fɨR�(1�T�:�3�����d��=�����U�~�E�'�I�*븆��t�Y����*5�E��Ȱ���T��s��������I�4��;V0{�Ќ�rIL�ٍ9\|���<���������/��,$�:u0)�hD�0��Q=�}B��Ǉi聪0����W�6��a��.�0��v@����򳙞�����)l/��c�K�S��U���Ld72�}�4o~� �gT�I�FP�x�P�6�a���}����	�(��z35)v�y�s�/�l�|��2nk�tF�5�C�j+4�p��+�W��֐���j:�7#Ƞ$Z��%�o�=��26%�e�:��7^/�Y1�z��_���t����n����FEQթ_�i9��%��a�gE?ȏ=�]/xC>� ��iȎk�+����pd�$J�yB�7�X;N5�2�����uE�����E���-�O���| �6A������f�B�2�4n[EM���M���U?IL)�KU�ˬi$��>���^W�5��o�z����-� �8��I����QĤ���U*_�pc�d;-$W�W���v*�O�S˃[%�� �k�)�n�CSE���s>ٍ�y���o�����ۆx���Alp3W%���in��Cp�I����x���@�ӵ�d\ .|4w�V�
�.�9K���i2S����tD�
j->��Ǎ x�2�l�xM;���JC^�=ls<OY��v���_���ycG� N)nK��r\�:� ���#�����h����z�}�0h�����:���.;.�?
�����L�X}0����C
�S�����u���4޺����T�\ꌂ����g�z�����.�͹9�1�ou�-�J�*���EI���O�;�L�
��#Zl�!)p�ޅ^��}w����N�VA@i��Ta�+�ʢ�-����1��+*��L,PM_���-j��|H�C��epRa ��syU聚�� ��fIU������Z�������딵:Aik����~�a�m���ϙھ6Lu|�!H�/M��~]UK6h��ng��;гS�*�"@-�Y����`葒�d������V�@()�7�j�_�N�仕Z��N/�72�XѕV^�˔������h���{Je�o�r�B�H�IGG��;�:��r-���R����mդZ⃔���^	������S�<�:�]3���9����x���J�rIB��K^��p��&q��i�����飤Oj�k&}Ҽjt�T@�	U:�8���z1��aM|0��"ġ��7J ���Q��=�L+m���Ar�蕸�B?�����A�K��_��U43��_=Z�Q�x@}��մMO�H-��#�@�+E�$�/��{F��ӝ��S��,��cfLT����\��{MH�) ]:Jch�*���b�#RMN[�B��p������I�.E��ch%��\f}��`��8D��/�J������̕9���� .��M5@͠O�pA�l��O[3�	D3Csާ
'#둎�S�`��`�v�����TOjd��u%!|�M��ů[kR����a_f�I��̢x/W�$˷ާi��wOY��@IjtO	ӹSk';_����#,'��.��S��k���f}|=�?PE�H������>��Yݎ`)$�%n�"�$�S��J�����9�E�{~R��=��Dpz*�f:�հ�ȟ#&ٗ܍M�E|��)�������ϼ3��Q�;�����5Ĕ{t����cn����yh��
א?#�jSzSs��wvުq/hv��!�ս];�ZxƷ.&��)d������~f�>/VeA�.SDܕ�
-�܀+��/�@����p�P8����ٞ��b�ы��fc9P���x�⟤�j�@�Te�� \�r�Mx`��&n+w��0���zH���K���ҦAO�#+槒g�;B������Ŋ�6[�=c��\|���$y�X=��; ˭(�@2��[[�z��E��
��z�@�Vc��T�+E�� ��V?�(��%�֋}�c+K]�c�.5d�uj}�f ��gF
S�Y�u؊��*f�V^�Cձ����<LGu�[a������zΘ�WE<�#]rB.m, �
��˯�ѪYg�ƛ��~�[���X5$d�����R�?6>/�9'��\����>g�0���&�>G1�<�$�,oNkǳ�ɋ��e��5�}R�$s?$5+�P���Ƅ��T���qNԾ:n%I�^������M|�&���O{X��M��r��7KQ"�ş�Ұ��,Ͳ���|��ޱ�S�M�wը�u����_�e|�x��7�8N/�o��]n����B�X�@߱צ�� ��b�qͪdF�L셄Ё�| 9�������Ų^�h�k�^���
V�:�\xcQ�g�	��T� �ny?�j0ʅX���j�Ok�7[pBݫ��Z��yS_b��o�ߞ(c��jc	��H'�v��j���� C+�P^��G��
�%��I!G�-4�iP-#7������A-M��n/�5M��['�$_�p-����"��]ȍO2�gӶE�h���¥�W^�4�����
�'`����m ���A5n��t���(���"R �Cw%T�1S���\U�����c*��U��k���wla:���4>3�ŀ������̡��5YiQ�����wT��v��Y����������L�p5�y8�=���:)�Ny@���׏��9�;OlS�f�-T��᱗�_�&��u�u�~�Ua�g��t3ZVn�Mh����5rz)������FaP#��B#���h�,>���rwPū`r����N�����)?�Õ��Y��'��w�3���f�љ^�q�Bo|/�N������ޘS���+�a#���LE`�A{W+#���� �_j}ja3��!#���ı4�Y�<�ڇ��|Z����ӥr�`�;>��D�4�Ų[����L6y����N�`�ȊU�����}��ٙx�z��*���i��2 �* .=�`��I����1�\����9c�b��kXԵ�&٭�Ͼ�*[��3�MB�!��-T��
Ҍ|�����[saR�r�%㑞��m��֒����N�φ�V��k�B��ǿW>F.�#$B
9n��)�7�A��P�B�G�P#�;߇92��ͅ���PeH4�Ϝ���W_y�_��)�u�8.U��K���bn8a̟`���z���=���`	�@�����@���;�A�ת��Ӎ���imG��p+#�9��S�Z�B���i��2B���nˍ�p���+U�(����O@[M�H� ��J.�!�L_cf�^�3�_��
��1~�[@�%�Y�e�зh`:R�[�b�M��� �������Y�hh�]�ɟ��7�� ��gؓO�m� RT�p爏B���Z.�N.A�˨1+j���>MW�kt��U����X�-���Ԯ�%�۹\fa�Ͷ6Z!,M=⻷��MqBh����H}��-�\X*4�����c�Y�y�����Q�#�C���2R�eO���e<�b.�,$�R{9"�+(���W�,��E�GQ4:,W��\�#�x;� ��ɊC���G�gmlqc��6��|�����>���ff�����߹X/J�P!�Ic�Ӭ������:֗y�5~�Em�	�mm;�5�^X����b�[��e|H��:��R�a��b��Ftr�Y�����erJ�N� �8gqf"D��_IL#d
��N��FZ����?~�=%ua@��&���:�����v��[�i�/�;�l��  :&F] ��`(�i���e����U�YA̼F�rF���'�ׇ�"��DH�'��V���_3��9uݒ�K*	����ͥ�����I�˨ŗ6[�¡�3���,|l�)vIwC���n]��Rq_������tկ�<e婦�Z��b���Ɗ�"7oU�S<�f�<�G����3�#�ͷ�Kb
�$eb��x����KQX��;��p���Q�/�B�=^���R����cd\������|b��m䯀��b.h�rWM�����h�o!�`�)���>W؇<�>�T�BKu1��5�MK���DWb�?Z$� _`PY�z�4�حn.ً�c{�����+;��c}�nVʴ��޵f���i�9���~�,��G���m�����+Bީ$p�'/�C㽭G��F��7�O�s��u,�6a�R5���T^|UsS�c�7�x�I��e��=t�q#��2��1��*oz�̼"��*���m*�����/XSUb��?}�w���zX`׆9��m=`��~\;�գN�_iw���,:�Q"�I	��28�}c�
B�| ��Ŷ9Z=��%�DܗIT�����P��S��'ȡo��(��O7GC��E�$���h��$n�
��0��s�-:k!|5����O�q�[�s�G��W��,=m:q��l��9��9�]�T�����iN�k*2,9�o�&�Q3���vڄ�wT��.�Տ�vi� a7v
��vI~�U?�S��r4�� '���ߣ\߼hQ�Ŕ�B�djd n}�� �'A�0��R7<g��<��-u�+^� Pp�`ȭw��IV���ޜ���h'3�@t��x�+rK
j�ќ���f"l>�������X���l��H�=C�	<O�OI��=Ƙ*eR"�;7�
����P���|uf�QObWB��v�?wb���no#��9���E����`��]������R깦����t5���L=oD;Z���lC��0��b�~��s	q�`0���~�ܹ��R������.DX<XU@�	Cץ�:����}��vK�1fj�9
%�^���)�1���y����sŚ�0b	^��EosR&�އy\���x����Ձ��ru-����\�H�Ղ�u������/�M�:�&烿��,.O�ӵ�hU(�ӡ�k�;KxHS�?ҏrn���Q����6ɘ��N_�o��J1백�h+�&i(�n�Q����$|3��9c��C��U����S�,n�,��(��_:1zv���яx�'��ҟ��L<!7� "]RE��]����SP��#�ź#V�B���O�3t7�E@$j�G���%,�6[:lC rLǨ_���DW�O��@z�t��LŹڑ�����aȉpN`�)�<r;��~�'r�K�8y�;�{ 6��h��
���{ƛP�&�4�e%�⯇����y����kY���;��PU��8{i��VZ�N�
���k��c���K�Ds���W�v6Ԟ�n� k���8������ ��zr���;2g��f��Rppmu��(/W��:бg�
{2O��2 �%����;M��11Ik���P�������$�S@u;0%\�G�&`^8�V��;�o��\����M�&��r�B�<���6�'$9�Dρ<�/L�X�����O7hi�'��ê����
�~x�,�MbՌ��Џg;����C�K���]
ˉZ�m6�c�������E4�/���,����t��VX�H���A4�� d����K�H�7B�`6]������0*)`�X�z4<Q�\w|]��{��F!���~T_�N�q4g���*9��ǀ��w�>���F.Ķ��eɡ���Bh����.m�υH�O5H�H�㟠	[�����	.���E�~�I3Ƀ"�4���c��!8N��ހ��Dn����Ⱥ����պ7S!Z��; ���e�̂#b�%����]�c�5eX�t04�"�w�L+��"b(k��δm$3�������r5��:�GB���F��l���!7�̵�C26�k�T@�G7��`�\fR#��}X+������P�(�A���k��ih=����Պ�l^z�/�6��V�)(��Z�(�:��^��@v���y/�t�!�^g
�cR+y12w�$bM��N��x�q��f
�zݫv�����Ց�il�yZ�8=l�$�
�tC�:4,�?{>�h����>��WW}�v HEUX�o��0*+&�ñ'g߹�_��G��B���� �-<��ㅇ��۱�R5�ri&��ܝ1�(�P�>��NkԊ��s��O��j�9�B��t�/�D�sz�\~���A����~�k#SՂ��oە'�kÅv�o'��+/��;��!�!��"t��Z��}���e&WBlwu$��O�=.�U<�[(��rb��$�IŐAw-	)����xN�|�M%S>�R��w\�T��hJqWƆ8�l�����P����'Y�	�6�i9��s>ٓ���q%�K��T|�6�v mGr}�DbЙM�ަKK[�pv��fA1�@]�(:�a4��Ki�o"�/0�e���%�Ny�z���sH���d��e��~S�����`n��2(����;Wrވ�nht�L���h�3%����ş�r����<�i�v>����fan�h�]�d1V�%��~���
H5/}�8��'niR3��w�y]\��'<�k���"��S7�߉���)9���\��ɸ�&!�@<ٞ��:'���V�?�2���^�����~f���0nl#3 ��L������(N.� ���)���/�ܶ��B�q����x�\���6nA�� ?Y�͍��'>_+��-����J���kӭ!f돺�P��!�%�}'��L='�	�}cB8��i�{��F�8:-o;��;�;%vx�0rM(������ɠ���Gn1���u��Xp��mH���p��M�B�Z��[*�6m�P���V���s�Y
1��H8\�ȃ�=���G���d����������:��_p���'L��ҜRA�H-��IFG�.�0l��1�=gBc��x��8�ư$�^�15D�U�<��C���{ːV���PԘ4�k�s��`o8Zl�P�x
>8t�P�C��kL. �����z��P�\���M��2$,�8#���e� ^�a����x�@?0Z�Q����n}���.��۫����i#w�e?��)>g"����(��L4����s�-p��s1ٹ*d`��O��a�`���+��3�P���ƈ��Iؒ_�T�bA��i~�����*9���W�����^�7����Zc��1�{ϡ�����r�G�n������p��ޮ���x&�k;^z`tQ�q\��H>GA_�x�t�[�����(ԅ�17q�q�'�X�	��6�9k�)l��A'w�=����T
�e�I'��	xy��5�	8�/�Iܚ̪��H�%ǀ?��-��RǠ���&P���2j�b�H�_��C�Q���OT:RH�#:���3���!o�����bs����W�>���ʵ帱�-���S�xU�`h�#��r|+��<�<9}�&��un��q�zK�<�C�sď�tg�� >��Ѿv�a�v� ������ڙp�G6ӗ���,6�Y�����x-����dU�/*�ao�$��E	�h��ug�;�S�%H�d�l���XG��WQXn�^f���Iqw,`���MhLUH]N��BX5��>]'N{�"f|�[c�Z�N�HX���r����ݠ�ˢ�3��GGV4ܢV' ��P�*~W�w�Ϭ/�0����l�I�xW6I��!�i,ȗD��3B����b?�D"�e~]��['���Dh�s_�r���$��cW�,Dz]{����f�q4i\�'
 �C���|
E����{�����j�$I��6�&FI���ړ����͘�g����Z%���^:�tʸ#,���?���èCE~(��%�QЎh^�ID�H��nW�sR)Ӓk��+�Z��оk�.)�e��F��ӌW�)>!�u�}w�N�㸝��!�z��,��L�\�j�7��H�k�[d�`�9=,<qd+�86��	�iy�ͻH�A����g;_~�×w��®g���5�ΒQI�vâ@��}�f.h�i��g��E>J׆�?�}@W��L���4��8k�j�
��P�X��<�c��Vʚ5���L�!P%3����ykJ\_
CӾ���ĉޡ�N���n���{^�P�P^R�:U�4��ކ��S�Ӱ-oH��c��8�+�鼅���{�d�6���n鹪�0�Ö3쩱~j�dm�Η�X�SvO��fM_�D�u�g.a�6:w�����S��^
ذ��i���?�wsN�����}
��3�+a�Q���,�_�&�i�����Ҋʥ(m0�m�w�F"([M�s��2
��\�('�v�
_��?T1]h�h|���c��N0�$�J�\Ie�ExI-�ܪM6l;��#�sԒ�\�}�"�Ʌ�Ah;�,kV�򿪅Ë��D�yg�.-^x[N�����~�Gk�V5�yh� ���5�9�E����d��Ra�9wO6��>o{\�f���%Mb��.͈�~��(�ڥ��	\(g2�V�gM4�.D�D���`�amexl�qJ�����!���@ğ;���Ob�1=�c+9^^���.��
��W'�񴍎2Ɓ��PH�i�0��NQ`��H<�
��	��ew��<��}��KX� ��!��A;��*u�?��v���4���l�r&�U&wߠ�>'��9FZ����XP��A/�o�J@�F�$��0 �z�hE(�՞"u���zH�-���?�I;�G��)�+Ĩ�x��n��p��'$��g#%[>�>�����b� �0��t{��,ex]�P��wYc�l�~��:�,�4��KZ[�����Nw��].?	~�UDϩ��$-!-���JˡV����r@NY�ۖM���w0�`3�i%���]�H�?}�~��huД�}�S�'>��w�4p��Ƹ�i{_;��{Q��t@�z�y0<�!�,ߟ��7�\�N��̈́�p�a��m6.2��+eM|c�l�d�c��5�`L��i��39��幅#+��>�ɒؠ�81o+]x�7��׻������ta{�tI����[�C敆S�z�`9R=T�;���)��Z)�����W�(Q�'����@a�R�>���%�KKg}�;�mLQƘ<ȑ�"�vgz=�Ȝ�$�Ă�������@mU�a�7xi@������IY�2yW�A8k���J�uz���ZX��BO8�.�O�,�G!��� u�>Z�/�E�d��BncaK�.ț�E9�Z�j
��fo�h��./�%��w	"����9����5���f&���ł�=AҴÈΚ��)���%u{�4:�b�ٽ�"Qt�I�c> ����Cm����|����u��L�i���#?-Uz`F���'��V.Dʓ\Ys����P�BtmW�H��;K�嶊�T���hr��:������]}� ��~�Ǡ?����r)V4�N��}1���" �ٮ�z$9���[�)Z���7B�1���n���Xx&�W�٧�
�4��i) T3�U��-��nAj�-ZH�ZE�'s[����5qx����6��5t�
Џ�ո��p�l��l��j�H�d��޾��D�g�wɭw3�5Qsl���J�*i��J[�g�k��Ysc!y8"x4������( 2�Q{@�Irz���f�<Wᤅ�J��Aԃ �q��{��W(e��Ah���B��{E[aB��w�Y�/�R�/�߲�VZ�q�	�,��%S��p�-cB�����h�k�懕y��Xf!��i����qʫ�*C������ԴJ�)���-?Uq}o�2�jm3��F
�-���Md����'Qr���1NW�:4�|3n�=F6kG���&l�bNb>^��Z�
l���?UbPQ���O�^cF|��9�}6�gO�S-ts��x�hUp���x!���
d��H9@��p����`���l�.[產&��ĭXa�"f�cws�����^|����� <�-��C����KG�W�¬��I�.=�ږ��Ѣٛ?CF�N	������a`�0~�����C��@Kܳ���]	�5$K�2��W�l2./BEFD�&"1��F!(��>�g���|Q3���μ^���v������fA�8�Ӹ���2�8"��\%1*�?S�->4��+*�kD�zo�s@����� ��2xF'����?���~�-f�T]�����Kf}i��^<��:+w����E�cT�j�KSo�f���S�zD��n��B�.ԾM+��D�0ס�#V9Β�;�$S�"�9����^��� �{����T~���WW�JW�Sd�k�~:�Ȃ�Hs��¤�9]ʿ덄��]�����T�a��]�>�E/��{��3f{a���YS�M�W�Ir�|�ǌ��@9���<G��T���+�Z�p����]4��8�}�=rPm�ib	-�'+�3o�Sڌ ����|v]g�VB�[��%��tY��I�$?��JO��WR�P�GÿG�\Hd�q�rV����,,ԌϞz��[�Rb��v�HEJ~�����ф���#+����gX�C���T�X6yv���
�Z���L�F�R\��˶��e����ݳ���Z ����D��<�yف`O;�~�dc��MN장C�quyka�y��Ҝ�����NӃ@�� �j�{@�"�H��p_ ���U�Vo��Y{�&����%�y73=�0Rs���	�E">w�7cZ�Xshksc�'EZ�0@�W~�V:m�������EӞ�($�x��ZݭҢ�Ӵ�c�ڀ���V,�}h`���N ��{�}(8�
�Nk��O��"ʭfXU�K�f3���4��'B��,GJ�)p�𠲝$�F������J"���:��3=�����-�$�Ml�U
��4_�g㞓Z�kT���W�	Q����ok��*�e��>�o�o�R(�����`��B�?ӷ"SWr#��`4�u�q�?I6"�`��չ�zL��?�Y�u��m���[>�ed�O�k@MI��e8�s(��5g�6��ݠ��Z"��k���t@�&��J zB|뀃rܨ�w,,�(�c���ؼz��e�{�`-�p̋i8�`ұ�*�rÁ��<g�"t.��h���"gܯ�k��Q��`=�&zr֌Dn�*Z`�����A�f��\�v�5�� Ř7��B����J��{�3��������:�p<vR����p�]���:3�dӗ*�)X�J���@*��&�K�'�7�!۪6C���ˮ�;Fa���H˂��~&
@�����~!:�Ւ3#���i�ن�=`C��{���ױ��1��DD��E�4��L�hYL�7�p-KƆ@�J�bӄuHa�O���5x����[����GoX&�ܟ����L~�!�Ae!P���7;�$;dI���z)b�<s��N�-u�dlK	�L�z�Ü��0����Y8��2�$.�U9/qU�RX�$��?P�B�qV��p���OM��Ĳ ؉�O�Bgʺy���Io��E��^Xɦ�n@���,bl?s9}�n9 �5f[�y���ܱ1F\�� E����Qtx��fᵶ�s�W<�᝛仪�܆ej��2���`�&��J����]^����f�8�v�3p��bT ���`�^/m	����/�����2n�|���"Y����D\`A!w������#�v(e��Q&�P�ϔ]��e�6ӆCP�(�<W|�B���H7ҳ(Q�wYZC�Lw��I#�[˨!�yS���T��I{FyK��I�H��QTfV=Z��P�k8m��CJ:�\E�$�~��it��7Q�O�On	�I�3q��f^��C	��-F�)/��+5-'�� ˒8zp�&�Մ����U��,�Ԓ��\����K���q"��_,M �ud������+%��@��^P�i9{$q(8�C�"�L�E[P��߆єh0�N
ļ�Ě?����|�^7�0�Ȥ|t׾T�tA.�y�6�^hx+MpyƲ��
������9g�%;�C��Q
$G<�ܪ�,���(;d9��cZzYډ�}%�
%Ү���]@0�8��Y��׫k<�L�9Gk94���E����.�-[P<a�l#­\�cs�i�Ս�S��xx��A.�_a��5��[�ii��5;��7Z�ځ�J͌=���ʴ	wk����gW�P�x�PfB�p=��%t7t7����sZ�ǁ'�]Y��'�05��Wơ�.;M{�Zޕ�e��Y�q��E�i�
:�5�p��U�w�?O�����`�rd1�Ԛ�m�12�C������c�xO˨ޟ�`q:r�)�󥂩f��W�6T�Ly9���I���.��s��x�S/DS���m*�Ki�]WY�̀iI�t�n�`����:� �WfZ��?p�ԅ��lo�?n��l,���:�Gt�����|`T�Ko� � ��#���"2�^_��'���~H�