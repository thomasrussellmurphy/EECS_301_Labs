��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�i��a
Α1S%� �uj?�L�3��TLei-3^5]E�$��f�A��m��[ۮ�{��!b;�Q {��-�4<�a~�������)e�j|�6��*&�+9�䒽���V~�Ė'L�1ɞ�R뫇ϋ���}�+���w{�^Ml91���ߣ@dL��;!�Z�Z?�6�P��f#Mw߂��+%vSː Q�F��ѷ؃��`enH*+���(KL0aFgF_Ȟf�4Z�ƍ�Ͻ7�?#u^��w<Z�l�l4������p��v�"(o��r� c�jצ�Y��S�Q~��7�����d��Ҍ������hG��9�O�Ǉx�|
#���� 9�K}���0���<��@��pn�Bx�\�yO*�<�V��HUH�|vc��F�v�ʛWd��c�����n)��k��.�c�1z�I+#�Q3Z!��V�H�n��w���w�>Sp�;�7��@VI��Xr$��( ����ر�������&;ڢ[�΢��C�E��쉴c���NF�v���L�I���! z?��(	:��l^N<W��g�q�&Z.
���\H�������Q���z�i�d��ʬx�ǚ�מ9��x���.�����^�O��;L�w���%��Z����:t�$X�]��֞D�IuW(W���D/�)h��sF�O�:
��8W�bT`�᥿ɓ��v�/�K������E��i���9|/�o�{�=����!��	�Z;���aE}?�7����?6�ss-��&���I����?ɀ�U��&��ʑ<�(��2a��p�Eė�>`�8��_��o���wJ� �CG.	ځ]/�O�޷m�j�;_?0��_�pQ�m����\%���=h�1��2�`� ���6�"�U�*����}<��
k���zD[���6�E�7�'����v48����Ln��`�YG�3x��@��|�4/�\δ8�"�����U���8��?kR(h�ozxxq/;���C���#�{�����=�@���U�q��B�.����_��ݴ�=�n]�o0��Gn��%�z?��f.��;2�0l<j(��N��yl���QAEP8�:'��M�)�����+c9�r�g������t|��^�K�����E}���c���t�v�BJ9���v���-�X��f�'Ʀ:O#X�jt��7;8�iQ�f���>�?� L�'oЏl\A7��kiQ�����V�"�̭8�5Nc�#����%���b7,3��4W%�����<-urǆ�}�1�u�T˟�7�i�F!���Z�xl)��8dǯ%�m^�4�<of�n��Zs�o_*]��큀$ÞS4 gir��1e뮟�2,?��L�lt%V�
�H�W)�[��͡et��&�wڊ*���t7�C���>�G3@x8�{�A0�3�x�̶�5�1%��}�nu+'~�K�9�0V/��:�e �5p���M��Q���2�~����m��9zB�YL��3L&o��qTq=І���c�<&I��C���1���b\3"��A%��~�����q�	��6�%g�A��Ύ#)�����y��~�:>	I��K9�mT,#Tىm4u�����S�Ea��vu@K����H�k�ѱ�����lނ�g�w	y5����4-,��ˆ��dF:�����y��!��.�	kuo�f�� �`=�r\��d�'�\n8=�(���rQ�S��M@O���F�u�,�I������/���{�^�<(}`�T����mE����U�b�,����R�{�8F�(_Ҭ
��'��w�@��t{��T�Ϻ�[`%@�@������.鑊N_�K|���l Y��9�MqtDf�0\P���%e*�}-�34J�2Wf���V�<C+R4e��s�:�K��l�9�Kb�)u��*���3~C�wL��D��+^��D :�5�v)��������*H@�$�z��w��*b�Rk>�~z��O�,�"��K���{HG&�};�c��xb�~-����'੸���5������$*�p�/�{m�Z�Ln��h���P���S�_&A�{��/Wy����^��!�ݚ�p��$f�=�G���	�2Ep�t������<૽Y@��t�W?�h7h���d��4�p�A�|@�D�����n�Į�xtǡ���M_��1(�9�(Kf9Y��B����.�����-�ί~������.��Ů��'@Li�|)u���TH��h�L��B�VTf�_p��������j�4N��^�hG�'5^�{���.�):I��c4|P�k[�p��Y�y9ʊx��E�O���27��J&��`���6��#��ޠԄ������>��uҼ��:Lֈ-)�P�Թ/z܅�L�����G�"zN��Y=|��q����&�C���h��-�X���gΡ}H�H��&������̝��M/G��e������i8�����Cs�l�a�D�"9�ŭ�11���6�����? ���`�K�4���m+1d���^;�"�T�P˞/_K�Sw%�'S�mHT����l$��]��g�%^037]�4N��`h't�I"Y�Ot��F��X�zT]��vj5� �����%'	���U=�G����li
����{PC��%?+Sj��m%�� ���>���[Xb�g�ءK���m�y�O�ǨEN�#�������.U����ܲ1s��+D��ŧ�h1���O։��Ԁ����^|q�#[u��E��3��$u\�罔�Ew Gț�B���6M���Le��c���M��W��L�'������b�.��)�����5b��^�檸k"����� �h�bK��#��uw����ߖ�����M��4�-�"��]P�j%�,+<7� 8A����#nר�L�����/O�J���⹣��T�T��sو8�����4���*���5��s8p�$&r�%&HC����W����9\I�a�9��#\�s_��ȩO�@ز�]_I��Йm&�+�w���FjOȥ�W�J���jxH�N���ϚE-�];���U�D=Z��jO'q�W���'����:��Dd�ɳ�vtr�rp�թ;ꕯy�_��u�Yԁhr�I�
���i�������CD��MCY����~����X+"E�|LW ?a�m�+��J�(C������m���w�dyRԡR��	��wl)�bUPb���^3}��9	�L
����W��&�D�xΞ���Ӥ�̵�I#Su5,�"��{n�De��#V��2�$�6ȖEF����k���mN�O{��@ �L'�����4�ٻ�?6�a�6�dy���!4�_�Ʃ���j����~�Al� �ݒ˽�����z��+��֮�0 �,���m����~�0�2�++�Gs�����@]��4n
ȸ3o`�R���&{�pSzh92��nY�RW�yíV�`eZ��e���ߑ�-V��}��Q�������:Y�j���_���r�G�Cc�^F���#R<1̤dl�9BϻBB���u��l�9�9��M_�
³���?�k���-�6
��{�-\�	�u{ql�ۈ$A�s_�1NF�?�Jy��x̡�yř�I��(��)���A�'�x̰��Fe�z>U��X���s��wx�����#?��p�>�N�y""<����z8�a+n}�
��G
�>-�5W��UhD�VM9��?*2$�.�w������� p3��-7,h�oڟ�`!��	�哇�	���þ����dv�1�q��0M+�w����B�1�/��2�u��xOq�>±o�.1�R"#��I���{�jI��l�5�u���l���Q�m3�҄�����m���_�#GQ6�^��n�[v��h��&Ry�w�����<�@���]��kK���o�$�.�9,~���NB�0���T��<R�\K96R3�5�q�b�� ~0���-�?;����b��X����,�H��om �Ua�pȷ�{�Ϗ�2atr�P���8�۶��A�[���"�x`�k��P��ڥ�ռ�L�<� )j�"�7O�U��A�炧�n7���Uɚ�����lҊ���)J ^K���Y�t��@��#%Ao$S��?vt$������~/p�Q��z������{�Mz�9�� @t<nw?�.�0�1�����O�g>`�������PE��\�e&���8�^��c�8��I; �蓋.�w�un��G��H���|,�y�XY��|B�z�Ym��'�(ϗ�����`�Ĝ��a1P����Ŧ�B��>j�� �V�OP��x���w'{�Jt�����W��p�]�Ŝ���4+�x~4&����2��p_b�aƷ���D*#�a��u�a"�>ڱ���;�WS�$#U eg4�;�ጚ��G��N��ꈳ�[ɯ�	O��O!�DF4џ��X��΅8�昂�s���Ż���a�e�f��� ���[a���J ����*�m\���%\�ߝ�~L.W�&\t�� w��c�״�aa������ur�n��%U�U?�\�G��Y���ݨ��!��0����H�=��d�Z^u�jCl��^�*��RK�2��C�I_��$�Mۧw"L�)5R�-�����B_�o���a ���f��V��տ�L�nc��.6��5Z��.76�VT"�JJ���u�~J^�L����&1�*%�(�a�AR[�+��hh�f�n�mL��L�nbnV���_)t���Ք֮ʹ��	M���uj�{k{E$.r�q�u�<����*"�܀ealy���0Ye��Ex�t��כ��B~���"˙�'Jtt:��k^!����ס�c͸�K�u�N,Y�}�5�C��8�Q<�)ʎ9K%5NQ���W�B�	p�����"�x�\V|�,Ug]��Q�`
���v����K�T"����Y�'����T��,f«yJȻb)s�q�'�碌N����u����kH�������,P����|�U�Z]D�kM3���u�%|��	:Sl�L�-hdi<���1���tC��K�W�<w�<������(+I�Z|8�',��Z���� ��#�R��]00%�P�y!~���'�:���t��9���$fJ�L��+e�P�b�6MR�1P�h��)Ti�UOz���!I�"-�RJR^�$����|�+��[���)t���Z�r�s��ͭ�6u�X;p�i2��|~01 �t��YQ��R��������I�1`������f�q�^N~l���[g}i�1�fNZH��=T[w�OG���Kn�c�Gmqɀ���'�ף�7\�r���[���+l�Y��<zC�;]�|�n�v�Br��5��l�Ap�8�M�S]�5zl�h|+Y�&i%�� ���X$��$�3G>���9����@ؓ���=2��,�
f��F*q�ל\��Y�i�(��Sn�
Z�M_����0�r��!��^�n7K$�̣�1����l��x 0^�,��b�(��Z��1`$�͟����c96 ���
`��zScd�6�FEǫy2Pᑷ}	c�A��ӿ6;�+-	�"��fƒm+dɳU��b=^�"�*��~�^hC
zWp�I�Ռ�l�����Yk���H.~D�^��Cf�2@Rτ��� ��ǳ���?��_]�nG�ѷǶ`Z~�u�o?xӾb��y���	䱔����棨�,P�EN���'�uշ����#�F[�xЪ�;9w�#��Ix�q�r'����`�{?U���w��Gqꓪ^�V�iÏ�ֳ��N� ���;��l<����A_�?�gYe�F�\K5T����>�������#�2���1kz�y�/��4��iA��ܷ7�iCF��߂��,��o�P
�����b��2���,+<j����N�-��Zgw�ߢ�'�����J^'!(#N��w/�	2;(�.E�&�λ<X��ؽg.N1����VRo ������}�[��	ZZ��Q��q��^�9�*(���t��a��L���;�y�uBcC�V�r�E�~��P��I=��NI+@}f��&f�rt6 Q�����xE.�Ws~k5d�Dx�����˒��|3�kZ<Z"g��+j��3�r�J�m��Jp��=�vI+Q�	23t<޻�=��ղ&�J���(�b)F2<�;D�TQ' KnC+tS^��+�F+����X��\R�oP�Q�'=��U���W�`����!mv G��sI�����U��.�wXC��6���gՓ>I�eZ�S�^��Q�D��FL�q�|GN�T��	E�G֪jD�P��_��ש�ou���U?�z���Wr��7���9r*��Af63p��'P�W!��ӕ���R��R`�_T��F�s�"|�&g�
�lұ���m�}9�u(*F����J=Ժʴ�����t���U<�_]߉�Ҍ��������}�v"�����_i��33O�ׄ� �
]��
��������_�I�o���>V��M0�,[ޫ
�0�{�Фf䟅\������Vin)2w��M|����F�' 7�M���HAo��\߯��T��R�a�;vD-r���D�?�0wT�Wا��;�X��۲D"!����o�mX���լ9�_Dp�s�P�C'ST`BK�U���%"ȉ*�4i#��5#�k JX�����P��U��Z�3���s�&�-5���q�#Hž�����'0���/���G�a�]u�V�Ҏ�i�mA�X��coN���ճd^B����%�������ş�����6�x���G�����\ww<��O-�a���1D���Zl���ne�E]�Ï��w9~)��&�|:N�����#^
s��asҿ<.0��U��0?���H�2�h�p����?�>
����� o��Vzם��']a�7kg��u�&n`�����,�z|���,�A��-ޣ�y�C:��C�qt42�q��$H����{|��;���93�`K@G���
 ���V*E�IG₺̯)�E�y��c#G���0�wqV��#$M�aX]@��G�9O8&y�x>�^*��4���!��KQ��[��_����N�pI�����>&��h��>I�;��LDֱ��:S�?��+?��D�%ċ����������6j��&
d�5�#�d�"�3ߨZk�V����8T�dɻI/nY���B�O-�����y����3�vw�-]�ju�iC���V'[�~(��(��u�