��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\���V�fnvx��ÍG_;�ȅe�~�>���9�>��Y;�0G\�#���q�w��
A_� ������ɨXv{�҉AR��bh�bF�Q R,�	�� �� Q�#g!���2j�KnEo�a�9��>9���dZ�Q���ˬG�nh��d�\o.���� 9��X�T��Ϗ+�?���8͎�[��[0��v�0��֪���wG�$�JfcD�u�z;6�.��hE��)�\q}�$w��Me�m26a?]��H��#/#��p���ː�h�B��-;e�4wv	��]��R����'�}���/���ٓD�Q�"�7��k�_a��@��x���S�l��l}*�EA ���hno�����������R�[���q~�E���m��1�i��@�Y)�fr�h,�wdaR?ƙ�1:��' N#�g�++��N����.>�y
��K���Kz�_�V��_]�1x�vR�]�9���ƕ�f�^�$H��Ȫ�D�A!N��j�� ���)� �t�hk�ZC�}P"�>�h�)�P,��bO"�PP�9	B~]U�j�1D��]�p����F ~��M��ѷƘ�bB��n�.s��~�-N�h{���ɯ�9��r���KA��R���f� �&N����a�Ϸ��=���'�oN���6��2���GB�;���'"��p������N�w�g��8��=SH@"6�nʲ�1۔�&p�>k0��ɩ����J�'3�6Ny;m#�opkP���i+�4m�{��?�I5ޝ\�o�zw�|b�7�)���eA�_z���k D�&�[��<�I���d$�,��đ$��.�}����?���h�mJ���|5[l��,�fT!T�R����۷#�	=m/���[�{�M�!טs�q r�*'^�X���/�}s��A�V��a��^�o����n�lO�����rw+��N��XY�:���JsqC3�v��O�̋,GD�Ȧc�Ƴ'?�䭸�ބ�f�n���DEh),�
�-C��+a;�`�|  ��Z���� �!9v �����*�I�{��o��� �Va.�tIh�j�M�a�K�!E��}��(��S��y������mG��5�T�j)��.H��������$� 5��cW�N��,?�H	6�!��\���h��5�ꎌ=��}:��4|?D1�Rw����s����e���q�#iu����q���7������ry�3I�����%`���g�
�9�`6�F�hsUed�:�I�cR˘�
6�,�N��7�]�iQ�����	�F�c��'���b�������S2t�ŭˍ����/kw�.���AO��Q�����mc��B�����/bWn���Q�VØ}��"_�	��#xX�}t�����fxS�f�9���Ǹ��/�=AMo;�C���5�A�����R�ptv�<�0�ju�� !J�E!o����TE�6��"���_^L�(��:n
D%~�}�傘7|�m���Ն�E5�Kˋ�ihuK�Vk]����бC��1����|���bh�H�����+�H\q����ug0���V�ˀ���-�١��+�3�uJ~��~`�F�q��q�:�8��/�Cj㘛k�Q+�%��_!Ă�;��6�C3aپ�#�w� �������(��\����r�r�0�-��1�v�����A�ZTѠ6"x�/�r3G�h����b��e��M�R����잻��k�M�����D)u��S4��ފD���$
Lq�8��`�۠I�Ih4����3{Fp�6�@Р��u>�/�Ċ@��+~DEw�F���W(�W�4f�eH]��h[Cu�����4k�[X��K��dn������d��d��>į<�&d��5B|�'L�Lʹ��Q����veHD)Z]t�@�'�Z�e�����Wԭ���Ĝ��o^�]{��Ȥ�ܒ�\}��oŵ�(f]��02,+ߠ�`_T�M����1�ߪT�ˌgR��x�~�{i�3`��$���t���C�/�_.!�D{�a�\��&�hqiW���/��{+�w�.E��ű���l	�8C��ʫ���Z>1�����j�sWA�j�F���Y�MV02#����S}R pW��|�(q�j�; Qs���X��"�JJ��խj��	ǋ�Cҹ?�ⱸ@�����&��
UC)��J !�f�+�y�?ƍ"@��3Z�K�l6نs��I]K�+���V�&�b�0�@;��Mps�pX+7x(��:l����WlV���➿�>�
�O��Mߍ��~U�U�>V�L-Ƚ�,O�u;�@��L[�$v�u0�2#�&5Qe��|ƥ8V�)������| /�෠r]`��H�c�2����~�kδR3�mN�V9��F�w����g�Z_�����:)-���~iZ��ӌ��,]8�-��d������3� �g�ߕHH@哥�s<��m]o�(��X1�5�@����~^hѼ�q�7��\�d���=�K%��*K���c�q�",�F8nխ��	K�f٨q4x쎯��������)`�d�:���e�y�3S��'o�ޥc�@�G�_�:e�b8�a��﾿���[��8����5���=H>�i`���,���B}��OV�Z��{�(�9�A��%���F32C��܏.\x����k�!,�\5վ���#���fce��_�KT�n�1"�NӪ��]�A^G5g�F��B�� .V:3-�W�z\�����V3�������Nٌ,�y4�_{P�(�2�J	D�b��\z��2r&��L��:�]���G�c*:��i�|*S�:݇�w�՟҂�<dM�r�{�B@Ʊ@ /(�M��L88����[H�J�#bA�/ b
�����Uc��=���ܑ�r
C�Z�X6=��/߂�Q�{ʑ�zz�q��G�I���d�`�`�D~P3�S�V�\Q���X�*9��#�YG6��Giz�
K)^���@��{]-�g`zX�3����an�%�a@}����{	0}�{b����m��nU�����.9H�|_�������U��Ѝ�{��� ����:Nٯ���i�vJ��\gk_L�i�������8�6�3�~Sh�+�K����߇���Ê�%��-]�����e��Zt��Ri ����QC��h@ξ ���+��P�l�a�c>�'1�rQ��b��c5�hQ:���0o�@u����nl�?8$��N�\���,�鞫}x���3�q�釙R<�Eg!qW�2+ܓ׶/�\/M�ab�zg%�q�������%	�:�,���V��%�`Y}���`BL�X)|���� I�Y�wq�1��� ��8������\A�Ga!�P���&������&���#����-oS�i�&gU�&� ���x9�ˮz8�l�����p�ӷ�ΧE�Vb�#����%9(�����ګ�?̵�����&���$=�h*�C�[�&b<�&�b��g�K�4��X����MЇ�VŶ_�<x�����箨��^���x|�X��R�σ��j3پ�/�	�>���h���V�F��9O��sg'V��Ѫv��h�fĹ��8��D�r���D�<{F�0�&),��\۠P%�9ڷ6ꋽ�i���F봑���i
ޯX-p�S�\Ri�W́b���Hcbk*(�멳�Ucd@iۈ߂����aNe�o�9=�+���}.�o���3�o]PA�_�:��[g��&�J��i��×�:vLFT��X�b\Y�{�c�BR&������&r���Nrhm|e��,K�b�&�Uٝ��3�ޅz�F���"=�o \]�ꈦ�lp7x�����^y���C}	��ym*�K�`<gƻ��*�������,���f�A�K��p͹]e��ay-�$�")��䦻�����<0ms����u^c�ѳiQ�%���������(�v���J�p��}_�A�P�O��:&�Đ���;��Yv�5m���γ?/;�O��6�X�=��e�l�w���b��'�xdn�����`2T|%�w�r��fT�<U�ۯ<��T�$�]��M�
a�c�~��I��÷(M^�6O ��J��׳V�bB��.��z��08����bY	��8�;�-�:�(�y@�x��ꯇ1���n�T�'��Q��|MM[To� �V8lE�WVM��Ϗc����E��f�%��b��W|��8*"�Q��i萎锋���Ӑ+��	��'-�!�����ba��̎�H@�+�l�/�����T�N���ʈ|�1��"�I��ᓝ��i�K� ��!�5� ݌�t�"�c��>h"x�.ܙq��.5V�DV=^Md��A�&��ّc۵��i�W��!�p�)/��<�i��B^��:��{y��YlY#�����e`2C��t�@`�wK��m�R�_�3��Y�p���5�$&�A4�E,�թ���mP-�b���Ҳ�n�����cF@��,p���1�j=��ĜH�9��Lt�-8��Q�B�34-�
��QZK� �CE�N���E��:<��}���R�A_u�����n|ʋL�xLC�Oa&�n�ͯb�l�������O�X�-V�Q1�M{_Ʋ}`i,����p��}$��\J��4�8i'R�:mIA���W���z<����f!���㣷������U�������g,|�%�5X���j�z���^�do�E�KN=M�RW�WBe�a�A#��|������HM���@�6�:�0���>�g�H�dT�[�7�C.�"����;�αX�)[f��D�b{�����=L%!�3��p,�!�u�����=&��-!�+�T�׮uڛ&/�F�m�Gz���pAfvͶάq�-���xk�x�+�`w�z=�gE��Pð����^�"��e���]UȚ�.wO�*�0L�s��?���_w4�>@�T]��l��T�u���#x�T�dZZΏ��� xDҗ'NDQ�?��e��4�&@�c�����쟬�  *��b�)������{.m����\,gjd�9O��r����yF��L��巔�4����Fa-�H/f��+�i�ӟd(���n����@�(�����aƽ����R�~V�0���g���)>g����G�C���2w�.�y�.��W�ӬU��
�~��y;#,M��z�H;Ǵe�������Qw?z[��(A�uB5ޜ�ct�Мp�r��l� -ز�	n�����H�T�.�l``�%��=�E?�v�+�̡�H��q��~�j�4�EҎ&����X��AԠ=������fJ'Ƚ�(q�F���jD�%c�7-�.��c��C���@<ci���z��p?�d�i+ �oF4�چw w���1��+��E}�ل�&?W�g�8�HN0RCn�Xf��=���O�m���"�y ���w��U"M
�~�G�D�ĚL��Y7�1L뚄�:��7'ݝ˗�bW�L\��ɔ��Vl$��_/�Q� B>	�a5H|S�-��*����0x��\������<'���Q�^��BM/y�ݽ�e��dL!C��3��` `�3�p��q����� �q�\��LQf�Ʋ���� O��ͷ%� �AL		2�,��T�(�v����s��^��ac}��=�6��{\���;��8ސ���́b3�*�̉u�8_e:ĕ�|�{W�]����/��?{���'G��rTin}b-^���e �@/�c�@����Q��Ԝb���.ظ!��)J&�b����]��� ۉ����8m_��b?�<���7��֜BB���Nȸ>����q����.����iJK[�9^�D�WU���04.w�͑�ڗK?����7�����S�L�л�f�J�K�m�~ �@40u�>pӥ����o����?ś����H_�N>X=AS"#�����[��/G8[�ie�K��(<��n��ib���F9^�-�)�����6J��hTUEnB��Wƥ&����x��G��$0�+��E��#s�L��x?/�|U��o5���#�n����0��
Mݢ�����]ZQt���jc���\�8^�����B�ޓ V���� x��>?�$cK�m��x�wilN��Ʈi�ｈ���TK�V6����E1f@>���II|�b�6���h1�٧ion����F�~�OO8������FH5v%��[�B��C�oF�,��*��g�׮��q�gt!��Y����B�˻sRA�>a�6�PO���� ��6��G�s�x�m>Z��>8b)Zl$j����:�������Ϥ��7Q.Ǚ���uT	Q���ɑ.��/�r���|'N�XF|����/��9��)�}벡�ʮA"z�s�����0��Ǵ�s�� �L��l�L7j�$�!:KQ�0���P_�#TKϯ�v ۗZY����dXC���9ppx�0�i�9�˭����%�Ѹ>x��ʵ,[�+����˾l?������=9E�.^�2����MD��.`�_^ZMlh#AS���:L��Za�Z�3y$��3������ 
�X�x�.i��Wv���0�D	�%w)��a�������g�?�B�z�u�5Ġ�i�ce��TpY��/�B�ԗ��������B����i#��������\�2v�e�'���3����Ka�oQ*���k�Q�U&�ݺ'DZn�]4l�x,R��ۃ�e	#ʉ��^�~35fz>��l����	����é��w-X��7�w�]_f�s�x���:��L�z@�GV��W��Ԫ*_���^7sc@�O7��G��� =H�dUj�-��x����T|��H�bD[/�v�w�	�h�h�	G���Vnȱ���]�r">Ŝ�UO�5�ϣ߱�����
�����׃�m�wK1��hPZ��1D�E�π����8���ǧ�������g�<���e��'$��2V����b�Q�a��T|P�Sm����bG>�����`:�`���a�����dkګR�򆶍�V"���iDpG�@�96�턍�؏Bn�I�g5i�#!��+I��mN� �*Z���<4Kc)�Fa���s]cwV�������Ŕ�����C
?5�r��i�"(�'�mE�Z���)�-{@@x���e��}���"%���ȯ��w*����pKn�`��Z��$�<2�n�]��_�YH%��o2��b�ZYG1*�!k���=$F���waz&��'i��?�A_�]L��g{K�u}?"�~N�-�{���^=j/-�h�	�
9��%R=r/ĺ��'_���J�'���C��K\�#������`��Iׯ�3���~���k�g���"���k���3�(N��w����U!�K2@'��#���@�!����gY��%�Vu��5�l�/5Q�9H2 �*h� ���*;{�0�<Rb�-j�Ȣ��{�����p>���4��Tw���ͰR��3�YŹ�s���!z"�xm�$3q<[�{7>*p|O� ҆�r��Ut:C�G@4��,����
5��=�l���'`�.�5��7�A������'��%Α�n����� v�Jx���Whe��׉�0;��T�� x>/<�d>�j�>P���	��@!�lFթ�*�L�d�H�ٙc�\�ó�e��ڟ�;"����^a�w�P��>�HӠ:8�R�����|�ճT�����{E-ٶ��L ��������F!�a�O��\[*�x!������!���D�Xh'�
���k�+hk8 ��#���hq���L��F��)�s
��9$���&U�M6'�r?�\�u�<^��8EΆ�1|������-����v���)�),�����U?s:�TXaΣkg�ټ
��`@��iۯ4ad��Qjs��4�E��HL� 2 =�3�u\���#�i�r���U��j%ټe@H��ȱ-&�/��� ��J�K9wBeA���D���/ '�ec�5,�:+?�q;����o���cF�䨖)�I�\v�v�?e��ĕ�C[A���4�I&1u 1s���hB�g��/=~(ɵ:A�OO��$������Wf9S�r�N�(R�:s�ū1�;�����lu�Nf��a=�/�yCv{~"~�2y�8�d���֪a�����V��C���_�����aP�x�ԓ��w�P����r�_�&�+j/�̏�H�a�4
�jL�Ό�����0�q�;e�	��L�ZڷhE]S�����r�D_��k��̧��ǆ
�0ɚeD�#'����Z��R�`8-�f����'�����~�������%�1R�<{&�E7����Ҿ��H[��\=��l�d(r����Rn�B��s"t� ��!�w�ùMI�&e��9�~)[N4$'�e��!����7or�?o�@�����)�Â��C��`A�J	��kӖ�]���*�7�z~sSK��
������g�q&�����K�{��<RK�b`<�n���>�:x<����܇�jD3��
'!7��k���2�������r_o~���1"g}ǜ�r��[͂��
��#%�&� ޼��>jOd�����	vKsn��A�b� �z;������[�ic�\���譾�h�����g1;�7������ve���Rl��0������J�`—M�4��`���ӐeL�w�Σ�T��[vg��]+�iN���䶦�43?+´�,�F
s�kxp���r%���@ ��ޖFL��B|i���^�dh`r���B[U3�~�m!��\�:rsg$��22�Ɛ�kG���<�K�ʓ;� ���à6$�@�?j?X8vN�9����Z�ܗe�C�K/�l�}b�Hn���� j��l ��M�(p��z0j�d��8=
���t"t���:. @_ҵW`ֱ_��4��5�*�?$d9	�r��6i}�8������S���bb�}d�лK�.ٔ�ϥb��B��^n�a������#7q+SC�Ch��0l����ك��Ey������g?c�8*�9����#���^�j����6�G�{�7Gd�-�k�.͜9�� 0�9�S,MZ��GTl��������N��U,�5zO*��6��'�*+.W������)��+�J�YȨQ�b�wv���=P�}VùH�0�Ŭ�t��2-��!��J�\��/kze�\����6��F�V|�d)��j��t�Qx�e>.R�{6������8P��eX���[�{P`9ɕTK2����}j���n�4 �\�G9��%���Ö�|J���u�(��)��W�,^!+�����1��xn��
�]M���l�Sn�"zv���xƷ����[���ze�:������}Ft���{R���t|�(�Y�34�^9�j���

Y���om^�0GX�h��3�1S����GiO�:w��̈́��N�������u��)/[2���Ȁ}�o�
ď�搲 ���[+�;���2Y|�ȧIJj�2��̌����hٕ���=z��Ԇ�BL�a�x�O~�Λp~z ȟ���S����IcѲ�S7���D��ȣ�ˈ3�B(�
uC,i��3��ǘR�a����@9+X��[c�/)Y���ͨ��s���������ril-&���j����
h���t.�v9�p2Q�4}����bb� ��yI��'�_%Å^R��D��v�5�p.��kǠ��~�뿃ìO����v�YX�;6���-���M@�	mf�dmE| #���rFP�j��M�ή�#�� Bl+*#%PdI{@�Ǣ��V$bـ��@��$\��I�;�8V��`�/�2�ibL��ZuH�Rm$͵����i�=�����F*�5�����k�GxM�<5����@�
¯;JG����d�R�u��X^���paǏ>�%	ry�Է3�����|�EZZ�q�ę���%��#%YD���8���Q�0�)3я��뀤�C~�H^��Y�>�D��u|���RM���D�|Xn7��J���\(��Ч2VpjUp�F"���2䤍��/��׵#�%��p����=��D��ē��.^-"�z�NK�~�H�)���G�X�x{L���i
�"k���l�}�/�#����?�J�^R�Vk>�Nv��A:Nk(�c�W0��#L�כ�����l o���\ۄS�_{;��
Gؘ{��c�qa� ��oP�����0K�k��tܖ; r N<'ݣf�Tˡ-T���]m�S<�d �5� ��,���ӝ��<DIK��є�]}z֍��?RCf��ӹ;�I��ب}���Rk��|�sP��GX��F%k�B�c�q50�*HYȵN}'�n��n�������A���5�O����8\\��'A�	Ӈ��t�Gcͱ�G0�:���#YxMb_�����WX�u[���{[`q�N���}�Q������t�t��_���5W�(����>λ�D�X��*FSګ?���N�4/mv����H|�Xa΁K?x�M��>gر�8�����+I�r=*ꏷ��a�8���T�����@�`@�o!����ݧ'H�#R�݂.���:kR�G)��>W��ǩ7I�ѳr ��Y�btK�FU���D�et�����T�B�ӠX��6�0z)��x$3�_��J
���ٕ��(PJފ{���R��Gt���)Ew�l������ k´V�tV�)���5�Oz�Fl�)�r��0.��K�L��!ķ�"�\����8�R��4�a�~[�̆JO/�sz��=+����������,�K�p>���;Oo�>^��/��s�oB�^'�ro��k6��Ip�B��X��MC�[�TZ3��X�y �ukAnM�=��/�'����r	�����F��M��V"ۍBV�Y����.���F�c��6��D����!C���qj�XcH��Ͳ��F ��ǨF�8'm���������ҦjL����v_tS�_�-����ܭ�v�}�W��jբq�C��r���O����l�����f�?����Ƚ�K�?�ME 6�*op��|P���T/��-��;��BFUN=�t^�>G!����5ªL}jT�W!i��36U��>K�))�W���	��V�ΙT�pJh����u�jd?C!�n�;9Sg���֤hn�qD,'F�۶����K{A�VBP��RZ"�0MW�1&��#`����R���"~3�q �_ ]J�V��%S���ՠ�	�J����j�,		L��X�+ku�.z`��op$��@F0�k֕U�z����{0ڈ)���q��b��6�(�_�a7f�L�����6\�t۴�XֈUy3<*�)��-}�DM��Q}\�E�$����[��W�t��hW�7��X����� 0&�N��6>�-o�u��ߠ��_����'�#`�Y�Z����TJ��-�*m26�-2��p
�H�i^4�|�G����.k^4kM��/��o�)z�W��މ�h���P5�b�����V������	�ku�p+�/&Ř��~��=�X)��.ֵ��^U��Qa�MN������$�e V5�AV�U0�\9:�ԍz�j��,vaޝ%R"�)W�|v}�1���(>Ȅ�cyd�;��$D��sz��