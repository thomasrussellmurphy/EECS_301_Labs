��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��I�ɖ��)�d�~<�*j�J����yIO�=�;��7v��.n�O�@���;�A\��Sw44Bp�U`��Kb>:��u�������q��Ǽ�<���v!�E<����"2�~�N����l�AnqL���2����i����������s*����V(Ʋ��^F�/�/ӧq�+��2�0�Y׍���U�WR�˵io�="ٖ��Wj �	ж��:��o�b�/}> �c^�O�|$/�ģS��mv	H��Q�lY�?��.i��>���&5��H��*'t�����S^�@�ā�g�4����)�0X��?Q���z�a |f?l��ҋ��T���V��I�	�Q\�'�-�d�g2����%�%[z$'�v��Y)G��u��>��	;��Xky0s��ca��	'��%J0��&��#Z� f}W����h&���]
�m{���T��/����Iz�?�3��K�aƽX^�]!<A
0틦�]F���z�����A\�L�u�O	�K^������s���qI֞x^�(��n��K'���@���&&oL�����4{��^�ԃ��g�n�����c��j-���P��ꟶK��0Y���5M���-�=������);��+�x"�ц8�������,�t���ZT�	����4���M~%��~��X�T13�D �,��W����c���������ү�$A�tvo�d�u�4��ڠ���6w����*Wod�
�+�?2I�� [2JLGo�t��V��g��:%�`�����#A\���2��e�9�E0(�
��R)��,5H7�v�C�R�L�z3��"x�3r�:^|�]l�a^��F��PU�2s��fA���8�)��X����s>(���D�G��}��>�����X_d��������>��!ۙ$����i��tLS����}֜�����h�ϑ���!"qh��N�*��!=�WVTV`�bx�N��Zz"�9���e2&w^"\E��;S�`���S$X5젲[	y��Q阑�I {�=���� ���I����9Pb�N�VL���#X^�������h�)P{πX�剼X ���y�P�wS�n�����f����ؽc�}��tD��5u,@�vPd-�ɐf�@�}�%�=����'`���ԕ�_�N �����r�,��
�M�uE�S��jwFo���;u���[j$�~ ��N`;���Le�u`�7���P�"U<s��� �pW���b���A\ R�R|J�'!��6�nx�m���j��L���"�+�]_�_U�� �����C�
��Y�"?I�*k7��]���a1;�G�b3����\W����U�8��(Ok|���<9��e�����~�&� j��u8��)��K|QW�g�?-@[�ׂl]������a[�X�[����*⅗3~��t�i�n"��N��2=6}�wyTM8��6��SR���[:V�^�;��h[�6��Y�8`6�>S�F6� �(�2hVf4����,�G�V=�q�g|n�`��G�ߋ�[j���'�r�
�Ϭ��θ��\=Ÿ́4}P��yǡ��%���&."-���[},F�lT��ߴ��+}��|����?\����X�7)0�m�ƈ����|�2����2��4\^�=��Y�F�ɽ��ڠ���Tun�����edz���PFL�&�k���`�ӧ?d����NiB�tGk��"}EyX�0hm��$�4��N,{3E`�U�xp|��k���O,$mS�����\UӨHјQ�u���3��J^����e�v�����-Q�) �<�����eHgk^4�kN�ԃU��v^|Zt<��F�E���K-����8i��^�zŘ�ھO�LB�!D~� �GM��k�\#�e6�,>zO߾y�0L�'��QI����?{]Թ[�m��[��߀m���Obv�.��j�_�U�8��E%�Ӽv�Յ�w�te]���O�t�K)� WF�.t��)e�~���sI�	���ш~���ω6�#���_,�u b�]�߬�|�L"2~��1C��un��:�
Ї6%+��\��6��C���2��0���shG�!��A�Z2
8��x0�_"���l�������Og!�J��I��eV ���gp��<Q��k��	�-ﲻ�_��I�����-%H�9 �^EM%�7���V���(�U�61���޻��fV��֫g�ɝԋ<�]m�@㴩d)*`V�IZ���&������༳eo�����0I��N�;]C;N�iܴ����K�:G��2��Ha����ll�
+P)<"fT�L�<�
�"Q�՗:��:��O�y��}�&��s��3��l[��z^�n�㮑�e��QJLa[�yA|���N'�+���iY��2F��-��["�
)i!��x�0�>�)��+��ƛsc�P���[�	"꼼8��Q'�]M�t��:W����lN���T�C�:��� �l��f�dǚa�����+<���,��{����Gd����Z�bA�g,�I�K�F��P�\�����5z�	�e�ZS�{�[��.�`�����i��d�*#�{���I"��
q���K���H�@�"%�
y��`ϥ�6�=Mh�V���K� [YrŁIaB�:���7�x�,1�0�6+/ B�j�h
��X3�~����}K�a��J3
C5����$�޴�oRcG�3ޟw�e���R�'�n*byJ������'E9���G9�Q����e���ޞ	��f�'��;�X)C��M8(����f{�����Q�aK2��yGY(�v�dE�����7a���N8�uQ�VEB�Ds=�/}F���B����Y����n �����#��)�w���?�����!��,�c��p���Ķ�.�O�3|�?�=�2u���[ulp=9��a��қ1t.9�k�Y�c���S	F����NB5��E|<H��X�/��;�s�3�ģ�i�A���$o���{:���/��i�"R��ɒ^ќHikD �R��#��ra����_�6cPE2ce�B��Xf�b�M��;ORH��<�ʘX4�#�9<HLw�&'r�?����w���ݧQ=�j�8��AqG5�\`�{�bEE�p����r��˽�S)ER��|
��A���������83}����RٳBbÍ��cz�Db����F����d��1����Hd#>��b�-�t+��&����{`�X �gu�V��
�\�N�\�B����:#���)�����`��E�u����X�8u�3�����:��$l��վLHfg��l�L���A��hi$#?7�{��Xo"ޗX��U�&��T,���������p��j/�p�R�Y�rE��@��lg?W3q2��g�)���� ��Іm:�N�^v�j� "
��^�~je����2� fT�?���+"�zJy� �$
T�]�5[�^G����G��r��z(�E��*4��k��p�(;M���~��q_��9|�ΖpLE+e�k% K2��?����ZF�s#�T�:�KXw:�%�J$S_&�<��(�� �Q9k��&tⰯ,-Đ�cZJiE/al ���8�1k���F@��8y{[�J��u2����K�@H?�|�}
�I9�4��'�r�^�d,���cņ9��VRq_#|�:��������E��� z�l����N;��Oo ��B?88��U ��G�Ds�I	Lt{Xjrg��
�+x�FT�a�gn�E���3L�Jɛ�p���b�B�