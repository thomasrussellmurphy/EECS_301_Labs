��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\���V�fnvx��ÍG_;�ȅe�~�>���9�>��Y;�0G����2�%�q�PX���l&���d(m�A�h��[�7����J�O�
q��]�o��X�$�f�/njy�^�%����g-��b=K�QKׁ/�^��4h�7"+�c����E��q�d�0�;����ؐq��'1A�t��p����̕]FI9>�X�0s���hh�����4��{�8��I&k�M!���o�\ھ&7ڹ7�X��á�g�jX����O���05?���ҡ;�!��<7�"�����iQ��:�X-���n���D1���5-:������2��;�U1s�PL]���*v^����ـt2p�������S�ܶc���<�3�\�z�J�U!;��TڑHR`�(��m�.��#}��VU}��{��-ɳ�d�m��>�q���04';M=WD�/4����S_w�z�Wgn3 ���T����`)8��!�i�p���`�����h����`j���/��!?X�~�=O�~�b,������v�bm��������#�~{�B���O�x>�u��� ����J����FDF��>)�ZA�icJ:�h�8%͌}�Xf���ύ��4|�	+K�����l:�����R����F��*�������a\��ϕ�0������2�Z���J��yX�ԯ��5}{�?D"��h~�< ��V��]����iٲ�d�	���GQ��������6����n�B�ؾ��
���?�T��|>pz:@M��p�'f0��nwU��m@�h~�$zi}PR���dz�?o��<��j�����6P�EL�%���+pY�=��Y��j��v��R��̢G��e��#�]�q���
S��,�~n	�UZY$~�#��Li<$�mo{:�m&pC���X'�{Q�w�$
�� ���J����مSt����b�?��A���� ��}�6��P2��~�i�i\��]q���Җ�#����U�^_���EXW(n��R�v�@�B��WVk��^΍�U2%�ꪳ=��\�M�yw�4�k�q������ed菢�4`.�����̰f���W���^`���J7O�8�*cGK�_ �ק[v`��`��tOB�	��bސ⦷����_q��_+�����(v���v��P�}�y���*�0�@=�C��b�W`����]�KK�+뽱���±�ݲL�3�,���v�ArE�����=H�W�J��&�j��,HĻTrrƿ����ϫ� �i�*�|?S�D��̘i~���d��C_�;z�)��� �W��K��Y�RPi��!��a{� ,g��� �q��^���	� �Y�u��
�	w�-���#CEx��"֒�hX��@�dM�b���*6EW��,j]�~����#i�6�` }�nC����9�rΠ4C$RЄ6�\9��Q�h�(_�?�4I.�j/�;��@޿��`�~��rjI�7���7��BSa,1���.?��5�����y�Z���uE�&���}3<#�G4���ҫYΚ���!&���Yт�ӾO��f���nt��:i�����bT�1�u��Krw��֝v-�>�ߑ����f�
����d�V١�w�+m�N��cj�6��7x��ot2p�=IC��=�|��A�a7���:p	dt�Ũm��Ew�����ު�U9J�ȠU��=~㈞��^N'�v7̱g/��e���Yd��ͦ�l�Bh���H����TO�4�z[6���>��=��q}Yd��B�j��0��EU)Cx�;)_��:��n �=0���'��� ��}�]���(q*@'?�}Ȓm����/�y�[i�O�:bZ�r�(�H�Iz�#Z�L�,G)u<2����1̨VC��X˟�������g��%����7�[���xJ�*A �"�g����zI`5Oy��ё�³��ăXZ���k)،�#R3C�d�6���a��9�c����m\�^Q�hLʵZ��]�Ƴ&�h�	����A�d����&s#)
܎�ކ�
,�z�3��ڞ�"�	c�W2�S�Љ�3_A�u3v;TfNE'OSϣ��J��!�W��#��[��;�|��`9����C�$�{o4[��or̃�h4�-����q���gl;����H{j�PȿH���b7�S\���������h1+���X�#;�HH��T���:������C��CSv��[P>�{�6���i���g�I!oC����͂�@
�����t������N`#&+�a9��R	lF�A����"-�Tw���h��Օf�#Kn�&@C�i�֧&s�j�=����
`�fq<�2�bq:�ż�#A��mɝB@`U��X׌&�d�փ�
�Ί2�bYq���x/̠(ɗ�:�+�+�N���}�|���O^$HS��vk��ӑ�/�\(���0�>]�0�JCڵ����C>���+܈��b�7z����q�\(�V?d�$C���]d�,g8Q
��i��$>Ze��6��Ѷ��w�Zcwt�#	�A�P�!o*�5�:�#DP鬚�pd�OoN�R�1���j0c�q�Ň^��� ��B�\��8s�D�&s��`MD�*Y�$��b��ķ8􀧯s(N�R:�ft�����Gi�~
O�I��[F�,W�����csd+f�^Q�u�hA�"�K�V�칁եl[�Y�6��Ɖ�%��6I;�h9|O�B`�7�E`�F,������`)�E�������i 
;��~��6/�\cŪx�G�����wM��ɴ~ۮ���a��ծ�#���ig>��hZt�U�{�u�OR���W�P�C��F��=�����0���<�`�}I�I�K�����>F԰B���*��R�+�TMu1"�����%'�#i�%ה�TE�a����Z(���F��=�R�:�V܌m�+9쑮ktM��>I}����9f*$��D��.�_���I��1,DIع��X�[��'#��)G�CF��Z^>�����>� ����9�qœ���{���E����J"B����k[^�HFF�eX��B�@J�oc�|ڙX�g�Юv�c���Q�K0�O��N�b�b���6��3��-�ҳItϱ��u�O��`�M�ڲ>[��x�=��M1iQ�w
_��8�@����1k���v�'K�E������W�I��Ä���&�~��_Qx�u�ȭ���i@��wt�^e��}�}��;V�a�y�iw�
����0�I�}m9���wn2+ �1I��3�kR���E	�ǽ�0��;�PY\�H�ؼ'��5�K�����W&�k��0+�����>�>5[�sw�]؀�_����̡�R����K%��J*h��>lf"��V��]���I8�h�hc���R�!����J���~�`!4̝�m'"~?K1����퐄mL��n�
�\��
� M@K�B7��ū���R�(�g��15<�g��
�����C��P
|��p36rZ[�\m��YFw�
��-*��TɎ��f���*�	յ$�~�8���)-��4�7���{&0y"c�9Pf��|�AB!joN?�D�LT��a���p��i����=����	w�S��DF�@ ��6�+�)-�	�2��w��N�|M�t�5:i'kNru�m~Ӗ3z��	_)���kM�]�F-0V؉b�V���*%ir�RڃK�_r|��I$�G��݈⫽�K8Y
�rKq^�KcR���"l���s�!"�g�Fs𐜮�#����^�@���8x ����K�%$p�W���zlsu'�m��L�5/'|nca>�6,�XsB�~��M7�u�@d^%���<��{̝D�k����pxVR�$]�����<������wEX�qu�K�n D��bP`)��m^���I9�.3o.+�U
� �'s��Bu������ߦ�^ٖd�C�i�C��ɡ	[���'}��v��C�B�7������;�i�O)pK�rh���e���T��������g��_���|�k5%o���r��I�gf��#�岗ndw>�P2���-�I�j�l3y�������v�����˄	X�D���i�����x&��:�jt�[�4/0����_��[4�fY`����M�eB?T8x���[�#]ɻ�r���)��\�e-������VN�f�0Y����Z�j�vҕ�z���N��U�s@�Cu�����Ar���}�� �{E|@GA����i߄)��c�RK0�\I��<�摏�Ŝ�֯}�`��Q��'B&�oi���8��Zsp'�	�J�--+e��ah䡗i{�ZӚ֒H��ֿ�lyb�Y�.�jp�ੋ�e0���Ft�2S���R{S��ѹy��~?a��𺱵Sg�Ԗ�8|e�G�w
ψb�k���Zݕ;�ٞ��ʨ��K��f�� ^B��3)�(dX�,K���0n����5���Ά��<����
T��2���	��I!����7��9�� ����Ҍ�/-�A�S��������m�#b�B�.�"q�d3fg�j��~V�u�[V�$�młl�G���[`jm���#6Tƫ���F��� ��/�E�HsF�|y��.��$�p��d/,��.@���S�ݣ�E���2�ۃ��9�=
g�kZ�&U�#�j^6z�H8�~LB�����[��1��7�0��[d��8��Aڨi��AeV���;�S�ۓ37Z�8 ݄G��H���~K�J��_x
�l�������Mp�b#���yR�ܶ�<(��s�U��V����AxmE��g!�0/,ʜc����W�(hlV��9�z��Ig�l�ׅdD9��]������vy{�Lp�<����\�@m���'�#{w���`嗲�c����ӘjQ�"�jV�E��H�k]g�qRt41|1���ro��p�#�p�5�\}�����PyXA���P�O��Ȣ
��4��r��X|��#HW�mz�)�蠗l�e>��L�6d4v�:/���a*`z�v�6-xMWR�s%7�Ì�2d�}���%�5��i@�!u��2���Y
K'
?�G�����bm�ֻ������|ez���w���xt0N��j`g֙OmX%F��Y�S��h�W|;Uw��/B��j�Xr���#�W<���㲂�g���*�p�ts;�\��R��w�0��H��:������� �����n '��5�����V%w�~�r����@��(k2lx��$��.t�ӭ�٢���)�
��[҉����Pԑ�6zEJ��p�-jw�®����̝I M�%P��a�``��M�[+ewՎ������R�A��GS�Ă��X5�n�])=e��E���R��'�=�w��%�m���'a��!�).��6)�9_����x�<�Fk�/�4A*�aY˵<��� .��O˩�;��J��lݘ�7:�H,�H8� ���ϱ��Q���[Dk����_�{��@⫻��D�Éĉ~BN��m)��Ϯ�!���s��^�j�܂#˺
�44A����r�I�ve�Nz�>��$!�+N!�)iN�w(U,�����r,�ʯP�ۈ&k{E'��D�u��@�_u�L1W`s<s����ZW1��(�49��l�~��=�(�!����g�_᳦R�[��i1�8ʗ���+��m���k ��t�3�G@�	�����L��0�$�9�F�m�`+�����p�G�c��r�נ#��|,;��@Y��w$�
#���](��v�ڡwd3@)�".�l���p�;�Q� õ��q��I�Qw[>�a���y΢O�0�}'��d���	�qd�h}I���*X��Lf�=�['�K�V�my��N�r�T�`�w6|�v�V��z_�1�8��-�?���:P��\rñ���ox�Osn�*����YrE	7���t�з�Q�c0�[\5C������~��J��t�+,��W�/xI٤�=u�z}��Ne�8 �� Ξe�0Nz�_��: ���y\~3`d>�l����j#�]�XNb��r@6��_���ʑ6�+���\tr�N�z����V��x���TmF[�9Z�՘a[�rZf���di��&b��WЯ�	�2�˰���$�5$9;حY��D��:�Fl���y�����Ou�K�5>��D�x�6F&}�=��ѝҡ%�x���_1���������Zkw�PQﷴ&�"
�5��Ɨ�tT�>m�[q� N���n�# <~�$���G��@)�t�T��[r�&��z�DQ�ˏ����uF+{�K��鯦JA|�c�y�ϋ��O*��<��ǘ
�a }SDT<�5��푀Xљ�{����5���.�h�1߱��ڬ�%�0�T(��:��$y��t�9�S~lY�ׄ�]��𘄚���E �IݻE8��8����z�^�g��p�:�D���2%4Y�Ӎ&����?V��BU⨯�#������}�'"��ɣ�̏���t�_)�ت����{�bC�Ȇ���!�b| 2�p/��q!�p����Uȴ�0[w�+�|��0��8P�F bp�^����F� �Mʢ S��Ͷ��"�_U�,�_p�b]a��Q!�������=7�fSw� u:�\7�4O��r�Zm��8W�L��D��گ��D?#�n5�𚺈�i��ם{�L��%���+?6�F�u��y�j�͊'C'��]������U�^����ǌ�Qm4�q�p����Q2��q����i|b}��I��j���kAݖ�[�}g��Z7�(ER*�D�6g�_8c%ң�^Bm�4�š�Q ����_���u�о���z7��}���l�z}� j.�W2& $z������vtg���C�+�N�K��xm���o�
�Wwe%Yޅ�x* �/����;s�� uYѵ�,&�֟}�#�qq���@aX�m��)t��x�M��g�qH��ŕ���_�7�s�������aN�,��K�-KJ%ml	�)�@[PN�kii�N���n��{���F�C�K\�X#eIÝ?)6�qi�ϊQV���i��k2�WY�r���,c����(-!�[+9�7������KP��O�,}��x���#����Pb=��/f�����Ok��H6�RL�OA�(��ӽ��Q����5���Ā3<�5O���,�(�����I�3f�r=g1lr���2['�ZEMP�H��ޣ�s�)]#��˧�"M�y.�Nh���5�t=>v���U��C�*���f���H��sy�GR�#���C،�T�ґ^�yH���N����Պ5X�g��D���T_�C����z�h�'�ԑ\�='�H¸2�����<��j�Ɵr��-�sw�>#��P����q.�ؖ��qo+���Ps��ΘI>z�T�P(�����0��$zc#��E>�\����U���QY�O�JQ��rǻL�4�hc��	�"��5=��-��'���?wg�$�'�6�(
�x.+��}�k��b�ؼ�aL[]�������+�W��4�x��.3Q��N�u���q6=���R�������М�m�Kb=���wg׽���Em��r& �g6�G������@���B.EF�aG�?� �g[���c�1���[��X"��"T�4Nt(�1L����C�Ab�׮]|�����÷�i��
K�1��c��9�{Q��SOA�؈2�_��8�ƧR�}3^\�ܭ�e�4��SR��Ÿ�n+���^d.B�� ��#֬��l..���������XH��	�Q�56�x��~�h�����Gny��/����p� ��3po1'���[�`P��U`�԰�^�u�Ybtȝe� !z7�bJ��+P�����Z�-���v(9}�&ݖ��V�ٯeP	E���(>�����`M3`�:�8dS����D Ѣ� 2��Ǧ���*z�o��Z�k�H�H״V�~5��Q�#�贂U�F�(��Pl	6�V9��}�é<1w��]1�`��*nB�l����
xu�[Ffj6���+<H���=R%��!gӱ�\yV:Z4
Ώ��� 	KT�nt7�d�K��luw֏�/[#�]� ��\�5���蒜2][|��o�����} #x1'7�´���}:�:�.���V%B罵9rE�W0���
��rȠ�j�m<���^��s��#��_�]�*�{}b���OxHP7�n�i.�m6��2��"J�� )�T��ʝ=���@�¾�_�0���?���(P�A�_��b�X{�3�bC5k���� 9�F",{����1��Z��.8K����ީQ\3CIV��%��n<��{���PkL;9o���D���ob�	���ۈ�K]�vT�ThZ�a�/�Ng�Z0^&L��j�w�øʠtJ�ǒ������m�,�]JO���.��l�E�)���7\I��h؍�a���B'D�I~M�|�����> ��-������&�}{��k?Pk�z��<U'�,sA�e��~�`�cV��5?�!Ҝ��OR�� �� �1�q����"�Y��y�H�T��#���j����԰�?A���N�/`$�����[�[�:,W6�h&��=���騶v��Ҝ��zW9��,��%��8M@)���?���Hf��"�ؾ��:H:��"[��uJ�v�c%��XP�C>B��A!�3,��Vl�#�� �\x]���*�	����L�e1Waؓg�1	>b0@�?U_Ï�j��,$����Ti4�}�����H��T`�ȷm�MW[	��cI� ����p��-4�h]�]���Lg����i�wHGRN#���x@���xT��<ߥ6�QR���l��h�L�C������RE*<�'̌L�o� �|_>����t���%�2C�5���,�p�X�l&�A3<��st��
�E͚��|g�bg��	@����7���r9rS��/��q�Ͱ�?i�%���#�γ�����0+���%��׌}�%0v��4�Ω����R�@d���R�˄o��آ��q7<�j�m0{ � S҅ k��@�H6�v�
�� ���irQ�q��-T�[�4u&�cW�VҺ��D��ͨI_��Zmڷ�),ؓ���'�N��q����Lc�3�;x�^��k��K�S[^��Q�{ A�)ɸ+��Z;�j�9
�e�@��}➂�+$ECb����6Tb�p܂-5~� h�\"��f�d�,��ӳ���]�E���9W��`��T� �b�X�EtG��Ց����-vf�-��^E�y!�ٻ@�޽(AƱH!�-O���1��/�	�,cb±�Yh�sȁ�r>�8���������<7㫙Aǟ�!��igΰ��K��/�lrϕ\c/��ӥ��X�i�\�^�!��j-ˆSG铊#?o*�Q����ׂ����q}C��^�)$U4wY2�`�/��`���/Xѽ-��\Nmb�J�~>�U�8w5���HvK�2C��D�p��i����Vɾ�c�����d�E;�Y��l�
Ut�8�ڪ��3${��v�
�YumtU��������Ɍ��ݔ��^�D�P���� x[���:L�a�g�N����wj���Ma�-�%�������^h��B0��pg.o�a �B�䠿�]jM�7��u=N�ګ"W����)
�M	X�wbjU�����W�/K��b�~��S�G�(b$����Ξ,���C�欆��S�G�ɕ�6!�v)5�GJ��ԁ��:*y���E)�ݹw_Q�����st��$l�ۆ�(���?T�q+c?�|
��K�3�zH&K��VE�A�����S��DAѽrD�-v5{�XVa��ȱ����w�4M�s&�C�晞 ��p�"�:.3+2�Ϭ�������	�q�c��V̡�gkaG��bD���w�'
k~н��^F����l�+�]c�<�7=��W��KM4��I5��/6��O���`��_��X��CT_��������[՝mRFX���jज़uUD6D^�S����.�%�����z|�7ޏ�"rjKM�4U��~hw%c���[���LÒ"KK��k��*Wd��1#hW�NM��CD�/�+����q{��%s�^��{etqA��s�H��~#:�A��ޅr���yc�_�_��j���J�����{��s���k�?�8��S�*��{:h�/��P��\G%p�SLr�gYY��o�/�@>1���ϰo���o�h(q[����+����a;9�W!�RS3�Ke,���������b���PIն�r Y��R� ��몡x�H����� �������z~+Sj2�N~Ɩ!�������=R_t_mU�	�9j{qi�S!�곭U��d�b8�x������&liXC��(��A�yT��3+�C����j:��MFY�`(���2K���yZ0�"t޵����_�uq�*Ikx�s?H4���&�*6�J~�5��3[�m�Y,�z�Z $�'�~w����g�y