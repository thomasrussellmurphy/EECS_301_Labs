��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|�L��58b�Y��u��]�R#��2�)�F"���s卺l�:m6ӕf~��AN���$�I��+\KO\��|�*ƮA�R-�?q��)!ڈ�l>��?q�8On(|r���?�T(Ȧ| �l�؃�т�
����]j�
��EB���ڭpQ\�<�����TS����T��Pf7z���v� }�Th���7r�+n����C����SI�k~:��7����ڃx�y���W�k>�tNd/`A����o���%��ux���sVxe`�R���Y�9k�xB�@�w�ti9^��Rvg}��R�i�}�{��VC�V�/��0�^i��	{�M)/��`��z/y�q�K�k� 4ٮ�0�SYM���� qa�Grp��R�y���Ю)@�b�֘���c�R��Kk��}<;�']�#	��ϥĂI��i9���H ��@S�KU��^C#x�1��C�����$ϰW��22����N!�'�?���c�}FM�(v����t�}N��W���H)xP˷X�B�|WU͒hH�*Y3.l�/���ȹ�{7�"��IȦ�k�H�U.ji?=�J���4�.sM��"�����G��`*�����S��:v	W9�!.�C�GNS<T���3���;�>B��o���#��hI�ؘ5��{�D��]��Na!�5�s��/PR�I�/�� �^�@G�;-Я��bh�l��0�:�oDl�k�7.�Zo��������k�:Ɣ��:Z��a��"b�0��:-����)�6��Y��Cb�W���j�B֠�)��~p9��K��|ĩ�[�'�&N���g<ZG��qi��	���y�'l��tM���&��ߍ�4��� �hx��e��X�Hf�6V ��C�z>��ߪ*���k�į�
1�������q�z�ƕ�4��\"��4��E�����2"�7���f2�fu7��f���D&qu<���It�� ��z<T��ew!�G@�5�b�Gߵ��^���)3׎�̪3��\�2��bD"�.u�՟�f"�!w���t���Q��E]N����t�%l��k'`_]i���ؠ�#�|9��QD����r��׃����:I�c=T�M=W����~w4k��i�J�imuѭ;~\(!#~��F����&�ǿ�?�q�f�b�����D�[|\-9�����q,:���0A���D�p�Ξ��Ԩ��=:��=b	2T0�"��3{��$�� |�&���|��(�a>��:�٧�����S5�
���b�Rk��m�,�1�P%Z��HT��#�<K8�&���r���"�A�?L+&�~���!T��iq�\L�I�E�K�*����l�,GniK?7��'R�F�� >��o����Z���/���흜�SN���-��Ě^ƯY2�3�S�g����x�8�-Scuh��Z�5���#x�?q��b.e��M�+F����p�<�(���:4E��f�����N�Ym0	R�۲���RF�ω�ۑ$�`u�$d`��K�C`�pח�y���]hc����%����]�s�(���;sې���όjT��?�^A&���l�t��ω\XAJ�͎܂
��OВ�����d��'�U5�8Zo����^AfK�#y������A;�6/�9�t?��qdC�*�
b1P�&�خ5G�)'���$�M���E����O��r+�8�f�"��Ҡ�^�M�~{���4��!��+�/�������OU�yZG��պ�H�rI����XG��tr�x���tⳢ8$�����7�i�)[�V�~�s�7�
�g���g�=��;_q|�ƞI�%,8���>�w*��ja��q8�T
��e��Ӓ���I�e�E9��-�	p�&��jͰs^]��)�Q#�;�3�Wο�4�V���;�`�T�O���X��#�`�8�:� 8F�]����,�����GB#z���+ڞF�V�i��z���գdk]���A��R2��c�f����zD�,�DSE��z(����-��vK�j*\�^J�uk�]Ym�,S��؜�^J,���A��R���U�aP=�YG�i �e���i�q��,�Ayo=S��֒�*�����{�=�"%KS��3]	���!�-���yv����.+�TꡫD=���Ѯn�j<A��
G�_���rׅ�_<��̿�����*�����dH�~U��%{ah����n.���S��$�M���a��x���]fz�������0�dO�es���c�sAv��n�>�a�`E+ԅl*��|���q�fU��	 Kπ���N�&�w6C����3>�{j]w��7!�MA9�8f��}�8�؄_��umu�e�ǁ��l݀�}\�U���C��h������ EQX>پ*D�+Z^.�TN�b���Ķ4�2~�i�44�ƆoӰ�?�U���[S�a�^���=e��a?�.�Rڕ̾2�'�UC�&c�ï�񨥩�
1��#�$�
�zg~Iz�{&��@��(L��.5=^���Y�ڂ�%ε��Q���@�s��g��d+v�=�f*
nc=*o�D  �;օ埞a�0n��hIV Kg���8;[o]L��'r7��?~	�����/<�b��_Ș�N��{�~)��!pl����A�"wf�]���V@�ߋ��a�{P3�h&��X
��G�"�[kW��cͦ�Mс�f�.E�	AHę�s��r�gFO����!�~z�M�ٚ��
܁)��P�(���Ԗ�H.L�
HQ�Խ�#�=��taj�V����Yv֮��B�r�eF�������8��@�/$�R`}�����F���9���RJrO#�dɐn��H5!��R%R��y"�O6�����6��/r���&�dcJ��2-- x��"����}���-�ґJ�Z�X6��}�tZ*�3^!��*�T�Pv��F/4����r��2��D���?�)ʜ"1�l�~�C�xݭ�����r�_�;h5�����w�h�C�EV맥Y¯�Gt�X:#p�A�m���!ԟ�\����<����6ͷ'H��~�('eq}!>�,�}p�r�t��,ΙH�/o]�[��!��Ω.�U���wbV�	�ئ�{�&@�?rW���H���(��.��;��W7@�4s[E��\�����7Tmx�����)����N�"��6	pı-�Ҿݢӈ�1L_7M: �#;z�<�r�@ÞW6!��r����4@�C�����s�}���	����x�Vԃ0�D\Wdީ�|��Ë=�/����m���:��LMJ�$¦5)�Y��$A��:���>�����r��(�~7̘/6s�Y�����e�R�.�>U5�0���ϭڨ������χ��[�i�i�ï