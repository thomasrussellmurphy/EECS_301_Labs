��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\���V�fnvx��ÍG_;�ȅe�~�>���9�>��Y;�0G.䭈N:�FyZ÷}��K��c��,j�/��Sff�_?JF ю��Q����\ѥAOqb� �\l5҆8`v���˼��V
	{��NXRB����u3<c<o1/�D��!��~�Lky�q��G!�%��/�)�u�^�9���$z�,ۿ8!�*���߼>z黺3�m	zms�M�%������a�L]n3�Ѷ�#uz�Fa#ރS���<pnh�o�soٚ��'/y	���#bw�W�}盪U	B[�1^ʹ��sAlJn)i���֌~���Grw�SYh+�+�nXɤ_�������liǞ��tfG8���u��9�Z?�D��]�)U�P�cI$H���$�ȱ<t'}��2$a�?�5�ޮ��6A�����l�S>�I{ZE|�&G��8x|������s�
�'���q��^�<��p\��K,����t6�I���:X�t���o1�ȰQL�f0�2�
r���+5��M��Jf��ʃ��t�)[��m����a댆��m	���ǩ�� �R���<S�C���-����4B���oR����![�
�!�"ĉE���Oj�M;�~l-�Y� �P����xsDjް�B}pT�B�Ö*��!	cm*�Ew�$f�������9�}W������b#��Y	Y��a/V&���d��;W�l��J�7��G"�=r��4_ȃ��y>�������K�$��+*�5���La��
�FH���������&�� ;ʮ3�C���_��h���!�Q�b6Ps��i�6�a��Ưh-I���`��������`�*.��A���*����u1.F낌v)�����̑��m������V��J-Cc����ݣ{dI�%�Y��9_Oar�K���.�h���h� "��0��ꢌDWݽw�`W�ے��[b�rL}x�~"柞V�UF?�1�zw�k?��豗���R�h�2Zq,��!}J�q�Z����e�3��a�#jR(w5�tm��N $���{2u��T�;�Y�?���E��BZ�ʝ/v��ӗ5:	*k
��$8R8˙*]!�F��iY��9\_%P ���!��?0u�Ř�|�3�d�6E�_ĥ��6��j������}3ƮA7q��2\��K
*���ʟ��Km�����(�S��m�1L zs>�]�fa1O����ZF�,SU����������{�,��8s[�롇`Q����!�g#�N�і�h��7�1]�"!3��*��s��y��yH|�����6_�C8�xx��=_�e�RH$5�J����f6{�.lT֗�u+Դ���ș�-# ��vQ��RM��Cb�,�34�LP�xj�dcyH���/�>I����n�&�o=�ᬽ
&x��ۊ]������N��\;�f���oU7�I�}�J|��X� )�VO2��9�Y�-r)�!mma��iT����|�~��q��}��/ ������Tؿ}�K(o	�C���!�͢_������ۖߞ��hi}���0��ʌٿN�k&L!�M��?oM٘2|B?vR9��� �悩ԑR��b/zj��*�t��n����Sᴖ(���1݃5�?e���[�����rÝ�Se_j�O��.7V��k���O�&"��l��z-H�8Y���4
����w%g'.�;nd�̏�[�v�t�:c$<��Wa0�/�>u/6�RJ�S�M1I���q����pɦN��c���4]����6:�[��D�˿��4�ѕ%P@_��0H
a[J�CE�K��E������I�鎼 �B�}�+�Y��w���`�`R��"�a�+�8����
�Fi�"7D�������i�{��b��[�BZ�M�,]H��i�@��j�s78�݀Ux��4մ���Ҵ-K�K����3��BC���~���i�4���xo�k��v��ӡ�����}���^����ǥ}��y;��y�>���T��jE�Nr%{�y��T\��LT�$�#A�5 ��)��G�~��Y�@iQ�b�ų0t�&O��"'�A�J����`V�n��wf(�/�m���5�Z���2�0��iNh�_���t��y˰�o+�&�#�""5�Ky�Mg����
������(���P��H��M�b�E��gܙoSø+I�����Q��g��p��E��Ev(����pJ��?{-F�!�H�⋙�����?g8.oߊ���e���t���Z������\K�?���"�QM���P�����Q�w��@}�ǵ��M����u��F$����T��~Zs ���K�	�Hc�{�D��jߥ�(�]��҇Q	�`�+��E����|��N�F�]�O$!��l�5"]C�q-BIE�5W�y��T�d�m�7[�P�:��*r���0��\����J���_�1ܷ��R�[�����#EU+"��:#)���Â J�=���D��3އԏ��t����E��aU1Wip����^�ׂ��4'���:�NH�Qbj���:�a	7��쨝�?�&{Vf��]�0_P�tOg��<v������H-��뚼cD�F��Gw�"9��Ը����s�\�-�ͨ+�X�C1}��g��ۇ��TV�;t��d�Ll)�ɽB㉆ㅣ :�O��{)s�3%�.�W
��~�\*��X.^���N����I~�����u�1�4&�̒��-���̩eP}�QxR�hd/49��=�A���sL��8Ӌ9�� fJ:�R�o���I���
��B���#�#	d��$%l������炔�q&����ơ�;� �Ʋ���WH������K}��\�=�㜵1��Į�:d7�#t��[�.��4�U�m�I��T��
ĩb�t�� t�*^T2g޿�v��۞�� ��l��f��Ҧ���4���JƓvm�+�aeT��Xhm֭>�ޓ������Y�Z���C�Y��Kf>%��~�.��r�xk+��~I�V���4Gq9V�< tFֿ|�9�Qf!��+)j����97�Y���#�h(Aִ��]ٵ 'y6#�v�7�f�`���gA��k&=���G�x�����R����dZ�z5^�,��c0�������pP򼫬Jh����> ��g����sW�X1�>��lq�Y�(�`��I�'�E��7���Iq�Я��d�Zq+zi#!�nQV�唠dK�ٕ��l��{�('�$O���l�r�-��Z�(�<�����?6�aϱ��BY��Q�T'qy0xr�`W�����O?*.��� �ܴ/f��}��q��E��m+�"�s�t��J�)/���}�;l��D/������J��@�`4�;ԓ���>|�B�^��%,My�g5��ۥ�����C�j�"駃5�����v��w���2_{.�T<p�^!��� (��Ay�tշ��b=L�z8��×Y焾��aC��'eX����rǫ#��J4���[8��R.6���Țz�艊������Pd^3&�@�)!3�%���̐Y�8��RG#͚��)�$�=6��Ľ�!/���<��X����S Z�Rv����ҝ�ա��O�h�e�ܜ��+�#�����B;���?�X{w�c]\S�5QÓ�ޗf�������9�c����\�~�`� .�J)ۇ���@�UX��̭޴\�&޹y��eg}�	&O �78-'#v}A�^_��Wa�V*	��%3�\l@�.�zD����]#D��!z����[ƈ͐�h�����6��
⻟}�Hr�ߍ�U��O���L]�`%�TI<4N�Cx�f^��#�&�/���o������ �{�'�Bv`{#�[�H�>O��/����E��*��(A�6�'�D�ʨ}Xh:��.�qKs[���K�`��������Rb�p����wVs���R�I�k��`7��I�G��G���`����M����=D���oUрp�1��D���7���O��B�E�Q�ɑ6E��n!�!F1��f�IVX�:籷$�7�e.��A�w�7�b#���m񝖢X��T3�d�Z���b�����}��Cl�\�̈n���oG z��Q�*�������멦�(�P��,3x��SY;�T�ɻ� �t�?��F4w�A�]�Ѧ��1�� �}����T�?�2�U��ܺ���]���jm/jh֯Lx@Rw�1��i��	�@�-��$�Vq� �݄Fd��g�:V��I1v��Ƭ�?"N������2���M�v�[�iN��!��w^�;S��j�h"̇>l�͊Q���������2A��{�p��?{kđM��D)���Z����.Vu��1�IBV?Mx�XCDʆX#�t�b�]/5oh���}%6��vh����^W�˸R�
�=w���eZ:�K:-�kW���`�DS����������N��Q{����q�Ia?N	�ź��``He����	��-� ����錋�����hS�[�����	��;F����(Ʃ��D�#���Qa��x��EZ�c[A�!EƿY�Q�
�7Oj������i#!�P��A��9/��U�Ggk��(ń���v�����G�$5��tZ�4��$$r��*>�0�@��~)�y{t+��W`"���uP��Т�Q�- ��@����=:r��z�`}jː�O���%?%^/iΊ�#�$(���ȧ���Ԧ�4�aç_���Q���!�r�[r1j�;�
��!�0G�m!:����Χs�,�R�ìؗ��z83�����1!��i��^�|���+~��-I�(���Q�E,2G�,��S;���O2�����?�!���B��,� ۃ1.�*�!ip�X�5h�оC��<��9�1���@�B�+�b@s_���%mv�2/ȿs�f\7�I�10��aUTc�}Uc�U=����3MO�O�Ws|F񏼕R��*��V�r<��.~?�����#��NM�^��ݗ�ɴ��Q��7��t���u�uQ?���k�?/\�Ke��Bk�6�K��2��y�~}G�����Ҡ�bS#��>��/,�!�5��5L$�j����d$8�O��J�͋h^5l��1%8��A6D�8/�:d��i@E�_� g(M�|E[��Y�?SlG����%pb���)o�{��t�^%�М���<���p�uIHx{T�#���ȑ�yU�c��:����m�ps��ɝXﵶj�ޣ���߼�=\)�&��~\�Q�{B`Do,
G�� +I(�� "/�D�Pu@g��m�X��}_}}´�J$�?�nO�5��\F"�u5[����u�0N�0��0�4x�2�옆e� &�ًU�q�}'c7\�a�rgN0�3�������q`����oe�8�P�Jx�FE]rK���'��3��d�2#���v��M����X[��
5�;������b޺I��ƃ�ܔ<��l�[��@�FA�	?���9�n�xo�@ׁ�WY ����ŝ���z0��Nr(�b�#��P��$�t�]�1(9�l#W��݆�5�Wp܅��z� "�*���˝�/kQ3���+p��g�	�S�S��A�9vA�(�S ���6}T�Ƶh�ߌ�2!�Ǐ����/�:�x�y���d�.v�;)PXSw���N[;J�tD'Z�/�� �=�`'�p������	��8�t%�4�]��*��z�I/ʁ xd��C�6T�E)��t��et����u��^j/X{#��
%�d�j��������=��<5*[���o�/ćG�jY��
�my7���^V�K����L՘��i�o�����_M9J��:��u$}�Ӷ�6Sۦ�|�?�Зf��k��aZ�f�}�S�����jYA��@#)ͩ�B��./>�����j���zp&g� x!�Y��	
(*5ޡJ����sjIS�P�|h�@�rKN�ŶI*�W��RL��FvD��:�\�9*���V'
i�=���:j9C�$d\_���+�TW���.�6C�A2���i�n�w�K��A���y�| �b�8r�ѱ�|T78�c����M�~^Cd:V���kr��K�>F&2�&k	��~F��y��9%lS���\�������paX����Q�xf��HH&���U�Yk r�����*�6k��������$gT/�+��n^KwY��}'R���"s���!��xB��ّ39<�d�l���F�(1�vVK�z �l�8~�E`��`������n}��&�n���s���ݝ&�'���iiz�v�0�Ǫ�i�*z�iZ��&�Ԟ�0�>��e��D���_��/���b�����ӧ��G�$�qc�����6R�F�f�>�y�t]7i5��.?��=1� 5��> �ղ��Q�]S)WZ�}�n@��A{_�(g�^Ue��$�A�.s3��������ۮaĺ�ˮ�Fn�F�7k�b��5B�5]>�� �!/MV��hu�iJ�^�g8ۚe�b��S��R6H�=̎ʟC�k�S�_�$�F�+nr���-C=m���m�Xj���po���P���}	r�����s�	���ٔF�	�9���͘�}�I��	E ����	�pY>UC1�bijf�����/� Z�\@�SJ�.st?�������sE�� "������;��ѯ����&h�}.A���<�����S\=���o�&�XI1av�A#����o�����t�j-��K@p>yv<�eD>���pa	 �̸XB�.?����\�vW^��v��f�g)k���:`2�����r���!<�ϫ��� �5�唰6t5O������1X�[��q�-g�:ڥ=�+��@�g�)j�k����&��p���m�{M?/*1��l�%�
B��`o�E��昷3���(B���&=���g �YK0@���6�-���VV!���w�W�*ZH0zE����[N��~�$�J�p�f����)�J��fm
�������9�v��_����ޥ��*�7�0���,��.NI�h0P��fBڳ���38W��J�Y$�@!%�?3�<�B�� �v��v��`��w��/e���8��bl�5���z��/q-(a��"�2R�zlƋB]6�Fj��,��p�@�����jBB&�.���J�~E�)t�[����%����yq@��"�]x���
���8V���z�7�\��(�sVڕ�ku����(��>I=��#h^uf�*�m&�Y#�|U!&�|%,FCt�T�k��߿k�^��l �ߣ�h��E�.O�D۞��0*d�>C�D>~�D�D�����ɑ��~��qM:��%0�A�9�K⊻�d�83'60��q��?�<����qK�A��n�����0�;j�Ւ�V����y�S�X��Ԥ�IF#�3v:���xȝ!v2��T�7PC+�C�(S'�����-3J�KeN�'ZK�|�eJ���������|Fj�{K6�e6�4��$�r ���V��!��d�8��iakо�#1@,/��Pa9��K��o���d\^��������p�t5�gqZ�:g���#c�Ϫ,ݍ�:s8�Y�nյ�N���tJ������������n��-�#��]�$Oŷ�c;(�7��g���K�?��m3N��g��5;
(��8-rY���.Y����v��>�]sO�	�F�K��@�L���	s	�Q��k$篭�gbhy ~s �0�Z��v�I_ذ�[z ��*8�v+��Mq����R?Jj�|�d����
�����$�x����0��b��-o.h���1]ٿ�A���I�	 �} ��m �6F~̃�)jo����̱�W�oe��G%E�Y�wg�N^�b;�$��e�	�T�|	�Y��t�:���e���'������+|HK%!t��n2W�������a�۾�r%m�}u4U�9%�Y�ۀy��P��[��n8}�~M)B���Ϻ�6��Sq�<�uv�F0��	Ab2�?�M<X�a��3�L�mg,�/���n/g�(I�Ɏ�^�;D��7g�������3��^8"�Ih�7U���}���X����&�D�5�{��`�+�Aٶ���\� ��TJ��ƌaU�gLQ�5�F2���Y[��RN�UY;�wV�_�Vimp�.b��$�B�C{�"�0E�A�D�yb�|��d!	��m;�Px1�Ͱ �f��v��bi�(Fg+g5*	F����U��O?�37�і܋]�9��qzX�È�姑�X��1�7���H�z/d55�b�.t�M�����˼O�Q�o�Zʚ��&���5�q�ù�,�� i���e^���6��Y�N��l��� \]F�t����S�:��b��̎��~�%T�ur�+u̸��Cw���BŨ:I@~�N{@0�z�"�?%��i���j��]5!n��GGo��,l���d�$tMJ��O++̥n��d�0�Ȭؤwb]7������������ϛ��z��	�\�(���z�w�����rWo����Aw-{�����"��`���`q�>��'����4�.�ўx����bOq�H��r������2q�v�� �!z
9�����w���=v%�	YE�^RG��I`���񵋺�~	s�j���Q�1>�?�p����S���	�{1�KMd��8�Wh���5S��%��� s_���kg&��^������q�<��L�"����Ѻ�`��aC� �^��2�Ґ|:�&��?�b��|��1�a��<� ƌ9x��xDP(��JE6��F�����Qh�0.	���g�!�8�YOY��s�>�X��:�����[��, dj���s-�D�x� Ȝ��ڐg;ju���tI�z�G������b
���Q7YȈl�p�4�-P+���ށ~xwz�	��>�'6`�����:��a�*W{G��H�)�[��W�Ym^���!�cۿ�2�;U݇ט/�OR���^?ϛ�,�����.�K��NAq�^��6 vJg�����%���٧�����l\*�)(f�����M:���`Q����M҄�H�d���Z���?�֙=O���Fd>ڗݫ\�b]���PS�W湌�t�l��t��T�ٱ���	��F6{x���9/9�H��d��Fx�ؓ���ަ����e��`��6X���_v �M�)d����t�
/�7����rS����0'�`"l�A�:�~s��ė1���C>F�UjROgK��ae (����3��7!&>�7�Ը�tg��(�F��������G�3+o%K���
�{&�P=�:^U�e	���(x�At,���_$�2/2:�(~���W��!�l[r��^����·�!�5��3�5R^�k=���ΕǕ�'�Ok�[R�r�b�<�y�(ڡ����4�u_����]F��;:_�ߒ�D���cd�x�n53����qe�J�c^�c(3��J� ��ご�B�'X��.��e~��^����Y�2d�B�J}Ҿ��~*A�N�h�)#lf�����L2Y�Ix��;�9�%&�� 0'f���ĳ��g�\LNx�"Թ��MQ� �NT�\���"�>�+��{���=���A�@�=p�u۟}P�e�#ʪ$�j�ŕ�:q	 ��jφ����r���-�oi��H�7���w?��Mt�e�W�R��)R�g�9A���T���K�Hx�y�����b��݇��Ϛ94t*:��sb�o�~��ZO!%=�Ɋ6T�1�E���D8��Pl�-�9/����\���2��2N/��O@j����$SC�A�jm���4�ȐL�}�a���(`!% �+ˊ��H^��:Bj��c%����#����F݃�`�;ے� :zz������� ;��}�yOv �D���u�i��&�I���E�}�r�;�g��	o�b�X/߀�)=���ŵ.= ��Xn<ɂ��G�a�a���R\ vG�WM�W��;�=�A�s}΁���;;n��0��I�Y�*�l)
�@�ΐ���=A���^`q�_�^9A�j��D�s�����,�U�(۫���Ծ��hP�\�6$����-�(i�wg5ْчm�찐�� �|!��I��*U���(�t�aZ�}͡~����@�xm�����$S�s�Fb��=[Vuk1^���ɻJ�)י�"���_��ƈ�I'�3Ἔ��Yx��=��o8�+��~�	�?DnF���s��2$�o����Π#����Z�������^?�p�>�ʡ-�L�y��T���.ǿ@���i����J��&}/kArHom\�+tl��H橌R6E�D/�TC6�]?P��1�8w}�n�a.�C]Y�1Jil^1t�w1pFǠ��MI^I?��)����W(�#2s"^[o��,����xy��u&��Nk�����@�&b,wlt/:[(��6�6q��":�Q����{@B����V�<�����������C��4q�g�9ߎ�d<+�����pُL��NF)O�HL��@��d]��͓�@d�֊��?g��m��%\�?�2_h�ir����TR��Ū��	�C�жS�Iv��D�C�o��ұC�b����?ܖ�N�*�wOJZ>���&����IK�b�.8��x�څ瘌�]R��Ȕ�Q�P�v*��x���KPM"�&�\7�u�fr? M�M�U��w�^���	�8��W^(�Q0i;�M_Cb<&����X�H{6������1~�(Q����X���tO)F��4Ax�(
�/�ݿ�7�a@A!�OX�4y���L�w��1��y���"'�/7�|t'�!c�}̰猂c,߶(q�$Y�N'U��B�lOeV��������+��(��~�e4xN�k�h0�����[-'x=�	�?r��������$�?3_Ӂ�L�&}ɋ�\]�]-�HK�f�E�ó���`��B���̂@)�0x�L�ďwb�7Z2�`t��~��r£����������6c��9����ϐнy�T��m6�,i5C�+�K�ݬ�&��Vj�WÄ���P�F
%�1�����B�,߿�/�3�=���3J"�G�{���o@��#C�x�N�����rBd�YM�Ȉ�@��iˢ;�<��Y҉{�˓T��@x�Ͼ�R�fY�&�� �tli#W#��SZ����bjǯ��#��iPѻx��A$�+�-��a'�&�I|G=�jG�f��^^|_Ɉ�>kh�׺��r����L��"M���-geW�$f��j���3�6`�l�8Փ���ˤ�\�w���'�=5{.������J���X��ũ@���~5�<�3�5h�s�uSq�l�Z}��w
G�Ie������)��/�nԺ5s��MN�������m�n2�����]��Mr��4s��4��K֩J�O�~����h
��V�z�厹nMKlF��+�|�� =����e�agQT��t�f��ֽk�	W�Y�H�QoE���ë��h$i�Vo����c½�S��m�+��eHm9�LO2*&�xy��w��q��&ÂRL�~۟s����5���|o�T��`�w�1�%�g, ��eϓ_�*�Bp���_y֏�W�0�k]@)�Ӓ,U�<��j�'^�he�p�
��o3����f�C���%�1���lt�^����[.N� ���>vdߍ�&����˞������,�h.Si�8��v�aq�cS`�>����]�q��j�7ܜ����/�-��9N�c�����)��!�8�x�j���������΂����r�T8܎P���"����O�Y�R̗�>kR�VMW��ͧ���4Ar�����9'pN5m�ѹ�֩R�e���������FH���[�j��=���qIkه��-��w�w�s��*!����RA�+��j�!�ߒ��;@^�~���J=���^D\{�����e6b�Ú��hu�� ��(�����y��:-l�KD�JW��Z�3�Y���˖B��2�jp��y��ir��k����B/��J�Y!\�ß�e-쎯�PA��p󣀪�`�+^P`�c���K ���PkZ�� ���b�����<���Ż򢰒�-:x3rH�O�p�h�ޟ�V�� �la8^�"���K��+�b�Z�QY����{zO�܁��gIw�D�w�0���Λ_��G>IVV:-��(2_��DQ�`@\������P�`%;
W���ދ��\�]O����o渞L�B�"�9SL�^����$�����:�W�P�L[�'w��ɖ��FV�"����Wއ�g)C�G��3�:kKO�}���N�����?����^p�!�N����L�u	�+fi�ʻd8Ct�O����C9(Wuvq0�b���r)i|�e{��&=��7$B^�T}�������#�+'�ۺ��{�Pe�r�g=�~�H쇣��I�{�D(%oe@]3�q�\m3y��x&#�<(1?o�^�.��P
a�& <.�;gxP�-�U9�J�9��|�����ʢ�Ϛ(|�����I��[�,�I`s��H/�ژ�G��co�s��c�3�I���(^9��
�L@'��Xq%�B5��j�3�P�O7�T�(/��O�󕹚u�LE1�����_H�L���0��(�Ψ�6=�����߹?d C�Lͽ��X�#�u/��g�&��$����h<@�
iT%Tji��*�������E���21.���'D��8|�	�'|�3��&�˴j�$Ju/��:�X�Cr�F��EX	=���z7�y���`�@b�	z�;gW�����B���3V]oI�bisq�Pz�ˀO��ә�x{���tEUx���L�:_���6	qֲ2SLU�ўgb��g�Y��g\��)�}t�b����,��W�Ĵ��/�[��w��7<̡h�dC=E���V�aw�6��!�v?�/��f�ۜWU `7~�鉮j\��	o!�
lեs��TPM��d������Q�:�XI��74qy, <cH�Ʒ �Z�����#�'N�$z�oH62"�r�7�w�0��_]h�`��꽺  �L*�A�퍢_�Q <T՗X����1 �u?�a�3݉(��x��
�4�&�`D�7�Z�ן���P�o���9�h��@�@��  �/�L��rfՉ������`�ՕJ����?��O�A�}�4M*�(2ْ�DX`���bF��/�͔F�+���rNnc��׿���4�e�>D�<�@�@�YP(_P��Aa=���'�gY�Z�>׺�B:�Au#ސ� ����8J�'��>�M]��am��\�1@�hQ����@Ս �A�Aj���e�Lv�y\�X�٦����BG���}ǉ�b: ��8�Ĭt����_�$����~]�Ư�h���Ɔ_5鿹0�0ϱ:�����Z��5rB>���V5�M��X0Uttnl�d�Ҟw�3������KT��.�+�`�#�?z�`�G��F���=h�V/o���=�� ����1T��垖"S�Y��6���A�������)�4ռ�t=�9�l��ǋ���Moc��˝���c�/�[��]�y(���S�H매>��BƝ ���V�z&�2z��L��~��Dhl`vM�P���-f�E�2��)�*܆"Ŕ�0��U��_L�h��F�ٍ�]LN�F���@�����S���>��K���k`+�0V�Yt�X�����l�E�*ǂ�`"��(�a�Ր���2i���=���z�9�C����5?񗜖]V7+�TX��j�X1r�.��L3�����Jʶ�M�&9�Zk�QJ�Ҙ�.?IX�6�^'�VL�K����3��<:(�>o��^�G_�U�Ȳ���s� ��Q1:���H�H�S����;�E�p�g�ܝh-<]O}i���&���{�]U��]���sl�2��MA
�����N�,y�t}��gA�_���� ����K~P�Ѝ���e�<�Y�T�v��9]�B^�߱�F���*��kd� ��enB:�mDas�@U�hCb��X	��R4�9�!5#���_��VlC�iی�hi�챋�Ӕu����y�"���/t���ࠞ6@�.'��.�oQ�I�O�i͈u����,6���=4���o�_��a#�ȃ�/�a�鿌� V��ǿ����p�r̩��,"��]�RH�/K��6�8�����P\��H�=���6:q�{�`��� S�z͵sɣܗ7|aq1M:#��Ƒ�ە�Y��,*3`˰�US0Z��;�E�0�m=ds,r�d|7�o��M����^`(@C��ߦH�а芆��I�wC�,��&*F��\h���M�VI�M��Y�=��#.�X&�3�p��kf���AM���"_� 0tF�}!����Y�Y^��T��5�K�>Xū̏n���Ʈ�|��/��R^�����?�FHI�jR�DɍY{�� x���[��|�$�/9d~�1^���[�šZua�]�����~nD��23�,���ڒT]�rv�E|��8�?�
�Ze���+�j�/��{�fo�Fh�Ք�^WDNk��÷؜��c�C���B�D����d�P������`��YA�2���/R!�Y��5`�HDP�] �I�yV;�}�#ߒR�u|Κ+����?#�|B���6z��i��^;ѣϸb������E�Cņ�bs))at5�MD�w����O2�UK�%��G��~g�>E*�d�l
�8d�@�	Xf��H��L	7�6�Zεj� ��3=y��92�C!U`V���%?��ae�#�"MT��Y�1��J���ù#�������Oֽ�)����e��8ɵʠQ�xk<�"���u�d��]������α Ņ�N�QX�{�ޯ!���Z���&��W6;�i��Ȃ��ֲ�1����"�:�g���nܽe��}�1���@��+~�ЖYZx��
4P�\2����7�d�y|I��Z�ms�Tm�W�ѻ �QGǠ�Y�O�%o�/^�m���:��E��{�e+�fX��)��,��Y\�k.���{#�]e\����XCOO�X�%�+���z�Nb�b9��l�ȋS�����v)�6I\r�kB������[y<
����d#�E����#Ϫr��o��mb��i&�~�R0�R��� 5x��IҺ���U��A�$ ��v���:�I� �})��J%�[�j?�lv�H�#R�t����t���q�hj��Y�|�#��ޣL�fx���ގN���u�K��q����es��\A('�w�%��?�ql���q$�o��ե��uS��^=r�#�r>J���z��ϙ������wt���s�,�w�F+Ѽ�Os&���/����\\��8G����G��(	�X��>,��	=�.|kr|�Y�b�y4�k��M]�^|=����V������o�<�UH\@+N�SB�د�u�c,W);d�N{�\��ND@��J(?�h�~�7���Jj�Ξ�y�!?2aQ�}�'w�#m���a�Rw�Lϔ�\.Meh���Z2~��HQ�=�n	��%�˕�q 8Y���R����3L�?�n%R�<�RM���S�'o>�����[4�Gi�{��,N��hg����.A�lP܋~b?/��ŏY6�,��0�����)7R�b0�K�^�P��^������i`.�m�;zh�=`[�W�Q�g�13��q���8��Hg��yJ�S����V�&�q�B��x�-���&&��[�F�[��mk��!��H���w^������Y~MF��H��E,F��)�  ||e�or�rr/����_
��|����Q��d�Fe����b��W����7=�������^��QKp}��v�%
;?�t���<0�4��f�'�P�n:������w/��cec�G����; ������v�R�,����̦��_�q�/#"W5����QsUs�N�4����eyN	��&���R6�����pCM����e�#�F�͹�{��#{�o��η�II�IS�S�\ӵ	-,C���v���b�w��_e4�ɻ6��}����-t���'�'��]ͳK�Ho�0H��9g/��52h�N�D�7�lP͔(�vA����@�33�J�PWnvJ"�\w����8+	ڋ�� ݠ.�� ��&����̑�nA�`�H�?^{6<�H���=�`��'RH�Ue����t~>���̟ޫ���3�ӽ�Kv(�z��.B_�F�D
3YCLS�X�G=#iIF�r��B�����\��Ժ�f�LV�t������^ �Q�
�"Ö�\�ӂ���*�?S������b^����;X��׫���:,��E����*U}�AM���9��q��fvHeV���!f{vCX�#�e�7������s�5�US����
�Z$�(5�ڰ^IY�����q��4w���K��6�_p�G���'fn��T�~u1X�MM��ݶ��r��ST���`�#��vߖf�zhtM4��	M���K��
��y��Ԋ�R����R�����tݛL�/e�k���Zp\yF|��}tY'>4�טE��^qW��w��۸_/��3�0��.d:Z*��q��i��5?>8���c��\hy{,�)��Bb[�,Ƭ���������-�������7u@w��~�chs��Й���s�*v&+B�WuV��))q�h��o�� $Eg�}.�����.���� _���!
����c��I�.���C����V���U�f#ZX��ek+���������68/���h	�
�dq���:�"5�o�����^�u�&���:��-`�ڼ���$�,nD�U���6���z'����M���ƖpOF�����",��Z����ӣƁ�/S�F7�s���9y���p�����?
'9�j�q
Ĥ?�Z%��$�e�D%e�2o��Y��"�y�S@_�L�:��.7X�kbv���%Dq����8�H�J��Ǔ%i�e������Rp"pj܍#J�X~���%��-�t<�;�Z�u��; c�tNᤫD.��ۊ�Q�x��w^f�nh&S+]�|��Ɯ5s6~�����^�b�/D {-���cb����g"�$q�n7�� �ߔ�!cݟ�[v��>I/IB��.�f��nF�J���`-��A�Q]���� �BfF�M����z<W!����K��f�#�n�(��$�Ͻ��ܧѲ���-i�7�j�+�v:�"�s�tX��e��x�X4�u1�Mq�}C/������e�|�u�z�_y��G}/�r}G�Wd�#<��#�Bg��s]	7k�����m)X�A�-��eeh�ڰk�ѝ��x�8l��*��5-�h�r�'o�,���%W�Ը�g����^]�F<�]xN�	R�Ή]/A�(�;���Sld�(��l�6b�ǚ�
���"䜻�T�|�A���u�]~��n��C����P�)Aé�V��i;�V�'�7�����f@�l�����.)�����;|�|0�&4�`S�/���g���������+ˆv��i8���}��e�8�P���#��^i�C%�{(��\��Oܫ�RDN�r�u8��:���(D�j�W7��V���]Wz�Cq���W��uaDb\c�}]�}lem$�D��33���t�Yqg��Q_E�ϖ���>��&���s��+�n|�g�tyؔy�)t�'4$�x1�m#+Q�s�mwcM��y��^�_�`���Cd�S��y���7��`������}�%w���s\��։� Eco����W���r/	>��	�Ҳ�A�*%$WP -}�װ&<-ŀ)�*6�Yi�*_)A�4�7U�g��T큳�ɓ�ٛ+ s����>E�n`ϔ��U�99��2����2K�?A��of�g�亽��0��6� ��KS��u�&�c��}�F̼�S@σ���ei��Kj7���^����^0\�T�P�	a>�|�M.uJ��)�N�i�������� M��,_1�)Cڽ��8���Y��8�Ί�z�c2-���]����=ு��x��ᇖo�$3�v��->|�Y������/сw���o@����]�"��掛?��9�E������UQ�F��<�IOрy��j;>͞�#~��Y�7T���KL��s�)�+J�iIg���t���?�tf����%��z$Hb#Θ�h�vr����m�m��gȘ��NrLc��������.:{�M�Ä�����篁��&<�I��f��c��MI����r�_�\X'��iƛ�K�Q(YF,&�:β#JO�����Y��ؘa���Z�]�X��܁�.罉���Eh��"Hj�I}�E��r� l:t^���	2�S��ߜȐ�[�$�M��nՂ�s�J���S#��)(�� {&f �Zp5����*G(:�g�xS�6{)snNŖ�/l�'?Ǿ��C�U����$.�=�iɭ���F�@�}ɗ�Mꍬ�)�8�)~VN���B6������5/��:O� �G��c�q�4�}i.�V�su/�g�vUs����.,%=�����Cd]#��u�.�BFx��]�-�D�a�[��BU��䐚!���p5�q܋��/<M{8m5T<��vD�61���º~)(���o���k�jȇN:�	ަ�a��u�����^�rG��L�B;ϪK���0X�/ k�v��B����XPv����}��!�kV׮�-J�؞���$��$'�����T��J1��0�H�4%��/��S̭����2��17qy+����T�N.Z5�!߫�Ó�}���g���`2�8b+
�|4��1r�#6'�c�JH�O_�9
�`�Zh���?�7� ��XdŒւRPD������W,]Õl�f~�ٖ���QL�w�"v�x ��֏��4&-*-pS��z�:����=�Lr�i;�B��O(%$G;��o|d���.ג�JM�Fː}:���ѕ�mu2�'�D�HR�Nӄd���:!���̈3�6����s���ߐ��t ��kK�US��p(��d��	fM���yʢ+D���b�#�(��`�!d�����E���b#�6R��]�.N
��r"��×��=�F|ѓ��}c
���px	��kw�����y��\�;�����kֱm�� 3>x���PL�Y����l%���Q��v�I���&�#����c%�,���\ ���jO:�8��u���Ν��Ȯ�XB���KG��p��R�+��
�*�� �m�j��e���!����hh@3�?%��]��?�X�=c:&�NjQϚp���D���_��O8�l��Kҽ��P[��m,���n'���n:�H^����Cᴔɨ���?���z7�WR~�q��M�iL����44�2�"������=�3�Rۆ"�U��Tk�};K����el.�������>�ƫ���ZL���&Y�:�'?@yα�K�*̗�r4^`37��V�^��"E�Ʃ�*�
�ރ��o��S������l�>i#��Z�&�^=�a,Ԛ��i�o?��sR�B!�A<��n�����޿������(b[^�ur@T��wЋ��r����]9K�ip��cܴ���CƆ,�~Ւ�\?�"�
���4��1��\�#B���j;ku�a%&�v�(H�,v��@��iK�aD�O���C}�O�������/p����/�|��yK��[��隉]?с�WJ���YH��C��Hw���W�+ϨDF/�z)��=7K`r}t�TD�����tp�v;��|���h�?2�_r�a5	^r�hwo�����V�0��zb�s��8 �'�EIC�>�f����c�5�|-��Ž<�{P_&��t)(L"�ͥV/a�2�ef"b=�U�acɴ�YG��V�X�-F��>/�or�׏�F�[��9;鬈h��h���Q	�8Э��O۪����@��(�#�J[V��W;�L������W��{��J�r�@�t	�Y�y��&� b?��;\4�AƋ<n����Qx�FP/5�����7�N��y�D{�z�;�:]�+�qMg�sYӣ:�x$.m�6ꫦu�̐3w!�� m��q� ��#f�U�@�5��ݜ{�!v !��7|�̤��M���_�΋/i�~�$�j���o¬�E[��]���P��w٦�����3u�E��šb����%g��c����Z�j�O*��~,�:�?b#�������zhFkpP\�#b�����D=�R0|����YYR�ߞ�OĮ��)i�#篲��V.y�*4���&��=�`P{Z�-7�+���U�\�䇈E��eY�눯?�������
��7��D�tĠe��b��k�T�s��Fܹ��z��(]�]iDpN�)?d�wQ�"0dR��CxN��5�O�^T�`j�[�1u��q��nc|�"Q�Gf=ߛ8�J�5�P�Z�+��z�S�^�KU�MKY��`�C_�[C06����X�n�P@�G5Z�A1n�Ƈ/ʝy�B�#\��.b���@��FI�A�!��+D��>ڄ-���JW�0Q���9��sY������p �Y`��a �����[??Ba]�@+L�t`�ڊ�m�p�eT@D�>�ƨ��G�i�	 ��ق���J���߮�l�LU9�}<��&�7G{�936��cY\ �*�3�9��7��,�����JdPO�i��h�QKj>�r:�ѳ^/�:����цH�����_>�6���Y���ofЀدt���X�x"K�@��I[��2�^���r�Z�����,X�����բ�A�Ä�^IG�_��V	��g��"���h��I���1&K�������e�Xc�~5�	�
�g$��ġ>�OW&@6�����So����)����M��[$��8���ۜ�S&��+>�h��h�bޝ��ē0��t"���'�T�Rm��U����/�t֏�h��2���T�x^zp����"ˠ3�������o�L\U�ә�x}���L&�木{HM�V����i�=J�e1�W�6�{H�^�\U\w�u�U�o��L������mD�>X.��w3����۸��V��>���s5�xU����hPx�n���h�t��ql4�;>m�� �` �����=��ݕ�M
3(ki�%�^�z��x�t�f͂ub8J��ǣ�m����a��T!mW��̾/Һ��`3'm�39h7��Ts����|�I�e�؉	�7Wl�駾�A��uZ��t��O�Ce��r�p|ӛb}��@|�Z�� ��<��o�):��Դ.�8��'2��}'v(�����p�o~�V#�g�DU�Q�A/w�I������-P=�=�� j��}���N�{��!��6r7���yzL)4��yR-=:`&����X&���0�������ۊf���e/@rO�j��t�n�V��,ُ�{g�H�����#qNelR�ᮩ=s7��%B�#����}a��l�{��ߔ����'�Hu�B�L�"�+����?���Q���)'h�i����[52?��o���9�G��,�P���\�{4�`j��sB��+�� pR@{�����IUX5$H3����Ug��oꀐ�Ȗ��Gқ�Rl���)b�qJ��@��OTX8�G����;���*�+�	��`8A�a@D���*��Tk�k�Ē���'��s�P�`�q��#oLZj��M1L�@3s��8��������@���ϗqWs\-)�r��}�!�A���e�{�hQ��>.i���%�K�Ye2��bSIޟ�c&H��>?r��
�	��?>��6�������st��i�6$�����0C� �K
A�Sdh쉖��E��A���������%,�<4��F�P���EP�����x�����ZU��A�p�s��V~�yp�/H��X�l��R�ƪ�a��,֘���fpSÅ$s0��jjZr ����\�jA����ʜl\�!W�w�\O��j�}2Є��	6�ܜ���NN��tt��s�Ɗ(�݇�R2����4���1jr�YK*�e�8f�����IC�8b��8����OY6_��l��7=�@+��Ń�v�G��C��b~ԫ��+��O��*W`�	�Z�/K6��{�	G:�< Cz	"�;�<e_��7l��-��k;8�oҀ���AV%~��̧/��)��^D��W4��z���"�uõ���g6��(�9�L)SV?nc�q�\wC��_$�(�N=Y�83l*����{��L3�>��4G�0�$hDzC�J����Z�*}}�EN{=|�/�Z��2/�Ֆ)g1�Kg^�GJ��1r�!宑h��]�W��R�k���7�!E����+g|:�8��jn�_�R��T���?�Ӿ6�pR�e�I�U�%� �����\U�!µ©�+LZ��Ϙ#����x��i�;��F��wMzq褫LNF��J��1�C�wjӄ���?��Y������B�[�'Q_��K�O-)3՛%Ͼ���J�$�]���%�5����7�k�#׶`|x� ou�P�9HW�^Ȁm���tշ.�� Y�,�f�m"����/�$�U{����вrx�ՑDvS��e�y�dW�9���}�W����Q ��k'qą )�>g��V̈́����<��B����CR@,��k6_����C�4���JZC��6�74��E��%5�����ypU�+�FmX�⟩3STqJ�ʎړ��l.�'֥u���@e	`��~�uEs �PM�wA(���b���lt�%�6�e�����\�t��%=]J!h�I�������2֦BF�G)�KaF6�5����_]�L�r���#e?��I�"*���j�(6�b�V*Z[��!�r��ι��7����I.8�-`��9X=�:�ME��Ԕ%#
2?�6Q�Y�5r���\ݔ���oJ`�e38,O]�:��S�U};����3}ZIZ�QN"q�tqI�	���VK�Q��*����0�2��\E��i��=���˘ ���96��b@����-��2�����X0�4�O��-� 6J�b�2|�
_ DP�(@^�]�u�>펂��s�,�+�NZ�	�澿~N�,}��)���O
f��\l�5F!�GZò�Y%Y/�O�CW����{-k���΄���U�|<��)ބ%,���ʸ#K`�鈽�VC��.�Z(���|V@q��3����@�|px�S� ��<>C�V�w�C�fG��o�us�\Kw�ĩ��(ʄSq! �.�Q��|u�_��;鲛E7j>s!rs�KAc����-���y3�HS��+��(���)�X�[_\��D2ȃM�&id�U~\���]Y��%��%]���;}	mD۷or^�B,6�直����CF8���?�_9l�ppG�%��]ަ��c�Өd�Ԙv6�?��0�2!kw!�Xd�	+�?�X�/��zH2�m���Ԯ=��|�ȅp�}�.2�-�_���'���/?�H1���}�)k��u".��-���A]�c�V��_ٔ�o�]�����1\��:`��{�d�<F�)O�"T��0���j�qk�ִ�r4!�$��s�
&�ZDF�h���  ��pܒhY�ς�@u�HR�C�\�\Pk�w/����F���E���ؿV ��ҹ`F�)�܅@6�uҥ ��5�"�X�NH?�c5l.��/������L�=�N]j�8�%���?ϰղ�U4b �vn�Cgu:����b�ڶ�#s���QI���Ic �B\�f�1Ν�+5������V�UYo���cq�0�%��w������ih��?r���۞[��W��%���ĜTT�׵���%y�Z��ۮ�6�.��O=A�>o����!d˸z�������{��\�"H8>�J�fo��Pbj�h.��c�%!%�H�LnX?�����a�ǜ����O����N�Y��S_VK�c��Ht��?��������/��u�H�<�^�\,������'�&�P!c�f��e��Lrw�u�[փ�h���܈]ц��s�,8?�嘼}4R�S��@Lc%|P����*l_!��n�'��V��Eتn�d�`C���Ϧ%�m�b�� �w���IĊ�,D"DoP��l�g)����N��ػBQ��t�5��$��`�5W#z)�_Ǭ%��"Ŝ�M�,���lp9-k�-ggaR��������$�����6g 
GJM��̀t��w�a��*�ՕgW=uV-��H����Ę�ޓ>�2#�NN�D�ȸݽ��i�ݻ��� $Tl����b��Ur9V����h��H�=���G�-�T>4�՚��[�O�qD��`�
�!鏜�DV��/c�[o!�x�~�6f!�8���P���@��ei,ݪ.ܻe�V�F3 |.3�鷊�������������JD*��m��]m	���ڮ`����3��A	0Ƃ�k"�)y:����0�������̍����V(�?	P�0)�|̮[�Wv`���Ϛ�/�8���� m8�~�2v��7&{�Ϧ�2�����7�J�A�4����%[{�$$+���['��ש�n��F7ɤp�z�h�Pk�A����&Tm9a�'���3�����[�E0?�=�D�7L9}�.�Z�.?�|S� M˷H!��l�;�ЎM�l�L�Z���82���S2z·�����D9�)�C0�!�C���T���]p����W�S�*�M�����<�)�ˆ�/v��PRf�3�&�p�=�Ą^s�ƥ��h���u�8L��Ux��/�\&p��;ஓ�� �Eef��Ję�T$�gC�9h�'�*gWT��4���R�}#?�7�8�@��1�{��`
��nR��� B��X���h!鞭���Z���=�ۘ,���8�.�gj�&7�����/�R�F�c$�'Bm:Tq�!��q�w@
L��I��C�ۏwh8RgW;�w��@\Q)��¡��=�v�_{���$�n�!~k���o�j�� �&O67 7:]^K�
����&O�%~4j��%b+�Y��B��2}�Yj������_���w���dJ�Ύ7-u�}!H��R]���B��#�S��3Vj�G���H��Hv���M�m��Z�5]�����Ov<�k�əhHX�8?�U7��`/��V����װ�0<�u�S�r�4o��B�ؤ�H�F��g�����9��?j��%׉]�1D�N|؄0��H���d.�Z��j�+]�o\J�e�ǧ|�'[e�u<���W�7�.4����f�\��߀)k�rГ#�� �sK�S�+�
q��k��K I�O�ie���v�׌%��~��D�����]�4`���{Vy�2�~��XU8+g����5�j��2Ϝ�k��Uf��_J��PXi���#�u��Ф·�r!T_C�%�Kȹ����ڿY燍zR����[O�ۃ�6]6���S��2��ezmg�m���w�Q�E�2#�`��� rIe+N� �[����o�x,s�lh3��R���(��U_%�?K޵�v�H�<0�Z��U�-��5� ]��z��]hex�j��;*�zZ?��4��è�?ð��aԚ���/L�{Z��J�� �BW���d:�SvE�ؽ�:��a�Xd�&�D�,xK���P�^C*Rdi(���p�Hw�Wڻq���2fe��ir�R����\�9�-(����h����S�_l�����EwPL�@D�]�D�6_*�=W;R"�,D����D	5-6Ԣ�3^�:�8FN}���d�c�ӧ�Ų)�.�W��5_���6�� *��8�!WT��ܑ|����L��24nt>�]�g>�Iz����1U�,d �n���&��<��� 7ǥ[�*-�v����C�q[`j���A�IX���_Ì�\������;ޙ9b	aMjG��k����HVާ�N���Qx@ُP�x#G�M4���_:��JI��˗,�����x�Qu�?�E��M�`p�(0��:.���5^�B�p;��a�3b���F������o��}�q٫ ��:�b�8u�$�-��La	N/DT�V1!T������'�y��,���)]J�x��-��.:�b�t�Gt�H�k��{0Z�H�y���0�w����N���hޱ�E\w���%e2�j�{�O���xȗ
U�\c~ŕ)��;�((5j��'�>��l��.���{<|��{���qD!x�5��N<����
�k2��\��U��pm��)�����&y}���/�J�6�ZNFRkd���_�P��?`��U��Me��}ٮu�g*_���ؘ��js�P�k�LWܱ��;�+ײ.-ϠR�	h�9��.� u��\;��֎�M�߬E�����b\���K˱v��k;������ ��e�<'�})�Wj��� u5�ębV q����U���C���O^�p�_)��[�pj���x��s�u"����V�뾻��u���ƞoɈ+�+���{<�jC�&���<�5��S�+�&QVx��[2�m��+$
n��l�h4&�`d�?�۞MՖD
�)�jn�W�Ҝ�i/8��|"��hS��1@hTSu1��% �Qn��+�4�ө5Tਡ�"��T��~�!SV&ة���Y�0���u�I���r��Q���Q"�o	\���ٝ�\*�gcĎ�^ �������r��^L�X�����*,1�b��?bWb��9��,���w%*M&A��W�g TW9��aHϠ�ť]�Z�]ls��QذSj9Z�b�eG���x����"-W�g��@UQ��BRAހ�1�?�q��.]&��ֻ����4�t�展\�2B�v)�c�cIz_X@[�,NbdY~�ް#O�N4�4Di�\X�K�X�0y�/ژ���Z�u���'9�� �w7Z������h�6��GU	++�.��*L�U��G�M|�P@�&��,�%�����0�'?�0�Y�-�صZ�Z\4{�J�%RDA��CN��h�Ԥ���-u.`+;1��:�bTx���|�4W�J����C�,ց��s��+�A�f�p���;�ߧ)��d���U�n��7jP�-�<�)�
�pYKn�����$���H����>���7��XA�i��>��9�-�"����V�K:�i[n�����c�i5�-��^X�hOJ�'�~TO $�]S8Q��7��$���#d�u�qri
�"ʇ�B�`U�H
Pu�����qaTY�Ѻb�^XM��}`�
ü�Db8\���ũ���G %C�V� �S�NL%{X���K����x�x0e|S<�����]@�Tj|jN��-�49SX�_aZw�Үyv�	��VMm��s,��##@#i�����;]q���pӰu�'a�g���+ʲ&C��A�] �(�	�y�㊕ج�'Bޜ�;{&�&�CU- y��[�>���&Ԁ��	Ģ?�s�^���cn�V�dـF:����2�dEyޒ�wH���Zh�JXA�Hꒀ��e*n���"�	��M�&���lc���PCcІ�=������h	�$lO����-\wܬ�/�c�N*%f�nQ.��taX����V}3���,�L]�AN��o/�7"J&�g
�:t�K�wHɱ�3yJp6/�K���F�ĝ���Kqj<	Zos��}��?E��9�RF�l���#�i�{'N���7<�h��]���~�c��C]C�H��va��D��g�h$Ӂ2$8����S�@X�m%�O}+�Cj��^��X�6o��P�����B���W�Q�H�9�ez�`"Wov�T�Gtx�8Q�Q��S7����kL��j-�6�(F��Z]���0�9��������(�&Հoeb'��I:������N���\լUE���BwxuZΰ}NB�2�Dh�S��+Q�_�����)E-)
$��m�G��J�)f/G�w�V�
��^:��Ļ��B)x n�d9�l��$Y�]����c�>�=�����O����Pre�M���W�6�J��`�mb�Դ�b:�}�-��|)�7�+�Y�d$z�}�,���U�(a�- v^=�IÉ��GA!�����V���h��x��L��p���DG�v#�,�f�#��m�v-{ڿ�`��m�jH 	�&-�� ��V[�$�T���шt�fJe�e��\1g7�CLrگKØe1�H$�ɦ6|��FwS�u�reݙ�F�Wx�؎}ْr�*�+���*CZ (��XUW��ҹ��vn��W-6��W�n=Jؿ�^Έ��k���q��69����2�6҃��v���	9Z�ET��*G�u*=K�`��$���!��q���È�)!������jˤkʶҖ�;>��zV�P,�T�ү�%�dX�amqx�ǈ�0jF}��vDk3̓K#�n+�,"2������iE/�G�O<�V�qni<'i��r�7������R��Ͱ�50�d�����vUg���h��ӝ�S<\lb\�G(
�)�o�L6B��i�s�*\�&�R�s�Y��� �/m4�^�+�!�����J��lg�u9�>�uQX_.Ѹ��l\ي�ӂdҼ���ع]2E5֦��Z�K� ��|߫�Zw�������0w�NW��>�"�t*�M)eŲ[Q9V��X���Z'EO�jn��_C���_��T��!��P�(��*����)+g0��e9��A��w���+t1�>��_e����̥k6Z�o�^��+��8;��G�����X�z���u1��:4�*`]y`�������[!�Փ-z�9&��12�S\���yH������c�ɱM
�G.��2U(����-��G���uo�b�iz�K'-�2wH�y�~��	Յ�i��~X�}�O�Rݹ�sS"U�����~J�lA���h��Q�1b��W�6���/���Q�|�TH�B�1!��KW~[~�.it������#wBV���hv<�Z��������K��.��M��m7�;���[�Ez��7,�_�eQQC�wd�6�/GP��	G��g�ˌ�@!��<*���F�8@di���/{<�1�&��__��q2A�]�#Õ�{�	�c����= x�D�y���y��,�j�R����8���g�glXχ|_�C�o���IU�{�O�ߋ�5�B3����U��*�.�w�>�2�B~�ӥ����(\Å	�zyb�$oRf+�eWN�FT�x���7L�ΰ��r7�	���|�x#����w��,6!��DO��>�܂u��T���z7�G�����b�Ĭ� ���O]xh�z���	�K.��N��OS�Sf�.95 �f��&��_.x����׻b��=��r��t��!�0y�0_�~7�WX?ǹ�<٭W��ă�!P�W�`5����I-�"��(oi��;*n�;9bIh"�VӜTIɴ�˦�R�)�t�D����}�@?�����h��h��*n$Y��;r��M������|�UIÐT5F`c� �Ψ�G#��1B������uy*�?6���:q�օ�cK�.T���)�.f�,$�/p2-��rG��">4Ò�c$m��'�WԤ��z�z&��W���6?�'�1�@5�w`��6���"�mǢ=]�q\^F6�lz�AҺĉn*�[2?��PF\4�I>�;l�Ooir�nV�#G)e��B�L��v&�뿥��gs��G��`��=C��{ߘ\�l�W�_$���
��/ܷ�tQLI";�!x��/��ҡ�S&���wuBK��5��Kq�K�@\P[(<�u��O;GH�-�Cg�=e[y��Vv�^n2h���67N:�����B'�s�C	ĸ���G�ۑ^@[�G���d��9C�;gq�����#��M\�	�����?�!������~]���)W������lB�'����ь���N�櫵����84�AH�y�����oloU�W)E��Հ�h ��V��h��̀��'b�+7�|��x:�_|�я��'Ȫ�(�{'Uo`%�`���>o�3���/�jT)�ي8�X@��kJv�]����7�Љ�ٗz���:)�^���y�kRS �F�ϋ|#r��Kƹ����X�6d��IԉUI��M�I{���������x�w,����W[۸��;��6��l�����"�`v���M�c�6*;�ب��a�T
�/	����y��3��d�,]r-*�O!�_)3������&�p�O�w����Ƕ�;� ���\s��tc�k��l��Qʡ�"6QN���N��O�[5��ƀ(�o��\�e�ɴ�@�������$[^2Y�������tcpp�X�����=!��$�Hu�����g'˟ )viALӲZu�B(;2�r������}M:["�OÉ"��L(�2-�6VHA�Kzݽ�삚�?�m�f4�:O5m���7DՍ��6�;�ٯ�W;f
t ���gh|rZ���rR�����) �5y1>O̳"��>D��J^Bd_��(hҟd?@�m��ą��H@gcKU� :err�8��5e�ً��908��ʴ�Ж�$G��{EM��T%�@E�B��$+��]W����p���ִ5=��]I )��r��ݓ*: o7��tgլ�-t���$�|��F�ؚ��"��T�����b�[�b��~�D��#�5g:<�`�<4����̐g��/�^bFW8����4��2 �&7[�26�ݞ�K+�8go�7�LQ���)�d~�z�+1��D�f��=^1�\�'fn�v�2��sg:vW�֕��t�^AQ���F��a�̌�]��} ��L��u-W�t��>�����vXz)�X��F�Bjϰ{���}[���ZZ��B���͠Ͳ�fH�l�3�L�/�W#�f��4?�X���|tM�����uMvo`�欈�`���0�cՁ�gW�_��W��,�]N"Sbw���3���W�[�ٓɖ�L�ݫS�AM�M�%d?�C�U��8׈���q�/h��P�k�w�O�I{�y���7� ��9����l���e!4�L����_G�>���su��N�Ŀ��і��p^��j�J�Q0���u��43h&���#:㻟�8���j�֢,0�R�s���H��U0e�.tYk���'"������"�D��[����ZJ�3p�7w�����gn��>��i᧡v�\��25u8�Q��q��s��}��V����/¡�uɞ���6sw#������R)��I5�g���!����C7��w���Z�4�{Pd�M2�����pp�t���&�-�`HE
N���ʀ��xd7^��0N������T�����Z�Po��&q�F��n���x �D(�Dh5X"ݰƕ���ͭF��b��LzU�'Nc\�p ���5H�­.�I��Q�cH�-�x� Q@k��8*��/��_�b��.%퐃;x\���Aje)f޿ou���|�.Ќpz����]UKE7�N��>�RZ���?��F��uw�Œ��x�-sCH�֬9�L;Ɍ�'x���J��o9|�?j�)%p���t�N���A�CdR�?�q0tW�=4e�Y��q�N�WIi�w��@��UPe�*��p�ӡ#&�G�e^﯄�?��2qz�Y=���"�]G��{�l ��Fh(Z�iǇ�E��9b�-���ua�15O�0��C�L@Xy�#`l���=# ��(�f�ۗw˙Q*ϥ��8.YrhT�Ԏ�N;�����E51n۹�>���ܩ�T�| FY��\>q�0��Lڨ��p�Y��*@&�4�J����Y�����n}B�v�0��t�Wթ�f�2|k16�?sq�&��B�ݞl��s9@��װg�����I�m�
C���b3A���4|~�& ��67�"���1�Dcףo)Cy�q�����[r'(�������r@Q��&�17[o����t����B��<^��������FVߌK0�E��#f%^�Ǿ}���$k��B�㡙%�}$c�(Ԫ�^��fEa)�s�b)p�&���[���F$��xRrL}�\�aP�U�^�m4�d��*�/c$I�hU^�Wb�gڟ�7����&;�}SXZR�)&ZQ4Zc���fi����u��*�ۚ�;�p�8: J�`���|e����d�V�}!p�P�v��!׽p5d2����ӳ��G�2���k�\�5�TP��њ<R�"�烠d4�]�x���hxp��ld>��)l"���Q� _i�1�$K��k��d={(L+Aʘ��rN/T`7Xp�%�E�ܕ���=I��_a<�RK��M{�lFL�
�-��BK�	HN�v� ���-!�;�_�������J�u�_��Rh��O~@�y�Mm�;%�٫c*�����62]YS{f�P�	����ߜJ���c���C�]�,��):�%��L�@�ju�w@��"���x��"r�V� ��}P=]������{���+�u���IQ���&���G�B���k݃%aN�Vp��)�]�U^wq��i�獃�Lh`.�<*�����*�x�ūA/>�]�)�ˉ��9�[�$����7�L�l����e�t��e(g~|�ZI+E���u�MQ��[`Tj��K���/��j:du�QmB>��0�1��L��e�-��ݻ(�ǰДn����9�S���y �%��&H�����y,��ƛR���^�m}�d8_���=����w:��J���Z<�q�}0��;�-�[�l���ˡ��[Cg�x�B���J����q�����\%�H#�*k.:���z?�ޅ�bzN�IsC�.�/�wl;+|s�r�Bu,_i�PL��}eQuzPHuJ|��T�gl��`L��s�q)K�01Ht�6�Vo5Y![no-� ׀S��蒝
�:��!S��(z�������JO�n?rR �羘�<���Ж�+�2b zʼ��dWU�W'�&3��}k@_��JlM���{]�`.B�o!�(�p�oK���l�U>���l���1�P��R����p��"�9�_t�7�|WaK�k�qh"�N�>mZ2��� :�M�xu�h̜����ҏ�e��Dt|�������*��N՚���&29m��_Y��^��쏹o��ъ.���*1�VG$^՗ٖfZ"�+�*P���?J�v�3����� %J��CO�>j� ?��Q�,�|e�'KY*����y�ۤf)S�=_&�]���7�X��J-��z�$h����TQ�R��؇��S��YW��ʿO,Wޫ�,��j�Y{K����?=���v�c5���4ڭc���W޻�`�8��ݠuGj/׃Esc��V�r\p��K�/"J���p˩��Si��%�
���#�x�QcCOTWh�� �W�;V�H3<��fjK��unU�[����-�a �&a(<�?C��]���/��,G$��I�Z���C�f�r� $Gon�8�ؐ�k����z�7�s�������Y�tp�W�6&�t;�CJ!Jj�HO�(=���^���,U����4#����vw?h?���q�]��;�ÒU�Q\շ���V((���P��һۺ�^$+
2o�?y��%P޻d�m�� �l%�E�5�'�Q?�W�k�}]"��N���H�y�����:F���ج��siT��*?cI|�ٟ�޼c���G��$ro�[��D�89��J�VK����.=��,H��F[@�	޿"�N�tg��Z�m�� ���n��k�8�)��Ta1�=mdC\�5
"L�]�ȶ�	2w�Ł�ƹ��"�o�y�\Ə-k�����vԀ�����l�pQ���*��@�@���5��b��pՑ�j�_����$0��B�ޮ͕ע_�g��'�)��|
h��^�e��7Y�o�m4ALy�;�D)�ta��Đ�K{�Qq^s����q[J.s披�X�I�	���I����.��}��8�Q���ؠ�tK=�ɒ����\��f����O����dP��?x"�Z~yw�v����3!�p�� |�ڐ��kr���;��l-*�z��i�g�Ӹ��]n�zL()��_�O�GJz�N8_e�����2�]��LN��QǶ�G}����Io �9�7����8�+̬��N皽�^���|�8�I��S=4e��	�vl�����F]KW������- -�:�_:����E�4�֢��1��q�d&�0�X�v�y>�o�B­�w�e�78>�4Ґ$��S{�6����~�$ҿ �N[��&��/��j�� B P�K���P�����a쓑��� ��|��vC�y���f��P��\.�,cw5#��N� J�t!ep�ZX� �� 7Z��a����׉�+4p�'8�AG�ѝ ��Ӫϧac�la�9C�Y�෉@ m�PAhS���SS�,��*܇n��6*(c�G����� �s�Cef�?(OO�X�����y���Q��
�S���-���M95(3�5�C�;a�=����Ú��Wj��U�d�V�!=,#�4(�{�}��!��̸���k�J U�pk�̣�^���9rXVCE\?1�;|;�	RFV���vQ!@�NA���d�:����U�я��f�f�#d&U�N޶�%���U�&P��2�d{	R��[1���h������������h��8���A�����$@����4m�D�9��,�-�q�_z���OS���奩ܹ��ZAO�S��>�b�)�	� ^��4
?6HۇxX	5���6������x���90㣕�J�0��^��3>�>��)�JkΆ�(�����ޥ�(���ޣz=k���=
�������#^xC�������%��gT��ʸ3Ӣ2�(+[F_�鸍>!��'��ZB_a�HV.A�\?-�a�\*cc�d�I���71]��Q.�*"6ı3�R7Zɭl(��N
�d��Q�
����L��r�"���n8�!������)F��#g���D������٘��\R
$;�&�����M�gs�&v�|O?�6t���[�ey�}�&��B��E<
��S��!��)�_FM�k�뾫��
��!U:�+c����DF_e^��^%�(R݊����< ^�vbI�6^�U�fM��_`o^&'�rʽ8���A6����`B� �g��i�H�C�ص�������()���1+|�wL03��1��J {;"4	�I�pA��p��[��X�~C�q˳L� �AD�nbh���`���.�8\캘�G�
������[�4��� )dOyU�EW�E&��p���7�.�Ջ����k�fޢ����e23S��<�>4&hYyk��<���Zy.�WD�PZ�!�a�V��R0����V�5�Ӎ=�d#���g�ωҰϒ/���YnVT�X�f-dĪ� �-^B� �0K�`�����������&MPeY�`}���&5C�!b��RJ�+)��?pz|mj}A�bF
AN���&�`��?�B+��0����o�
3Sv�}�:D�c	�bN�'�l]]�!?A��ŮW+��ܦ0^�kԺ.�s*���c&Z��	�>@�Oh�#o�O!��Au��cA"�������,P�S�
M��N�+�P�����u�}p_ơ+	]*x��R�ɪR��E���O�G��7�����vZ�R���>���:i���u�x�Z+ݸ����;p.+)H=�_��UQ�չ.��ʓ�$���.#�jNӨ��`d�:����T��=�V�RD'�S\��}�.%(��#ېC:}^]ar�;�2M����U��G�,,�@�w˔ A�GG�+l�lj���D���� �oϒ���ո;� ���)�g����KWF�Ŋ�E����1�\�X�|�QA��Ƥ����G
���눼��ߞ4������oBGO�ݳn�I���z��j��[�̂oE�[�Z�D�ke]f��;?{l�E�1@��"�F���F�ă��&��> G�*�sؾ� �Q[�`[8 6gr
�o��t!{;ߧl��9�H('خ���8Hf��� Lt�P,^�f"�t4Y�jޗ�ܛ�{�F�p�+��>��-���<����_�CP�{��"����Yڱ:1R�v��bhmc4X��p��/?�ٽ�gOUڥ���R���/�ˊm�!E$d.�C�ְ�Pp]�O����Af�xLp���.���7>�\M
�<'_�O�ԑ�#�:�3�E���b��/G�FN����2��6�C�R�d�&Пs�%O�T�6��Ro��Ak����h]ݭa���I�����.����U���z%��`��I 92L����b�_ge��֘�X�ϐ�F�v���q��y��5%{�P��T3�p��Sb���*��`M��?��r!"`�ٷ�U��t��7Q��2�v��%H��ӓ~x�eIS���M4A�0�_#q[+��5��ݖ�Ʈ�e�:N]�)�{�ε��"N8<]�)X�@M1���A��o�aq����'>y_@�;F�b���n��}qv\n�ք��߯�<a�ި����jF��WT�q��8-`����������V���RM�$:;�W���Vtp��cg���UrQ�W&�]�T.-Q��Z�m�#P<����%ֆ�-f�};�I�� ������5G�T0�ں[b�NR�
�D��h~į���n{7~�����'�{��ASż�̆�`Qy���I=~�$�V�Jwքa�|î�m��Z�ZN��	d��_9�}p�s^Dp���F�'l�	h`Z��o��T��]��%�� <2Zp.o�7~��[S�D���1����4"
`��Bz�%5��X����uZ�ի:$��/F�C��g��N�͚n��
��Ƌ������B��T	8�Uf�#�oF��>��B�c_e�������;A����d�9#[�hq~�U�jÔ�n���"+s�f�n���)�x��0B�W麶������d)�t�-�߉d���x;���9]RAl�x�.T�%���~s�֘6pM�!��Gό(���Q=Y�U�:?�(u��Y8/���q3ҚP��׳�$|�Q��d�:��lf���D����w�&�z����^�(�v:���K &���I��|���h=�!���i��X��D������	[��*ct32&T���7��(�;�3��w-�VO\U!,
ܧ��ڞ�f�{���i�4����ʪą(�y��T�QO�$��Q�G�� sٚ���eR�dv������A_~���ʱӦw�@@a�<��O	GSX�a׏iv ��I���C�E����o�!����3�cËw�Vë�{�����w������z](>�O��d\��,���pn�Y��lX��z�X\-ʞ�#��C��4K2`Yim���K�����@�̹�}��īLT#
�O(獁 J	3�gb���!�.������q]GP�<OM�޾�оq�/��S+�~�n]�	'΍�)�3DE��I�9�C�	�I�ч���k�t�>�b�/'�mD�kD/�;��'B�R(�Sf�a�T��x�����	#X�@te����7����� �|7P�e����i��[�i8��N=B�T)ǘ���8��] �6<
C6�E�X�c
�W�N�/!Ү�k��M�\	U�P�ӕmhdd�4Q5�}���-揸�6���e�@׫�N�%�4�3�zf��������p�䃶:�
�0��1A2U��)e�m�zs��	S��0<�Y�u�H�
k�_�)��7�=�d$���>��DHdB�f�V���}���oZ{�����N�qg'���L`���Vb��s6j���/������S�p��[�z�	hn-�7��"^�$���C�m[n�zN�ŏe� �6^`F��昁�WR�W>�O���3�F��s�$<Ȗ^�C��q�1y��j㿐��Q����[�=0XK�gC�S��^6�("��,S2�ޮ@�L�J<�Dw�l|;=�t�x��+c��o�G ���g=Zn�'�c�;�X6���o;�UxN��a]���-�[�2>^I:����?��w�הf�5SI�fE�<d�����5B-prv�H��d�Ã�Ć^	�ݦ��j�������W��y �j"�a_���SG�g�9�������ZM�������������Z�2��7�0�[cn�ǇjVCB0�~4��`*T���~}8�����h��m��T�R��{�³.�v홚Pt1�NhJĸ�U5���;(�BKw;��Zp�P���^�G���~	$|�f�f���S<�P�ʤ�m,��Ei������[A�>��,������ �|�t�[��*;�2B��Q!��Z���Z�%Y*ㅋ`ZcެitqS��cH͔z���,?$ ���ۺc�vޜ��Z�5��̝6�d@�#1~����>(Pö:Q�w%�E�	����
A3�ݞ�ҭ�b��<	y	��hl.q���)֌I�5 ��/C\Xl��OmTh�����b��Ǝ|�oj�P��!���漖�G�2=q���zLK�M�{d����}��Չ:��Ok,I�A�q�һ���YO�mSs1��B? ����S�+έd��T-_�]�˞`���u3syE��1K���l� �K���<m]τk����&�&��=���ȧ�&�.��!�܂*����4�����QG;��:(��z�-���5 C�Q�o<� ��Ix�}����U�,�ɘ���,C�z
�����ͣ��S��h[�V�Q���~8�Yh�d�͑<IGe�����2�V��	v=�y��;Y����C��:���H/9��Y�r�]�c������	AGN!�5������ŐC�u5ޚ���3L�+�Q���w�6��مh�~r���*��p]@枫����S��b�C��$���k���QN*�����C0F�𓏓�T�vOgz��ES�{&,Ou�
�b��E"P�k�:tG�~��>]~|�~��[��`!�H{�P��2�~k�ɓ5���`?~8�?Vc	���Habl�������J�mnX��=��Ҙ�U��əS�3�>~���\�1�IV�w��**�P��n��Is+]�;�J����Ώ�����#�\\���Jk��ZwiV����!��?�j�c @�R:�8�+B-�!��Y�8�`>�AR�	L�(��_���V���p�YE7����|G�� l�Kݠ��Fy#B�V%�-�бa�|�����#<�L[l���U+tG�	�+�T�0nPAw�ЪKF��=�t��Ri<�̋���7A�9�Yz�K��P�\$���7�f�ށ�	8/�c+�W�d�]�B`�IcZ�-n�;��uy�{}�v��(V"é)�9�ۋ�I�	�p.iY�)*�^1C���s��� *�(�Pv#��xn8�	����>�k�ER<�Y���546�B��d����EL-zǃ�@`�UɂT��B����E�J�� �s~�����^"�r0�X� ���������ܝL���i��YJy8)�or���7��#�o����������9���	��m����j:pꖉy��{�Ն�5 h��Y�,��h�����C-N�.���Q���YG'!�<��qP7 '�{�V<�U�y��Xu���e	�rv��(���7ԕ]�Y�Ɔ�K���p��\��N\w1�`b�.�K���o�*��]n��b��7*(\��1��Vq��A��.���X�:6��s���R�v#�5.��`ᤅ�) �q2�@��0T<2Av�R�И�Gv��I��K���ts8��*ƁE��M1���B�@��B�sVq�U*�Ļ:��7�~�Aj�a���o1y��&�U�(ƞ��z���G2�E�+�'��Yɚ�)9�!<x��a��@4�tl6S˨F�h�_�*yHd�Z�},��[[F7��d�ҕ1���̑�+6(����V�ؔ�ua'�9�@�g&�j8� ��2�藪��r(�)�0��^ڻ�Z�+)��� (�ܳd^:8@��Vn��A��c"Ø�p�/��2F^ᾌ�bi����`�5B�W=8�K@��P����j)�����t�F����?i��{
R�U��t�"遤���zu����:A�sP�����]&@;�8�����W	�/�a��d�s�E�x
J�~F�.�9�>��������������/	pQ�g�Hr�͜�i��Sc��Nn�5�
LhWZv�s�X�Pz=+��7겳��;��4����x�����'��DRuAՅ�	u�:+;���2��-��Qϓ'ZH� "��k1G��I���\���x�������RA�ס�黃O������e�����lf�*8��
1`V�j�<��RuU��.��f*L*cqڡ(�ёJJK:�QUF ���e�g�!�֍*q:ze͏@���R�/�0/�/�\㌍5��<i�_'��0���P^�\L��W�hs�F��ms�E&B��= ���촋��nC�x��>���c��*�:� ��\ ��;ዶi�>�.q����kpIF<�������Y{p�����{y�DMS�E�%(��r�L�\����>�@JI��Rݺv�o��"�ݧ#5~��X���WR�@F��);d%����WFy���q>�[26��Ӭ��'֔ݩ�?y�bK���5�a��0�Pq�����Tx�����﯎��ŀ�|:�������ux��
��i�
�`	Js<��
"�:Ȱ��9�ٖk��!�xk�%��tQ�~�7\x|�nkfA�i~h��9]Zn�lkx���I��o�\���U�7W�Щ�ǽۛ�����fp�ym2�oF�q�x�	2����+[�T8Yܙ�����b9"0�c��_���ag\���¥sR�Y�[$�ǵ�hS�r1B�y���Ѳe=|ص^u�j�>����!A]��/w�mO�},���I2�p-�*oĀ*�2�fL�y�k��b����+��R�~:AO�h�$n�|�P2�ݦ3���g\��S���v��a���$/2�r�u��xo�m�r.[�U�a���2�N))�������#l�-��JD�Z��ã�Q�}Mn��1�y`�/Sn�˅�q�y7-.Uҟ38�V�q����qT�B��� ߵ��׿NF��x	6�v���Ɩ����I�EH��7����o�{�)J�
�9���z�#^���3b8�"EqAM�^s��ŇSc����n�{��RV������G)
����a9���(@�v���6=j�v�������ʽ�CM�G�x��z0y����#ڝܪ�J)m��U���n�/�#P��C$����$����,�Iֱ��)PO��2w=s����}mr�$X{}�Rw�@Ĕ�x���J ����k�]��9����)��K���ղy�ܞP.�_�}���FA�W�e��"�հH�񌪗��7%����$x|��'m\��ޣ-D/�ł���)I@��B���s�� �f�L|�=--*'䈁 ��	`���ۃ���x�`�D�r��(u};UOr�?G���F��3�A3��=�	i_ɀ��p|��)|:�!����[AO��M��v��X�!��v\��H��	�=YD��w���D e���:��M������cK_�EO��`[��+��ǥ?��u����.��\]��)�=��<�H���DF9��	
&z>3}DU���ås֜W�=4:�PF�',ӗHkj����a�u����T\}XP���>�TVJ�&�f`f Ti	O'�����J�����sVI%�n��J�g��r;�p��W�%���b2��j�U�?<��1�Z�P�����e�G���BCDq�:��3l��f�j�7��p��C�M�`���~ֺV2x���:�xT����_p R�Җ_�l�]�BŊ�=�k+X�%�G�rl�@'f\�°��T�M��-L����ZEh�%*
!
lJ/p63V���1�:����n��<󂼣��n�eMo	�A<D�x25�i��3�xGs�7�������v|�Ū��������)�h҄�$>�����{@E���Y[dq�_8c�$��vzk���R�ؓ@ď� o�.�e�ٓF�Jw^�V=���>�v%Q/!yxIB�Aw,�6!��M��q^���i�?�A=�hb��n�X�B�T*]7+d���2����,IU���䒏�&CA6;cv����,{�>�C��W���������s��D�/QԎ��o!�8�{C,�%�U��o�A��nq�����I���	C�5^]����\��|`��U&eZ���M�%5Ev�Xk	�G��h����[�"0?W�-�k�$1`�l�f���{�f�7�&����+~�#��5v^����@�I���ʩ��>�ׁ��u���q��-�CC?� ����z�괆TX�@��Xͭ�EҢr#x��{T��3@���ڤ��nv�Vj)������`]�<w��p��d7Z>��Й1h�7!CCG-��D\�-��Gr\N�w`�����Bo�ޏ$��9�u��.X�b�'��]�=N��P�
�:�Bp˞�_˹؉��k�/a���;��w�I꣯���#�I\�A9��!u��_��"�w�����QJ%�M�8��������f���^M'|���R�Wz�[:�RG�*�lY%�z�\��.r�w����pwy��t�U؜>8��a!X5�Vz�w��)��Uօ� ��f�3d����R4�$P�qi[1J�83��Cܟ�k�@��g��v��B��q=0���F�#A�.>��!���`(���#��-�B�ַ	}��?ԟKXǢC��NF�n����~�ƽ҇���v��MR�uɈ��Me��8�j*�����&]^�`��*���p�V3綃:�_f*~�y�4�������"��5���<�'�ٵ��g�0���-��}B�E��d��4TL�Y,�j������Iy雱��k�4qq_���|s>�{��);�cY�[��S���D��
�[{�c�7l�������^����y���䒊�ݷ�qt,�g�7;6��F١��~ع��@~T^�
�K����j������BLf�5u�)��)rr�&����!1����2���b�	y�_�� B��������le���)�Ǒf"�8�����s`�ُ�a���3xaڻw@V��zh1r���}���|���z��ه���;�7��G���+(ij�k�X_��k-��a�6�I�_l��-WU�󕈤�:R�<���.I��{n��N ����^5����c,OW?��#h�x��}���۪��n'o}�
a,.���f�_���,L&�{-��)Ǫ��ڥ���5�^�"�AA
��J+5�PԪ���ͽ킛�p�H/;؃���Jr@W�Ɛ7>�d�f�k_� �E�l�a$}��m�̣-��Q���`�Z�={icP�7X��i�'����`�)�$'��'Uwu�8y�Q��T=9i��v٥2t�\��U*�\�a�D����9��a��A��'k�=ũ�߉��	`��H��\3T�i�1x8&@���S��*���.�'&���N� �yU��~h"�A�u���r[=��	��E��_$u����s�摿>s���mj�w(k��%��@�[��R��KS�
�шf�t��"�ʇc�QU��ߗ�̻yB�|E�~���T,�F	����#��O�w�DAZY���}�<��tp�Q���$%3ԗ�fO��O<�m16�|��U9M#'g~��f�v�N@��a�K��K�PIq+�~4Y�����+��3J�����'H̓�{6qެL�����x�\t�ҽ"�֖J�H�Х34đ5��s�E\�,���P�����2ߓ���}��ED!�l���;g�ք9�T��"�s��4#ٟ�cB�|^"�ݙ�Q���k�I�����^�\;����e�
����爤9���||���+��Q	�s�#��M�܍���4�����	�z��#������i�u�|Z<	��x�ʰ�FD���ʻ���T�#���2�9J�p�����i7y)�<�4��˾N��
pt���u��w�Z3��(������'|���2P6$mI!]Y}�ݰ~G���)��LR��*��s�²r�R���'�����%
K��w�3� {�i�<~LWG��.�Q����8)��N
ֆt�5.�O�3�R����n��^��˵��}��:��i��ȿ�J�J��%!��a��.���.�\���s2��7�#i�?٘���)���?�0�n`Kz�o��qw��;Ӕ)ZGy�e���\y@�H�v�g��ݩ�=p�SmB����v��k\���Y���'�|�V\�����[�ֈA���RAk���)��#���s05�K%�tyd���1A���C��\bN��cj 
=��������ݍ�d^UH�n~�m��	f���-��\p��XYwvV;��8���.�:SL�R9��F��|C�{�Fٖ����Ĵ�+,T�}��d�n��!ԏBee����Þ
�W�w��>82�a�#�*Z흆5��)�P�7ޣ�]�U���ş�%�	�vi9��8�m�*H���g��r4孆��቉E�xHL3�?�溛�i����k�j��w՗@��8���ʝ��$�n��?P�V�*���^HP��KIXV���1.}( P#�E�)א�+�CE���g���@�������K�ޭ*ԣ]M^[;��R�\=7���e��t�eW�uc4"��C
j�3���ٖ�-Xw���/��=�X�ȷ[�3*eO0�F�E��EMr�>�N�6��A�Q���z��X�	��>�� ��D; g>������ޖ��؍�=�޿*�"�\�Q�~�uM��]g��AL��!�,�@a}5���.T�F�_�>ާgX�_x^��%j�LgR�-�==��W$v�d㉴T�;ka�K�f~�+
sw�cf�3C)� ��S��FZ���im��Q�N[1@>*ݻ �v�d�k�9�����y�yD�Q��Pm0@���1� <ZKn��D��<�������x�b���T�K3侭V����2�m3�Ƭ���*�?g��N>�۷�V���al"��E�
9�Fގ�SC��mY��=���6��R.[��?�$����ד����Z�v�/�d;ӹ���d� *��!]GHhZF����v�'t�S.�0m��K�:�3DJ&����'�3����&����qd��>��N� ��E}�vTM?�S�[Q�������(��Pb��´��4�Jh�n#Go�RG�����:���e<��G�g9vg 3M�������k9����aE��[W��̖>���:�!��T�Ĩt��I�q~gކg�&�m�Q����^��dt4��\{��`�K�X,υ��s/HO���9	w.�*�9�{鉵��( LQZζm�h�y��f�X\�V�J��5�ox�������kt��2WsY�^a�ԕ+oM=���q�C���
0e�r����������7��I}��+�8�4O= �2N;���������B�P�욗�if���e1����fyY�[ɑ��3�K�-2��Q~��no�H�߶;M/��0��͏�3~ΡQ	|�W�#�yY�ӧT�e���cBH��ʪ��J��h��;�]����j#�s�68 �h�����������
��CQ0%Uɇ����S13�6����1v�G�,'<'��f�ţ����.�h�eJ�8�e��>�}U�JBiڨv�Y�I5�񑜬��!n��`t�N� ����wK/AQ�8%A�_>���^���IL���2��Dv�h:��m�ZU�ȑU���Xۉ2�(b�� c6��Z!9�賱C�;�8��OZ$6J�w�,L{�eP�~�Ij���z�=�B	8cd|w�]����j�o%�B�*d�ȇ}i�V@?���+����m��>�3�G�͑�.�]8}���5���Axsp5� Fn�����wv��)��f�~ ��>���>ɗ%��1AAu����(���p2���^��x|��ӛ*�@���\�F��N^��@S��H�9OwH����w���6 C�NH��I��#������גG|ϙaAl��B�\����WD�+�'w��a�hقE�\�|޻j1�^_�oP��&�>G-�"' �]@�Q.�36���~('�#��F�<���`Wė�(f�s���*�G ���B�#L��#����cj4��s��ySh�P�GN#Fp�������ӹ-J$I�J�iƲ�f5�f���gw'֦Cg�[�Dm��u<�_�/ $�`S�bHb��|+pOF�".��	�9
@�lcA>���K���b?t���d�"�Sӿ��_/�T-sW]�x���S1���['-sΗ̋�ˬ4�.�]�|��Q���T&F��r2�"�����;�����	��_6�%���}��4�F�1�DDJ�P�J���xvK�9j��-}�b`�7L�8h�Z��v �����/L�׿�Z��5��@��kB0u��}RaGk�E��(�k���mt���Ҙ����2�t�<ޯ��cn�l��$��>'����3���
O~��( eI�F�W�b��ӸGq&��ߦTɄn|z��Bz
���q�9&4.�;J����������%�Jk�g�>ox���MR�ʖ�\M	d��J���c @�����O�ө]+K�g_IZ�w�5���,ޮ��N�$�f��&��~dy��ؒW���?+�"� ��;���<~�R�	_Hxb�dEx}�%Ǵ�_�]rT����(-�i,)~�c�\�#K�J�M� W)�۪7z/D���jD���J��ǚ,�&F�[~/��:�I�������^����G(p_LX�?� ��H��0��F.�V� #ײh�%�:�~zbB�	����&4#B��H��7��Q	ec�+WC %"6W��<�{�(K�n�9Y_�m"R9N�G4SQiD ��y{���?ZA|�"_��� X�G$�h�<�V4�'��cag�I�SB7@�����X��n���Av˽@~uri�ɛKK��	��q��q������wҋ�N�.��x�9G��|�e�:Wok��ȶ)�%�bd�u�����4ZJ��w�aP��_���N7d�#�dJ*GG�ore'7ǟ��N��Lv
�����'��Os���x���]Cp3V�#ˏ0�T�0�kEn"�w�[���V�f���	v'^����B[��[n㵠	/wj��%��m�aD���Y#v��Y����ǟb�nĄ8:��`�/��ZN�=z��Zh/q�v�_��٢�Jx5�d7
^�Oۏ�$���E�oGY ��$�(�65���yΩ3�w������pWO�����1�s�[铷�\%��*��GV�rH�.C� 'Y�p"C�4[	�U|h�������&	��ytV����2
���N���U�T�\V��>[���t��;7�[�� �	��s\S���6���7"���ݗp{��y���E0�"7yٳ7�ą���Q��q���<(�Qm�$M���ڭ��M���7��y:�K��r.�'܁�[Fǧ���c����P��~5���Zk��D��EOGj����C�x���$
B��(���T���͊'��l�^5�yްP�z�;��0�Lo�W����r��R�f$F^���wث4a��#�	Ç�\��5�Fsi�v ,�d���k[��T�ǘ-M?����[f�ڑ����pz�9��J��w��턟ߧ�Uֱ�'���I�"1/�>Ƣ!��h�B^S�e�i��I��ᆙ��5dM,�Wx�t1�k�Q���Ųw_����O����Ewmtݵ�Slɍ���f�8�'�W�/��j�%n?Y~]���tUG��پG�t�ŉ���Й�\��0Y^���7o��A:<x؎&�T��)a��J6%\a�4+9��{NQ"�0�	�6W��1�UbՖB�8�As�=W�ڷ�|⡛"��2�,��F�ˌ$T�
s�<�_?�tK�w����bU��!�C4�S��(���.�?dm��}�Lyԧ�Y�e��K�k�����,z���Zd����	� Թ�h	2�&<*�܅E��aV�#r*�}Xm�S8l�tYD���Y�{$�K2��`0-}�9�@���_-�I�a������+�i�߶#��za)��(�4���ޤY��jэ0��Y�Yzh�p��@(��6BtRR|\��j��Ĩ�׉�Y �������Ĥ@{(���������@JO0`�{��H�:F��K�==�|��E�?�Gđ�jO�w�PZ�k4K����CK�$��x�m���M���À+���m���y+������j��#m=.u.�4�u��>��U���{�Wێ7i=�\���koy�Mn�+�x�rO���S��Y�����Jm�7ځD��`���e�q���\�Yq�[3%�[�OR��
u��U��MJ��}�k /���po��K�V��A|���k��;XC�`vM�%�f(&����n�p�D�Q'Υf)Z��ԏy(��U�������5�X>���J0�Au[g#h��L�x�z�Jlɝn<D���mT��6�/W�ǐ�*�T�CXY�����ů7��2�(��/V������j�1�U�h���� ﾠ�y�%��֫��qU�l�W�`�W?L�8@�#"������x�h-�v�m:"�9���<�$n/gJ�����͖�<�7Hn�n/b��J؉G5�ϋB�")LĆi@P�p�Z��%�q���1��Oܠ��4�C���
N�s�����um3���C�9<�������d������"�?��&T�F4����uۇ�є'U�<w�=m"��S=�Z�:h�_J�f��Ks����XP��bȻA��ި��W@<�<1�6�W�^�]�8/ր�i��>t�($]�h��f@�
M��f/�� ��]�fn5y�%�O:>烝\��OY�"�T(����о��b@�٩��V^�ϏMw���ĎX���4>eYN2��eEPD�������=I�-QY�U�G���R_��F˓D��=/�U���{��F��4N2}��θ�{-z�,�"'�����X�1�*�Vl I�s��,��s�<�l��Jbg!(Q�$����K�)L��s�8'�x�g��)9:ZJQ��Y�X��øv�C���
P+}K�]��{�̸�J����n5�i��.* ]pF���FT�`��}<>mQ����p���<�r���������������H�"Q_��
�`��M��	Tᜭ�T����~�9g��H�MI���Q��	��ѕ5}�#�(N��P#y�]�U����{�B�QG�ŝv�	Qj��˛d��tK���&�E���"���C����@���l�x
�~�w4~�c��a$���u�a�=�s���;���zU�:����L�1�	��A����q(��`0ڽ����"lF1Ә�6*}�"Xb�!gj���JW���/�9��9�k!�n[04>�� ���"�������>at�B<?5�5nw_�e�_��l��>�������u���C>;�G���E}���'���M���D�L=2'��; �ņX]ړn��pQ��L`m��[�+�<���U���|1�9*�Q��yx]F�'�c��+\���:��</�A"l�qR�r�M���=!&n����"��m���4��j!�j e`;��i^�������鄃�/7d���H����P��^qs�O�XylSY13�fTG���Z�.�v��1�5:	>����YL�vr�%��"�M񸙈��51�,m{7�a �o8�t�ְ"�Q�Qlb�'4y�aMzт%*�Vl{�/�ã�����W=�F�����Z~�5��8�q������VDWy���������p�b0o�U�E��b(���h����H�+����@I#ea�u���=���u�]�l5�����z���Y6OW8:"�DS�QӒ��k`�ה/ ~z��^��z��%�6z���5�����|� �%���g(sk�`��q�Z_�0��1�ϧ��7���?���ZcE�<`L�)�|�~��'hw��|:\^��F^0��ُJ�~�Ju#���j���*8��~�mi������߅P�����n�^�0U'd�(���yb���?���,�L~4))L���7�߸5�R1�ܻZɴ������#�m�T�2:�_�j>��Ш7P-�e9�e��}K�=#�/�P�g����Qtg9,�!v�ŇF�pV�57s�[�8^&�����?���s����ofUr���u�A�J��O�����א��`o96���C�y�ޜ�&+3��.7����59$���|Դ)�<��9�Xhz��[����k�S&��� :���ܣ!�ź�tcc�-QkZ�┽lk�uF���C�����Y���r�.Yɝ!��h�=,8q�U�7�E'�m�4�
4ށQ��T�%��\�j4�r���˸{�Ƨ�(!������Z9��B�#"'���w����5��,����;_��o!����j�����1��9�/�E
P
��k�׺�	��1��h��x������8��æ��C�Uc�Sqt+�;��
��� �����z����̩)_�ld`ϖ()�Q_��!z���>i��XǢiwP��Kb�K���ǯ�L��M�rN�3����0͑�b�F��7�\��!,�V�D럍z6I�T��	��m@�ez�Ÿ"�/��4�ux���!� sً��L�TŌu�U7�g���HT�sc�h��%=B�e�%X����@�0;��̦���()L�HE����j�@8��b����޼	��a�y8[^��H�*�N�-P���:엾>.B�T�y����@�D'��Pj���ob)7��g)-D~�N�'ň�u5I�Oo��n����#���9���)� �z	�0�.}�8�1�S�E��K�4�F@ș.��`�Ŀ�d���7E����g���9U�~�	��L+���)3�I���&�`h�Cx�]�%�|;.�aq�њ`�oT��(J�X�5�M�Oi<wd�z3�,#�H�^��J��]�ZpoVv���	�~=���������Eɂ8�Ь6����I���	Yt�y��(��L��L�9�ό��#]�$#���&ǌ^���C%oc�e8��{�n�j�������D+\�3��@�܀5��:�P�8�Ҏ���g�����Q6 8̠(4����V:�����k�_}�c��=DzZ�裧���|�)_���
Đ��?�ɸ��e��{��e�py�ܰr�@��24��pn�$,6���9�АQVd��D�n��q}:�@�f�y���8��`�<F�d��6L!�iG��1p>S��Ht���$�_�
V��6d����B)I`C�YZ1@:1g�]3$3�������k���	8�7F�B���P�an�Z�8jE-�,�ZgR�]�!��J2*g��&j���?��gN�%�$p]p��=-�����s� �6u[V�,g��u�L�|]^�r&��i)N
�,�?g�X#qUyW����ǅ<�?��ݾ��)���G�q���}@�e��(��my�C���Xi��&}LQ�=0{WbI�1x����Ӊ�O���)��^�=e1�^�j|K���X�Gk5���8˘�gD{�&�4[˰��B͵���DO�#�����Q�ecB�@t-߀C�\�.z�k�;+2]�Z^�s�&���#e���B�W�ćx��<�<� ێ�^\�҉���6�z��)8SB�Z�n#�Vx������H�9A�j�����-�w�6�!*�(�I���r�K*��̟�����:8J%�r�Ǉ�J� ����?������V�����m=X�R�Ցzݸo���}ӥ=͵3�1��"B
_f�	d?��������_���d�����-F�W�H��w�H�,c!C�Tc��ھ�:q;y��拷���݉�tY宴�A�DgG����
����ڸ!�j�cq��eF�v�,
NEW��vE�tm�-��ȼI���-ebEߩŗSʿ�CAH�T���oy�T�?��iǝF�׎%�����ജ|A��&G��o9��y�O4j?�!7����7�G����S"��p ,T����jZ4ג&d[�xa���S�/�SY�wW����S�`e���=��!3ʙy�Y���b��ڿq�"�@=���+�c�ȸ&-p9��GGܛc~^�.	��]\�rQ9�ތ��j?ў�x�!$}�ԭ�o�s6[���L,��F2��<�>� +p�6=WJR�ޘ}��cx�Ϲ�N�ۃ��q�o�"�t�k�L�4ӟ�a��%\�x�M)��"�W�������I��{4�t�{D�!kB��-����ȣܒ�U*�_qIF;��OL,K�P8��Թ�d�di�+֝�D���S�� �S_{w�p,&�|��Ig.Nʐ_������e'����N?���nt)Ǥ����,Jt��TiJЫ�A���t�茦�5�ກ��F�"Ų:ɰ-��>��8|q8�j�ú�d�Bn�qv�}E8��!�V)�i��K��Bf�W�
A����p ��ODާ����귬�v�V�:��h^�ϊ�Ï��� �Ľq�(��6�C��j�;��g"]~q�Bi"ԓ~��]�4��(`��gd��P{���(.����]�v"�'����-��o�a�N��΢��1�ռ⥸ /����N���w~J��1�^ȏ����R��CL��?���x�vU��|0��ɗ�Y�Sq&��c�6���ݑn�~�df��U�U/���D�i� �j��ă�
k�Ҳua�(t�f��l9$��L�ȕ��ۻ�<�3�%��E���cV��09��Q�Y*P��p��M�$�Xf7T_����Q�t?��[a0�͍�U��
�\i��ڨ�:%}���2I��-!]��4d���t�9�9�7^'~9����7kQ~��u�'�	��6�e�v�p@črw�s �%#{�[s����;<Ϋ��@𓳶[�ޢ�cHC���Ty�E�w���I]�k�U�7B
z�7"�}��8(נU�zz�'��s,;,9L�\#_��	$�~�Y4��lqrW���ܘa���g@K6�x�@�+�/m<H��q;j�Q���h�K��8k�]���2ߝ�}8��h���@��#X�R�*�U�4�b,�ch�tX��b8^;�M>��3�gPl��ن��m�봹���Q�:G���U� ��C:Ys!X�@�ذzǬXy���!D��>٨�|Ȓ�eA\K�g���G����W�d�|A毹�H���0�U	��a��bv�U�ܻ��y�B1��킣�SB@����Y}\�hQwh���2�J��U?��U��%�vN��j�b!�8қ^c;�����\ߥ���5�'}�`5@q ��QҖ�'�<���fX+sD�Ye����?�	a rq$l�q(�
H��y�H�T��qE\����3��[j�	m:�>K\��}E�\W�rDЫ�+c��΀��YpϿx�c�T�����@^��hlӊ�lJ��:Y���F�t �)�ł��gR�#�7�!*�*L9ٴ.\+�h�7�`<����{��~�����+��_��/��s��ەn%�-i�B�Ð�kp7t(��l�{�� u��D�djR�!�Ϗy|#��S|���N��V�S8P<!�ȱ^��0�����ȁ���K�ߑ�'(�DA��3�5�Q6#�Ϛ�����H��Q��10=������n:�u��Z�����~ob��p��}��P��Ks��� ˽ɼ?1m�1 ���Z3b
(1��NF:V�!P���Q���"���l&���nk�n��N��@.�(��~Yс�����'{�����Oޥ92���S����BY97�#aY�p,��kE�	���1��ϧ"�@���Y�2C������KѠD��3��:(tK��F��^2dk2�Ά���#'�^L��]�t�g�P�-���6!
F�8�C��V�W%�'�p1u,���͘���y�cݸ��}�y�,1����E�0p���.���k|k�7`=��B�ƫo��p�w�
v�s93��:8us���]��WL�?d\��ȿ��|����1�p@5�(�g �b�:�?������� �D�O5���,+m�\���P����	 p�A|� ��������1k�>wg��?��ku�U�$�C[0}�vp��%A�ɍ��_�ȣ�����\<�!�((-������ONU��pD侣H�x9cJ���#��o#�8"���������5DӶ�$��,Ī/�=����N��5N��j.��ꔋ'����2���� �Y��R��̼���"7�h82퐘��P_����Ne���1R~*�7��ۉQ�- X��w��	�����qtP��K^��C�C�,���JЄ���?YnH�4F��z>����+(����`�_n�.]�+�a�Ʌ�>�	���Q�5��֛T������V Vf���E���p��2-"&�l�HZ`�ϛ��@_���!�����<�p;�w�������`��o+��P��F�ٞm�?z��s���N���zR?+=B�ls�O��׫k�T����vi�m�L���@��at�=�.yf��T�
�� ��Qv����~W���Hpo->�M���U$�c�{<;C�Ͻ�^vC��|D�/�dC�k��,�j{M�D���#�I��޷�R]%L<;�Ez�Mhݦ��8d��=�?��x��ڰ�V�{%�y<�(���=�緦*O�tT��P����*/�= M�N���.!9�o@�����p��M6��=;�Ji��6�?��2�^-n'ΩV��ֽ%�3FO1�G|�S��a(���&x����b��»_%Pl��$��ϯ��J �"��O������w���Ma�i�"_��i�75�{������N��=x�QI:����������)�	[u�>����]�Fd��D��KOX�Q�/�r�!��W�WӾdM1�h�`<1ɔ�뗣���@G�z3�<��w�P�ن/�ߠglAo��&^qL7F��A5� �MC�r� ��M��XA�c�(��C��5�������W~����VL\�cRc��"��3���&<N ���^D���X�E)B�S�џ�����WirqF��[����>�2��L����v��ix�4P|OZ򏿍��8�:[�Inд��:��'P
_�����=�.���r�y�*�UI�������d]�w������1U��r6�����ԋA��)���u�W#֫~�����E��ax@����I���@��v�DI���� |1ku�X�C�}�F��x�</=B,~��U]uJA�'I��!Er-<0�q}��:��n�}] ��w����G:�
�N��zN�t#61Ԝ��&�8)��'��ܙ��G,���8g�,I-��4�(�x:�vRF�.���㎕?P
}�_E�XȁKF�y"랚�ej;��pJ#��Kk��s(V���������"��50�J�I����C���o����'�: ��)x�`�����/44<A(�����h���1wɞ�G����b�}j��#��֎��OB���:pb��zB��K�1���o^BL��H�l`?��(��Q��-���L���"����\�.�c�>�*�&;���_���u{�j��zD�����2��(s��:3t�A~Tm�
;����������n4}K��i&��"��2�0���Z�!�h��Au,��ND�ʫ��/�J"2�e�V�"��ͮ�r?܀Qk|�2WnTn|�.��S%�r�c���:�=�&"�h�b�k:�4����sm�M_4�⽽s���N� �l7V�F�����)
	�&;�:	U_Qk&+�>�<j�����7҄�|n�j�{�ݴ�^ð	y���W'xW���yˍx�K����� �U�����1�c���]���S>)�/�?
m�9���e/�^��p#�j�Vw*H��&��\= ��eg�ܯN8����7v1�F(�����,v�t�|�G����%�6��#Á���Lh��$`����~F�WJcc�u=��w�)� �I�}PJF��
.4����ӿ��֬�X�n�8��p;f���ܮf1��!dt,C��c�ܼ�l�g�6��m2;�������oՠN�����{� ١�CE�RF<ؙu�q�5�؝z�_8:�m��:��>��*�F��v�E'��4Mo��"�Q>��Xj��eX��U�'G�(O<|B�� ]�H��#;��Yո�Q��q _�b
���L���ϟ��O{�!@�V-��S9���=eB�qv���v�û\��4-[˿�Z�C��~N����M�_v��3���^�)zZzD�R����U��A�ʇ�E���Z����8<����1��M�*��.
�ojT��I���ɂ%�Y=
U�L*����?��B�M�x���Xq�B��ϩ����G�촻��U⤏����&���OZb1N���!�D�[����|;���L7#C6��`�Jؕ��W;�vT���!۹����0�?��@�jT��v�#Jjږ���w6�>n����4�w�xdX����7�-g�T��2����]���3�`xe�d�"����j����%�/ ii{��#�g�=�Je}��3�(s�f_1_ק`�ޛ�f��+�D6�Щ{#c�[H�ȪP�7o����^�`F����,m�c�9�)��7ջ�����A�U5v���d�r{����w$q�m_�QM_C�9�3�0����*��D- �K�H��h�ዋG�R(�N�6j���b��,f,ڡmVy��`(��r��S�~y�A�J���),�\8�|^:Qa�TV�����T	 �2��V���G1�p�&���W�þH ?���38#�	�K�:� ��)P��f��o�����|��&J����I��Ll�jr��Ti�Ќjé��^LVM�{�qC��lg�����T�A�N4�:.gw�����@�Ga˧���L&����屰�9s3'�A��::�]�s`�d\T��zS�8�˱�A�)Nu~p����.�8�)�~�:����k_�������*��w��?5����#U�̆Ca3R[� ��?8����.��o��1(R�銲[�LɾkldSY��K�e�5�*nU���:�%iP����*C�����z
���tw(��7a%��HE��L���R�\9�B�sL����J<�܇�fo�7NӖ��Ģ[�)�(��52D���w!Q$8�w� 6texL��|2�{�޺�Ct�k���03#�sC�HiBg��ݥ��(�RR��de����zyg�fQB�̑:[u�6�F�ݜ���L>$�-R���;ζ���xU��~Qߜ���Mj31���J��{'-_��aY {&@~�e!l�$�<@פ
�Amj��]=Fgd��$zDn�^���l�~�ɽ�^&`��ƚ7B��N����b���K.�~-�0J�e����䒒��6�l�����g��u���6�@�Er2 mu#h��S��G�Ew]"��9c�gmÐ��ջ�J���{|���aD����d�1����F�h�':�G�R�&�ϓBvm������i�s�A������O�g�����92�labw�x]!�TwF���D��>����66
��TTB>~��p��I�q��ߐ�+&��H��U>9˕�xaZ5j���QZ��Kp��S�l(�����GR�n��	�Ht{�s��.�L�ºݎ������
�]~G��7�5T!�C����
��y*����G��M]Xt��Y�jP6���4��	k/�O����M'ޔ*�؛�Ȓ��y�1�Vف���&��u�zPS3���k9�j�e�xY,��̔<^���jn>�,jYr\^�"�i��o�Ϋ���=�����]�~+CT�!Mm�jz-{7p��s�@D���W!y���ـ�10T����*��N<v�����:]Ӕ�\��6a~�K������	S6���Џ����q���-�;��KpL�l�C�6WWT��r�h����������zh����@c�YmuSz�V5Bg�Xx�U�)jxE�f�����㠨U��2�jۋ��P����H����up��}�!��d�W�D�A;�}��N�GW��O`�⸲��ȳz�(;�M�X��A{#k�����C����mB1���@r�� ��Կμ��8�Y12���ln�b�2=,}�q4��I9H_�^LB��G�����Qݤ�<k*b8Q�bԲG��v��tV�A�m�~;�?�b�<�ʡ9��S�qs8�¸�'z�V���}N:{�ܓ��W~�[�q�(�v֬�@%#�����`N�ŕ$D32�������7x3��t���
�-N��o2N���C���Bw��c
ڨ�mApGnd}O�
3�=�D���o+~Y��!��e-��T{�&eX�a~��"@�(X���`�7�E�fu�v�i"�������<�C���.�����+6������Zpxm������?_�`���R��10�L��>.��=�S8G?�Һ��79w�T7ڽd��	�ϸL�L�1c/C$������,+(�*��p� �:b�g�ȵw��R�4a�Q����[L4�o6D��c���VI�@,e�1�W/�����xA�i��Ĥc*2׳6-��(&�r��3	�@2�%wg�Q��9ۄ���۩[uw� ����8p��{��I�JS���K�ǜ~�|������g��U
�e]�T몐1|�D�v��o���)@�i��w�:E��8���I)av9~���0�$ø���C�:5F�2h����F�m��ye��¢ �E��˛=/�� !)�i�~"��,�O��ΰ�fX�Y�?n���aj�J5EP,�<5բ���5���ͷ��U�-�W#"f��f�vq�N�}uLY�W;p�VM~����~�k�MR�{�>tj$`�'Tb(o�9�J�(T$�s���ږ�Ȓ$�Z���)뽕75�\�Ps6���h�˵�f����ʾ�k�|�]�q9ܖ:4"�Es��h�2�#�J���s��Y�T�ܨ��b�+A t �P�Gc	z1�ڬ�� {�+$P���X�����$����y����
����N}k��'-�>��},�r6�.�K������$]͒��)J�Mn��B�ũ(C���̯s)X2!l���aGsN0��]f�LcȞ���Tn��0\pWt���}!,�"!4�qX��ƞ���uӁ�)HM��h?ٛj!b��|�
��B����˫�8=�|=�i���X=�9�Z�ע�l�]�@ �8$�&������8��g��[������;V?��5�>����E,8�Oޙ\/�ɰ�Vq�l�Yb ��sҜ�;����*.�K[�̠�@�@%}�a� �{`c�����'gq	����k�	��\?�X�g��J��+�d5�|ʳ���I�4 �\z� +0U��`(���_v��-�uI!�T��$�Z]y����,��%��E���\Ԓ{�,J�ų4����D1��
���5	HоF�meS�0N��l��UŊEVǁ�Qײ�,r2�z�.�H�B�lƇL8�����^%kna�^�WS�N7�1��b�`�s�"�*�¢�)t�Y� �S���O@Qչǰ#���ơY)oJ7J�h�N��l\y4�������cq$|�yf�YlW�ƫ�&Õα�<xyY������[X��_1ζ	΁T��Lo�փm���RV�x	���5"͠�V��b��v����Lw.PX+�_��i�0���N�:��&�"q�`����\c�ey*���`B@z�f�^ �0 4&q�:���h��zMC�N��ݴ9�'Z��2��*Ne����/�&�v}A:ײ��0��{�8sC�YI�lˣ=�'�\W�n��}G�B��(��\$��E%"�on�f����v}T~��H�yO.����Ԙ��iUR��뫆��T\�U�x�^���1eE3���mP�zPeK�qHvK{rι������{��e��h!$��4I'�Y?�C�R,����n셮{8u��i�`r��� ���΢�6h1��d�,$M�0Q*���e�����C�w�M�9w�]���0�@�� �����!�o�7���Fⱃ
dݯ��b�`�b�1���A�0>�����b#��c����h�Ш��0��=��reޫ�:���4g4]"��$��Dg���xՔr-�������שО:o �4;H��k^Io	�.��1�k���F�q���tt�Pfb�`�N]����Ɇf�]��a��l�hZ� �/���K9�ϸ���y�a���*���3��%� ��=�F�QfѨ۸�X�{��$��3��t� ��:^�������P7�X��<�����e�n�q��2���"Y�,w��B�]�QJ�:*�M.��(�)#!}�Cf�b�[ou堺7��q�L�W���4ZN������m�Sq�*5k�b$v��Sq=4��Aw.s�|x#2�z��_��� �t���СZ:9]e��RS���(i8�N��^�i��K�ĶD�^�~��h��)Z$#?���T�3V29@��=2�%>C����}���&��zX߿I�M���ZV^����b�0�ɾ����A�	�ٙGr��*B��~Y��u��^fz>��+�T�0��.y�aU�7d����e �P��N��8�ń�*�a[ Ժ��{�+B��^�r��
B0[0�˖q@b�� 5��0g�`Σ(_߹F�	����,�~L�
mE�g>(���x?��H�K��>���rO��3�l��{��Y]���g�g}4��=����p3��Z#c�Y�L���1xG�#�y��6 � ���|��t,���ke��4�I����s��.�|��MխQ}��t|��������0�fW�E:�h���@��E��Q$y8]|p�BV��FZwb��
󱝟E|��g�u��"����/�~�-e*��@����"(٨A@bd���k��H(b{cu�!�5�|���_�OwRX��`���u�cf�d��2��"�~Q�
.��sU���O/�
w.>x��~�JtS���/0�S�j+��N*W �－VV����?�<��<j�^Qc1��}�R&eS�(�Hu��糋�i�ѸW���:ƿ�r⁜+-6��<���d$�\@���ߝ0��"����ڡ�{/[�Z�ӽ�U��c��u��`�+��"�nx�6׻�����zri,\SDp����k�I�S��X��� ���;��՗�~�z�шE��7[��-����0�nSv�4�N2����ժ]#���}���m������_�7)eH��X��J�,>ɬ�k�%�o0�ĝ��6F��2 �S�>PB��;jP%�$/J�^�"��UJ�Q��W��<�>�Y����@T�w��;�.%�����r�����M?\û��C�sզ�׺��a`ϵ�*����U�egL���'>�Gӎ�:zr)_�#qq��� �\O9ݹ(��q�>���Y�T�q�lcJ�Dt���Z�W#+��
��)��hEe�U�1�YF?�˯�����#gt�T2*��$r��{��d���9Z�%���@d�uq^��sWL�fS��!M�pk �cD�Tݖj�����KԴ�;���tc2�'�M��W�4�]���ˏ
�Ϣ��D��܉_2�1�8~�*�z��W򻁠P��%`�\Ⱥ�S��{L�m����!��!��V����6����?<-�YE蟟~ ?���:�v\�Nn����ƹ�%�R<v�_�.�)RVu�9{=R���FB3n	�c ;�w�>.�n�F�v�pt�U�g�˿��!^����#���|��B�e&���up���h��V������,w����D�Tcir��>M��ď� ���9��I���OX��F߀��t`�Ba��tN�5@�m�榱ڞƉ��1*��?��A���9�H�ӛ�XE,���lˠ,�����vG.s ���)J����#�T�eiZ@�,��H(B������/N�����҃@��w�P}��k"61�V���H㛉�p���R0��piaL��ĉ%��)�����~�_]�Uy��i�X�.>y_;����B�(x��J Z�)�\�tو9���i�%��Y:�_��$b[i�&�	��}��R�G��5��s�t�.�4��7!�̤+�=-1�I����}I�B���eȯ�0ǭaM�Mta��(CDs�\Puf'3F��
��$5��D�;�8�y�0��4c]s�; q��k�4D�
P��0}�$��_f︮���oE�Q�D��7*�o������V��*����5��|Ψ�tpo�{�fA�"QH���?'�^og���4���ߍ�o�%�[EK�7����޲Ytz~��~_��P�y�&t앿�����tLBَS��➖��U�@��7$�$�"Y»��V� �U�Q.�2`8�|%�R�O$dDK���H�m��'1-0t��"�����QH��k�Z�{�a��3�u�/�8�HϚY�(bz�/@����ژ��Y)ׯ��@`mg����Q�<2��j�M�&��O�>�" P��y,s�4�����c��q&0�"�0%�:�R�O��"6( �[��a儜�M�N+���>~5a����
�a����������n�����q�nŧ���n1�е���2sn+��F��\���2���w�E��`�b�ʜj��f�*=87�F�]������UUf�՗�"���魴��y��x.�I$���i�#��v���4�c����h�8/Yh]�%l;f�ܹ�t�� 4:���Kg%ŏX(�I�"�bE:Н���-������ƛgp�X؋R�$�3�
��s�[�r��D�?&$D����svH��"�#(�x��F�!I�
Fd<�LF�sp-���s��ic��u����:�٨R��?��Ws����悻��Y۰P��ll�����������U�r�:<WsǞԞ�_.d~��qc��S�s#��^�*A��6@����"�,)�G�ב�D��^<G���S��a�h���l�å�aO� �B����Oa��O�v]J�¯>�	{����<5�x#�j�0p��]o��U�"׾����]�Ҏ�S��4^�Y��x�j<��B	l2ӽ�h����x�|�����ʘ���U�G����Ky�F��I-����oac�k���`�;!�R䍄x��B��p������6#�q@���<	�N�ʯ�����/�&y����d��V�y�y���yJ�'�q�����Ɏ�s��vǀs	+�F���"� �=������+�,D��Cx��]ֈ��5rZ�{ ^̶�j�S?��(���}���jM�JN�oizR��<D�G���񮠩����JI3�%���t����
D�u/_�ts��<bc
��罶i�4:z	V���{��;��M}'=L��e1�������C�	�a���سl֬�"&MO�Q8Uz(	#�	.����,�M��*�#y��X���Q�-3} Y�?bS������G/�$�]��p�Ս��n��x��*8J���,�����u��wL�����2�u2_����O�ї�TLIz�z�_\�9�~OK�r��	sK�l{� \��<I��0��|M�N����z���~��J�7�G~p��=��;��͓����Jf�~�ǥ�ͤ]�l{F<���Wį?��4��ƭ%E���6��mm=k�￼�����v@�)w �#�C�������v�������:ւ�����˖��t:B���u4n� ��FA��*pQ����}�7G��h ��� ��� ���p�4S�*jv�����Ί]����ge��I~Y�Lɒ:A��jAK��5���Z��#Z�~ z~�Q��Tȑu y7�)�\#�F2���5���|���"��{9�J����y*@2櫧�v�3�t:K���<i$�1�>l	��JcO5K��:V�o�U"]�������Cp�4 �Ep* ����c͗�!Ka�x�|�.��&���<?���2���J��7��jV.qE'����s9v�J�Q���V�c�K�r�&��2�me�!1<)��gb�3�� �8��|{Ӂ�{ ��2A�:-����a��5�q`88m'~����i޳��HȲ�4GU��;�_�1a��z��B��p-�;G�P[�P�������\)�'�.��I�S2�/����.�̲�K��a��x"�L"S�~t�׈>�i��H�גUN�>?O%�䥜#�li~ߦ7�[1BA�0�.0��y"YvY��Dv'����i@���Ú8ܧ�%���C��(��#��vD�޼��N _�bM�c�148�r���n�?�*��dH�U���: ��W��D��:�3��b��\G��d�=^�3d���a�o.pJ���<����a�q��b�a_�h!/���Gr;����>/ݠ3v�
�����o1�u%O\�d�� %"���O2�7ŝ-�%)��>q��$,�[0�h�?W�l�wrqF<��ߢ�k�ڦ�ɕ��=A+�����{��޵�Ƙ���k@ZI<����j����Oo���[�$�[ڲ��7c8�;"_3�"�FA���ݔ����N���ٴ�B��!j7�ݧ��G��a�N{���ڿ��� %Ph�e�:a�5y�e��oE۞��~K�-����L�J�j���/��o���q�~���2�W�Ë^�ǁ�ã�ꩨ���j�0���Xh'!�!v��G�QY�����af�Y���k[���+���cs����	�ً�c�q�1�[��@j�ˬѻ��"-�[�?R�͏�H��*tBE�L���Ŷ�.���K���ۢ^���]M/�$� C˨�ޢ����V?ۉv[�Y��O�5����2����n�iJ+�������5�����s��D����b������w�
�ؙ���y�\kZņ�+�uxV��M�Az�F,U˿s��H���f�^��-��/	���#�PfdnT��'�v7�n
~,e)��GA���I9�.ط7w[�h6�����CY� ��o�1,��Y�1��;�%� g{��`8��;B2+2rᆙ}A@�m�bE�]a;���r#�����  �R����]o�BG��Ӈ^N ϓ�s:��4�W��CI�0�	EK�o��8���{���@cE����ƛ�K�uYP`�=CRR�F
\
�oV�󎄶FO�|�����"�|��}/X��vV3�Bo�U��Ma�$M���F{��}C�����N��
2	Y���1���}���y['q�k�n*�r��A�V,3D��e{F^H|�m�r,��ۚ��@8�Ģ��[j��n�G�I?�0���]�V8A��8�{�6�D�R.��oe*���q"1�s�P��vgj<� hr?%���pit9��p���������%���Ƃ�/����ˢ�6�K*�K�"|1?CX�3��d�7�Ճ������=��\Ғ���k�[I���{f����P�N6��BE8�Ǡ-�|5hX\���}�\ɯ73�{O�1��1�J�KI� \ť_��:⢔*���O�皇|��:D^��i���UXA/�n2Ή�Ml<v�vq����]��?�[d��4~
�*�C �K!�Q�I�Q�����Ɉ^'a1����- ��T�lƫ��0� .��0�:.$�2��k�$�e����8�+��bݗ�9b��lQ�o�VՉ]zQMK����\֝GgP$����p����cփ|pIۺ'�'7Nt̙�UJo90�7#']t�ǐ�*���ydtX9�v�ױ�db���/t���6��y�T��lT�"4>�^J������R��X���-nhPZ4堵�wz��� ]CQ���?��@���P��<���)��������-��-�����fs�\�*��p5ϫRj���hh��J4�ld	�!��ǉ��&�O= �^ȇ�,<�w���۫�P7X�Ӝ��W�P�_G���sm�?�4����,�[t�Y�Lq�>��5v���/"����iٳS�3]����n�}~�$/�m����|��

׎)L��G���/���� q(eX�n�����݅4� _�wq),{���TU�o�+��`�i�h��>��2��7xdu�w��e�1e(7�(d/���@�����Zz�#��wn�A\�sM!#��!�mD���.�h��Ɵ���q��^��q��U�0W!y#�j��Z����S�y�f�7����Ҡ��GM��*�~8X!/���s�{��x�d�>���0�X@����1��8J�l���F�(J8�[4{6A+A�c^��P�q5��zE���c;M�(�z�2C���hގ<I����Z<���6����OT0�c���=�miNL�Z$�r�6I,F5���G"�b�3�|T�z�p����4�2�ZL��Dd�ҋ����лr��~K��c��~$��M�����#7�#m ��ټ��'%�R�\8�j@�MQFmd��l�X��-4�����uym����_�n�e��t�|���>�Z���;��}�
ئY~+�ʣ1j�i��
@�̉8�)��A�B���ip&�i�R���B;�Kl��4�K|�����_��<D\����lAwQ9��7*0k������Kw	}��ܱy��'�T2�:�k"��($�:�i ���DX�з
�Q>�a��tԽ��
��b(�LK�!�����i W��� �mx�q���}P�ۜ�d�ݸy9}�Lzk��mo��O9�����B���	���e���x3��!�!Ώ��|���mc
\����N�2<�$>������ۻ�``��S�]�ۂ�Ⱦ0C}�v�6��:{�'9�m�@�6lmO|>B��_��i<��n�]�'�B��E�|�*�����QM�D'�3q5�~���5�Ҹ l