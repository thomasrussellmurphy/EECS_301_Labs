��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\���V�fnvx��ÍG_;�ȅe�~�>���9�>��Y;�0G.䭈N:�*�>^��V>�6XVuYM�Yy���=�a�FY�����,��i�ܵa�z �k��ϊG��-"�.\�CIr���q��y-�JJw���Tdz!�߇���MY��^����E:��R����{7K����P)S�$-����sA��*`�.Xs�?��n�t��-(�u�X\����'�0�ެ�������#��Jk����ӹ����C,��%�2��ڥD���u�$�{��՘��b�bd �RN���5z_.D/Q"9�k=gB_���`l1�心��3zx-��'��~$w$�T� �ɇ�Ho������m�Ȳ��S��}�<4�JC��,��f)%��fT� �Cx�<+��Wc�/i'_��Ș�E1�mA����4�2�^��N�B_�ɐs�B�Q
J���l���0�GD�����,�]]V�UmH�#���yg��*�%�9�4Ud�y���}�%O��&���L�A)��̞�lڿ<t��[}� �Ņb���'��U�_k��4g��t&�g�)�������Vm����>:l��|����C{-�7�&ek��s���餁b\�pŀ��>�Jj�ϐX0�4�3���ʒc\��$�Js��	_��GY�\f6j(��^<��nC�%����\ �r�刵����{����7�����k�̭�����v9�K͏�1�+�=�V�	�m��I:�s
��ɶ>6eA��>]�P��lMB� te�e�I���ш����\ETV��d�)3��T�丧����<ȧU��:j�ڢ(��f�F��lbV2N�`�+�iD���^�i9lT:|�u��t���:�W�]x7��P�q��e���v&��mpFG�Ɔ�&-����"�=�xŒs!�-�	�۪BEl������
���z�ݧi�/wf2Q�~Kb�z�ˆp�k:��o���Լ��%rҐ����az�8���6$h�sn/X9�6��E�@i�~R	��U��@��)D]�g���G���Ts�`��:�쌿������Яgs�����Ka��?t������i���'"2}mq�C��ԊY /ͭ���![򪌹���/3��P�ֈ�q�Z3�i%d��GW\*L"�'"�
�(�_A\[fG��#Q᠂��^��n-'�u�Kg��~�q���g8�5Y��5��]�ߧ��E0�yo�Ȫ��,�kV���?����W�4��������n�p�_�=s�&�"QP7vY:ދ�����a+2x�͞��*v�ouo/��C�H�l�ۑ�f�G� \�S�cwX�5���
�	Kha{�L=C�ͳ?P�c2����� #!
�~i@��"A����\@P�|~�0����7Qs�bfȗG� b`�t�U"��]��ZT5����T��egL_qY���yP���j-�t�с�'�!���ةs��`��Ƕ���;�ћ3v�6�<��ʵ�R�v�����n�d ��Bk��$���IxP�8Vn�d˂�wD9�~I��r#j�jS;��4yA`M�"`�w�>Z��1��@��q��4�2�=�z�;��41>&b9������di���VKP��s�Xz7dD1`���bjJ��'�K�h�g���Y*��jn�b�0hPyw��+sUg����x��zC{��O���h�K�L��T@��)���re)�)%�voٞ� 8�~�����#��%p���ӱ���;�/�L��w���V�Ʈ���m[���8�ys՞TL�!,�Ox �����C��Jrs�$Q�w��g˛nV:�&r���89�F ���0�\7&����,�;�����T2͑ �z/J �*:�!!7:����pC���u�n-4}nnw[r�sJ���.�0��[������^��VV���u}a�����%/O�|QŊ^��KY3m���ŞQ��+IrV�O���r���T�F�}ݭr{ͳ&?��?�W�%T���c�}ȭ��p��1�d�JM!�7�ݮ��|�d������c�}����^�s�U�_5��:�}re��E ���g�h�N^gً9g_�r��q��� P ��z��q�(���C�%�����6&p6�L^sC����!�ٞ��p<@�<*�{�)2Ә�M3�%�iu��864�I�c���S	{���eyOp�?`��8�kd#Ǹ���5�u\�;��@���la^��si�l��?*F�ɐ`��(��b	b'~���iF8c�~	�ҳ��I���b��~��Iu�1��c�xN����+�qׄ4t�tG-��-#0 �8h�k�-�㮉vޓ��
yo����3�aLr&����4} �ɱy	~�~��:+Ȗ�~=�~��^��(��x5�naU�����*�6��gȜ=�H��8�f��en�4�03uefݸ��|z������I	+��	jb��D6'��`�[A�^a� Sd�/롢�9�@�f}��ܔ�c$h+�&�
V8\}9�27	��ǃ��4J�q���<�z�8����^N�~k����N�����=�!d�n<lC�q:g<}{��>C�/:�//��ji'#.䧸����Qޙ��a#��[N��f����d�����i����x��Ơ���ٜ>�����-���*�gq`�"�
��}�ӫ��sO��i3���zz��=��jc�/��z��5�h�;������?/��2��C�}�>�J�a�=�qw���jM���=P]��%�Κ�m"_{��
.;���v�;]��Sx�&^`B�Е�_��*"�<d*�����$��M�H*���$�Ba��s-��pL�Ҋ�߁�4[��J}��'k4�2�߸��?�jȅ{��wU��AÛg�,�&�1�Q5}j�@��!�g1��s����E�	i�-�L����p�d�����`�b�˂p|Q:����X�2�_�@��b�P^�^�"�P�]���_)��YM�r�x<:��P+˽awa�8=V���c����h��01�X�a8Ы3*�o[����5�Cïa��Q6��Q��`h_�)(S�2��w����ti�����i�S��'�"������&@qJ��4&�+XJ�Di��L�1�y�����OG���ܩ��0�10.�	�A��v�\��ev��*��4�P�(?�s��#�Bj�F��if7���~Sp$ZǾ�-��-+�.��5�u6�}������\�S�U��0; 6�I쥘�5f~��6EkV�e��m��󏯥8�R�$Pi<�O��ؖ�j�T|_P�KX-�&�
nE���Ԗ�@a�������	�kHߎu=����@7�.o�Q8����O���8�=`)ٖ��Z+L�n׆
ű� �B}!W@�6q����`;ţfC(p	��3C��x��D�cB[�#"� �I�md#?9��H��m�t�V{7Z�Xw�ș��iC[_�I�lߔ3�I�?��Lc�E����蛒��Cp֗M|��X�v����L6m����8�U(�x�He[h0|0��[FA]�mZ/��?}�I��<$m��!�
*$�P�A�%�
���H���ڜ�7
nh���n:�/�cY�MFE
鏢FVx����M�ޗ:��	6�8�CM��RZ�[½��7�4j&ٱ6�'��b��2t%;�I��.� L��E<�9?��GKy(�+���{*�����xIǙ�:k0v#y֛���i���Y��R��Tv!�h���:!T'�����F���%��ev$�^��-��ջ�5���mN����d�o���}O���т�bŏH�ơ��w�B�钜�<�%��Ƃ5�L��]�F*��4����g0��Mxd;m(�2ݨ
| �RoR2���;�͓�A��M�<U/m�!Z�X8�⛔C������_���I�� P�o�D@6�����5S�`g_��3_b����ɈV1���	(=����̓2̷s��+~;�*�}��J���*H���#Nt�9�Zʇ�n|j��
� Ҵ��@B�#{�V�^<h �E-����S���V.�+�,�������� �,��s�6�Lek+7N��>�C���BIZ��N�{9�Ǵ_O���b~/�l��	h,,*�_M����?\�}��&L�Q-���o-x�Y7�#B��-���C��bUVQ!J?g�}��!�:҈_~Rq[�8]��e0.��}�(�o׶���`�˭ t2�I6��F4|X*�ׅ6u�\�[��E2��p�P�~�&2�Q0�4a�r�A� ?(%����|����{����!1��[��@�Qjb���~�
=��.,?pE������
RG��ζ-�L�ƨl���)Y�(���h��a?1��R�����31n������|�n��X��?j�Y������s*��hU�������K^��ڪ�Z�$p��ܸAl�L����1��ྮ`�<��4}9DL֡�K��~�و��L���9�`�pǘIe��ԅhd����m2������OC�_��;!|�oN�����3�Zj6�fN{�(&�*��4=z4
��&H|����}A�_�}W���bJ�(()��K��t.d���?'K�����������Z��L�?c���(�(B'��_��r6#�:��G�o��J㲦>�Ό�Ts;��9z5��`�̵F!�� A� ��p�!#�	(&~�O�n�5��R�L�pT>y}@D��k`�����_OjJN]<c��[��E����9:<�Mŉ|v����$P<
���y��>�\0���rUO(l��6�QsZ*�a�O��R����R�x$̙�1��;[Ix39K���n [Փ�Ҁ�T� ���=F�B�h���l��Cv�:#�7���|����T�<9l���СX��$�lR�!ృ(x-�_v��,�����݌c�&
�Cf��!!��y�hY~V���'�oɀTHC�4TkY�EՐ�#�w,Nr,�Y�:p��C�T/��}D�ɺ]�MXeĽo�rhM�.?�5M B��B�inD��9�*�>=F�怒�<>�� m��7����Jj��=�I�7�-��
w'�cR��@�͵�r�L�P{w�F`��=֡���:y,?An�t4��w��᳇夷�C><�֊�wN�Q�d.>=�D^ӱٚ���r���Z�8��G�(h�R
?,lu����ȗ���e���q�Mh��H��;��ꄮ
��F ;Șo�0�x}8�Ev�C��'�R���[+���z��1�o� d��4�|,�� �3�^�}���0C'���uJj�歜dr�=G������f*E���g&�E��S�Ȝ�u�/:��;�[����g�^�g�-�'�m�<,�q�Uv��װ���-�Fq�tl��k��?u���I��q���Q�v�Oq)
S�i�_@�Z�H�4'�}���O86�V�Ҕ�)jRUr�@��T5}�� ��x?)8c��o0���?�ٔ0�Q�rG>�x���xOx�a�`R.��Z͉��[��ϰ&ޑr $�,4��T`9�D�w6~��p�-�Y�N/��-���zH���b�Fs_v��A�/Eܬ$Ơ?�ȥ�
p��D�*�H<��i�]>!�&7~�(�is�܋S�(�+�kEUμU��� D#&��p<@q��ٚp����Mv����	�>y��XJ�Sj��m�̳AUg ��j�mw�R�E�ρ 9�K��@���.M��P%���I?|&���ꅎ��9�R�?&j�@s8=�������ڣ��8%d�^����KX�&N�e��x}O'0@�\���R8�=0�5���_p�.M2�� �[����yx��v�������L[k�P�7���E���$���0���xLOo/V�7G���5���ֲ��BWJH[5�-wY7o�6$��N�H?1���X7<�yy�(�1O����(2AH
-��bp靄]c�GJ�M���X�k������yȂ���]8�K�H�f���X1*ጬmhd�F)C�%��=3�'�����0k���._�6�"=$<M��q���1�����ـZ�l�W������Etk��;����O�j$Ԅ�
<����/�=�sXk��(���]�GP���Ԑ?�ݔL!�)$Dx�y� w�w�4��7N`�K]g�	�2DN����2NG���Ƞ����[���P��ҏ��`�����	�x�3��ڞ�#�SE4�`�*%Sp�Һ���\\���^/��]� *K�O9�⌍rR�8,�8EH�.~�.v�r�gP��f�{Lnղ!
���q�$N��k҆�L�o�\�l%�y&Ч��a|�A�|�R��U.z���E��ő?K/uA���������⡽��q����`c��W�Jd���.��;�~6�uB��o�̏�d&�$�)v����!�!i�[�sp�t�� zD̦���y�9�f���T7X�v��8?>��%Gp�17ؑ���eC�����1�[�<+{lzz��	q?h�i$Z�|6TZ	����z߷?a�b��m��q����u�r�4�@7V�D�9��d��CN�=��ũS�(mT*������M$ʹ4	\�y�l������\ĩA���5��I����0(VOe����T;l�#�#н
zf�㘧~s|HNahކ�G �<��jrLƔ����Uۉ���\k��Z���ѹ%�<�K�]���9��4	�hk߸��d��17S�-�2�����<M�����P2x^}��0��>.�;X̏���^�*�e�>���,�7�g���,���6Y͐���خ��t����T�
3�]kSЌ�_�H�BG|�K2�[�0�A��(Oaf��~��n�p-�����Ji����g�4�Os�K�F�7�ͅ�Ck�W�b���R%�`�R���}��[U�bk�Ȱ&1L�׽�Y�7+���F-��1W�h�:܍�n�v�q��惉�5Q���L�?iqd��2,G� �S��_W{]vW��qM� а�Cc*oy8�-ӭ��I��G�2���NR�i �sG	c��@�k=y~F�ڎ������#wr�ͤ��3C��c�=�ý�����a�B���&�پ�>�oI@�cصV$��AB1���0�Ү��%D�.�_l��b�2!�LZ��d����)j(�@�Q���~��vUl~"Y�[O ���)��Z�+i�V�s��u��z#	萗ի7
R�+�x��Ф�AA-hÖe+[��QI-� Ԓ�TK��O��A�j�P�b .��/�����+�w�5��<�#��W�I�(��b���:_$�2�x��Gzܥ�~�J	�=pki}��a�ak���ȫ��&���d�Q��3'ۮ_��1��q_l��D�V�0�A2~	����b��
���Q��4z�b��F�9�@�?�� �-e�r�DY�Dw�Q����E�,���	�������\��d@��n㙓ا,asj��o~��UC��w�kٿ�� �j&��v[T��5Z�j ��0LCI�;^����6{�e{�Tt�^į�x6�H�+��L�l]z�s�UAU��8ll���"a��\36=f3���v����h��U�|g��v����\�?|�0�rl�K%t>: ��/'�܆��!����3ӓ�
Y��8��a��x��B*4�U4v�%M�>Ms�nQL?~����A	���-�D	0+��ES�;��2�P���;���#JF_M�MZY�x�m����ǵ�P8H� ħ��ENE�է��Cлv�b����\ۺ�`���c{.�}�]�u��p-��rm�~�m�9�]�ؼq�.��|'�P��FN�*�͋US�6���!j��Dm��.�fa�R��������*�B��]3������5��\N+uJ�O�#0��TW.8�X�ѷ�+x�1��� �Lc�j���p[�����lJ|W$�������!��o�g��H�:�m"`}R�ja�ov�4sѻ}����|��W�H�XN�a�h�R�f>R����3��c�xu�gW���Y�ˢَ�����פ:yٕ�ڑD�z����Ð��tB$h8'�����W	C��|����My�mK���г��FmXe?����a�@�w��1�I�1�������������)����+ў݄�0oV��/<��$ ���3��-����PO��+�����-���>���K�������L�ٵ���'Č>�t�`)0wl���zM�����nuf���1G�8�hZ��b�*5�&SE�Ԙr��A�:��Y�iC�ඒ��-�g���s���ڒK9t-�TT>;VHE����9C*ۧ�B��|���	Z�.Upv$���Z�����s��U�H��J��d������X�(�"���&&�q�Oo���aW�.�"Q@�%:�|#�����Ƣd�8���|��U�Es�R�s9ً]@X�s[|3��񐽠�H����*�o��{|��[���c��zrk� S;������Y�="�G��G�Pp�Ƨ1~��椂�i�v)e��q_�(��/�.�Y)Gp�5_��r>dܵ\�?W|"6���}��н��wQ�m����Ċ �W������w�HE�ɏ��9�1܄�@#�5�ҽZ}�����ϳt�4�u�T%�OwI`*U�П�i��.C��{�@[�!�R�@;-���� I݋�më��@����S�F�Y٫��x�ʟ���
�I�M��W��ʹb����=ъ��lP��9a:	��P�oi�]���%Y�ki���b'���:]/~L��fEa��WXX�� Gªn�"��i���"���U ��'nԈO��ml�ģFd��j�^~����L�Ij�X�&�()O)��U�oyd����&��^^38sLV��R���>���4�u&B��pe�e��4<ʹa�m���|YI��\鵆��%��1��D-���y��</�ȗ2�+��biҋLPb�