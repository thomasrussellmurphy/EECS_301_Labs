��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\���V�fnvx��ÍG_;�ȅe�~�>���9�>��Y;�0GN����SlS��{����W�y'�Z`0lk\Y��j4قg�W���� ��B2�a�,��O(�W��[mmR�� ���:������)4�$,��)�c�����+	�)c��k�L��w�h�xYy�D����nس�΂oyt��z>��"U�� ��}&!�"9.k�Z6��ṍ����|�AT���k�j�G�Y�[]�y~��;�-ˍt��gQ�񿟇�aɤk��^l��;�-t���gE�:�t��TA�?����.���\L�F���Е
��Fh���j��gg�
h*;�ُкs�RΠ�����<d�M@�8�%s�S�i�:h���h�V��V:���4�	�gŏ���XM��}ى�}��m_�V�^Wc��{�!Z��zy8!n��4�C��8
/b~�d�X�Ɩ�P	)�����TVnj��K��|�E��c�f�����x��u��������Ij!C0c���+%=VS�5�bQ?�B_�l��C��}0�0	ה���`O����
p*���W"F!��j�Ud=@]�ǳ��		ԋ	K�%&7k����ǈ����:1Fy�b�%�2��>-�K*�F���"���"d�!�j����ܮaz������犫d.>�b�F��x�6q*޽Αx*�B6�bLzώϴ���oS���I��?A��p%𷆋'�R���5U.�{Y䒈�Rŏ��zd�G�b��l��3=���6�M(�=����W��.���Ut��"���FK��2��<�8!��#�*��LU^���yh[���.k����E�Y���|��(���?��3oD�Wm E�t��GyUU}a�"�	�c�QoY4�����-A���s�G�(Oh��v�����r?Zo8�A�&���yn�n���Tw�Ɍ��*y�m9C�� ��6�3O����z���P��� ������8�_�����)�s	]�G�U�
u�i*x�!�\N�ܣ�>�&��o��a��7Eԉ��i�_�%�`R�k��ɉ=Ԓ�/��\&fT}��d9���eEH2E��V��&ك�����[ÌJQ
�"&�"���� ����`J�xf�[m�%�=R�;V�CE�!n�T�����<h�����Qg�O^��$hc��Y��Q�f��6��Mm�r��t�f�~��q�ȬOhݻ�&��`��1 +G?QI�cwd�qp��?T��2�.��_S�6�
�vͦ�Y�_$���K�e绔��z�J�ld3u+d���y ^J�+K�"�Qw
}���o�=/��P�*�I� f�nN�3|t8���y� �ϴ������aT�f�� H5�g"��S!�����l�N��ִO�,����_nV�������x��ߛ���{ZK;�F�k?v�b_���x�Y7����P_��rM�Nu�r-�pOa����F><�V�J�`:bLE�/o>�����|��گ�BE��n����ֈI@�֩�]�$PkI�,|�~�U����� �V)#����g�H��x�� k4��7�iƚǱ���Q�."��1��lt�1
�Iv��d�YC�,�n�� �䛜L	zP���)&��B���~�LǩJ=5sԁ:f����(w��U�9]�$�PI\�c=b�:���r������D�i�� ����II������|d��s���46x�L#�2މ�����#�^�c1wC�e�����5��I)`>En��X�P�h	�ٷ�I���=hw�]qo8-��O6X�U��*e��+T"��'�c�!T[�ɜ�zg[v�xi�y�(,�<ydx�nKax�(�[��"��/��A.a���iBmP��s��I�H���-R[�r]��77x���n�-����-]��\�HB�����g��rH����\Mk!�4t�c3)^�!O!��O�KB+Ƚc-�|�jv9�z��)n��K�"5Z�z�a��p��n��|)*O	�����'�=��
ƛ�

'���?��
� �z!����P�:כ5]F���k*����i���ׇ��o̲�7��?����ĚG���m�KM��v�`�����M�]t�ql�7�ԅ.`ǲ�|���>��k�dF)�z�һ�,-ؿ�]���}f�L��݊v��)�A40�����0vG��N���,"��֊��ed*҃���z�Du������@Hoc��u��g��Y�E�d$�w�	KX@NU�dEO�@���^�)i��S��,8�Q�)49�z��s�p.|N��@A-8o0�;�r���Z:ͷ�W�嚜ʊ$�K9[Ѐ��#�j����f�jq���u!}CJ�����P����4�p�d�	'}�R�cҒ�Kk���Hi��oqK��K���Z�JLI���]`>��@{�dZE9�� �:T+&Y�jxn�����<�]<���v\���*�^FbK�ǚ�v�\��?.d��j�(�x��&��n���Ww|�����L2�����9�S������:Gh��V7�(�ٴ�Ծ!�-;��.`5�xV ��|�B����)~�< S!�f��]��:�O���lG;0׹�w/���1�� �ϛ��4���)S��_��� ա�X���O�~�:"��;l=����1���=�yA݉�ϲ�d)\���|�s�_��d4����	C�awu��8�Y���6�c.�zY�O��LY"	����4@�f�G~u*�.�%̘�g��x6����5j�I��+������'ԅ�-]�yh��	�@�X���cy�)��^�8��T����0�e<!pܦ`-�>�#��9��18� - P��;_)�y�홸as�8���M�3���G�c�)f���߸��Cxl
������[�\�����iԾuSs��sE�#!�����P�0��Xͦ�N�{�����{��MS|�sz�@:0'�tv�����:���#��d���L�������[z}Q��prHL��v?���҉�uD\CF��r�9���`[�x0/yt���"i}�4��P��qB���0�ڃ��*\���-f�ufv!5&
-��X��hLf/���{�/���Du�߆�3��#/��d`H�6ب.k���TZg������U8�ˠ)�$ro��O�LP���6Nw���ٚnj�і%�UE�iWG��`(�7 _-_����QBIS"�-9�e��'�4�-�2�l�XKc<=�B�ib��o��]L�G���~>Q�=�6�����~�h����Ƨ�I�k���5���������(����Z�k�u��(`�z î~f���J*��a���n"�r��5ل��nQ6uԋGǲ[!ʉ��gu�1��:VMw\ƻR��z���7���ef�w۸�Ơ9�3������b�#�iΫ�X�C�z�H��	BҶ�l��p�K�O�w�BH�hP7pv�l�䵪���:�l�:�Gg}!�6x?!�����(�u��P'|�+9&�B^b�/Q*S[�i1���G�6��N)7����L����p>�pw��oe�4
��Ƚ;i���O�R�<��=On]era�q&�# �B��Hu:�'P//^�g��}�Ѣ �bz4��(��P�S�����7�L*gjſ�[d�u1�P�����C�2���VG6'�w��NX�����\'�L���jL����yR���ĵ�	[���f8��zKS��@0�	^�;L%���<�WZFl2��U�u2�~�O�<A�n���)�?D�?L�SI��H��:X��m�L�r3�7��C�t^����xfr��7�|�BR�I`�� 4������[�ހMڔ��,��v�S���W��"W�){��#���T��"��H=�E��@"25.5����+��'�Y�ΜA�.xe�hb��̵8Z���i9Ag�][c^��v �V�b�8�j�;zYϩ@'�X�S,��z���a�����*�}�g��5P^�e*Մ�Q�A�qm@��Z�pDUx�#.����h������ ��,AL�uИ��g1J��U�"`��d4T��Ko�p֋4rt-T�d'zG��B�a�_��6�R&ҳ��Ӻ[	���t����wC}����
�I2 ��;{��5�_�i������A���T��63���Y��O��X��m��H��m�RC~z鸺�s��?hrbn�#iW��!iqĨh��L&��k��n�CO	P�y� �������iF�W��},��r����/cWo�����p��B�;>�u�C��	
 �սn*T����d��'d���=��}s� ]�g�ʖgM0Cq���r)�����i���,�.�7+Z��z9��|��d��ʴ�,�#B��h
U���D9�a��~=���e���`�o�.I3E�����ΙJv�%}1�i�?��A�}]�������tN��-���tūעKO�K��;ZЭ��]L��·uNLZ�3��&�Z�TB��9��I�����7�e���&�)ywlN϶�Ɛy
���b,��d��o|씘���jy�-��v�b��[�����m�a=G/���CuJ#���T�ɼ�O'C�byE����/pT�Z��a݆�P����1}�*���2<(x|qndA�[��j|���%We��cF�����`e�k�ͲÔ���W@7�y�pr?cxS��Vx��)\�:��L�����Q�uR7T��{�d���~���o�#�H���k�E� B��q�J�νu�c��{�=�18'��aU:@Deb����۠�9��v��sW�Z.��w���L��;���~��TM=1'����Ap^�ǃ�����Wײ��é+;�}>�m���GZ�M~��c<��-�J���%L(�������1.��m�h����T����PiXy\S�"����/~F���y��z����^Q�?�az4xI�U�ߛz���g�Nz��{%Ґ�R��Rrr��J�kDG�����e����p�.�B��郒����/_��\H�y�V��A�wV�
'��^Ύ��\���
�����ם.���v��H��tW2�f��]�F��	�`�[`���� D�]Wo�Py<���lM���ݕ�5H��>0J|�4fI�,j�om��p�^CPD��������e�ѷ��C�޸��E���P
���z|.���S���[�
_���bdO�Ϝ4��0b�g����� X�+�E�f�1IL��1+o�(�/�/6�4ٻ8Ձ)�. �@#�E(��^:~0�n��Q&=���m�e�x˹��.ޏ#|����U�&�kyh�o��5tX����z���͘Z�=�l�q�^I�j�S�_��5g�E]�v3J�p��k�`̀��+z%��Q�f������<�b�
�+o�Z�n^a�$Z�V�~e��La��.�̓�^`��d?̜�8�c/U�s�(����4�c��8%�����X�Ear�9�K0:��ok��B+,a��̦e�WirQ���z	B�bm%����ډ���q*�w�I_#�q&���9*�A����΀�i��<�y����l�����ݵ��v�f�RU�?��cj^��'�߀�̟�@��<k/��XV}���病��{m�T��@D��a}�Ϸ�4׏m�ni�4���J��UI�P�;]F�u����_�1�q�S�D�|�{�j�xC2�5YqŶ��D���ük�o�f���=��>��܊lr�k�B�6���N���@#X�Z��Qۖ'tg���=���T����;����Dk:<��ޘ>�1_P��8��6˄Ϛ����d�������,�JZ6��[Ո��8!��Ŏ�`���~���Ѽ�,�����*zk�����]�af53�CF���L�UĠ>��)�)O<��m�� ��=��_F���@r*W����Ze��S�����Oэ0M0�#L���Fj�wa48��eU�䞟�w9��v���Ě|�+�MgP?�!'���w���U��&��/�(�����r�rSPs/�i�6t��iȧ��*��$��+T7���)��(�7��8׈b�(@��
���t�ܢ��0Q�zB�l���
��o���g�-�ҏW�%���lR���쯑=�Z}�]��f���T$��^rg��1e��^LĻ��Y��N��>N=p۬���Ca�ta{��?=p3�!�!U[��>.�V����%e4p!f�M�v}��E�� /�m�yB���a~2Q�T�H���[�	�Om�ɑ�m/��h-_h���Mf�����H�/�}8��g�A�2�hQ����uwdW�W�)d�~�����-��`�fߕ;�Dc9ւ���jf{�Y0��\s�''�B���Oh'�g{q~�r+�E��2�ųȘa���%2�C��Ub*i����$g�+��꿇�
��ۼ������ݨc���
����_��p��'W�vC7�1�gJ�G���Q�H.s��m�Vʹ3I ��[����UDU�VUFxB\�^{�`k�-�+/Q7��x�^�s�q��iDХ�{�B4�=�i����^硡}{������7ܹ���!��E�hfR����u��T�`"=����|��Zʏ�� !�݆�4b[��2�;�J����gx&�b?�Qr�b\2�(�����*ƔD�/Z���E�8%�����ǧ�'�_P1�FQ�bg�ˆN��ZRN�lKD�R����&N��i��j�`Ū C]W1�Ρ�f,+�c�a�|/�O���(�n8ԯ!&l�k|��Z\5%��PK���A2�C��]�($Q���J;[fIfU��eO��D�N����d�v��2��z�Yq�4诟ӄ������c����]K�����z����\����i6�u������4(�~s��w�{�����<b$g�n���pA���P&� <o�F��=1t�\}@����ks^���I���>nA�y:�~�n�̽����莞F7ͺ��4���lB�n���>�P�1A�)5�i6���i������g���~J�jԦ�Nyޅ�1��C��#X���	�ă]�T�����5�v1������mF3���M�������9��eH_��^ޓ�S���t�>{��_)����M}8]��Z��H�zslp�l��fP�����~V�ُ�	u�n%&����F�˞L���_(~���l�k��@��L�f�������֍X�;���f�gj�!��Q�ގ���'�B0gc���<��P*�_�$$gTu���/��=��Ctu�O&�J��W���t� Ier��`�_(}m��2���u��'E��oΥ^^����2vC������Zyty�XB?�fHn���9�s=�ֶGsq	������4��Bۃ�B�|>ٔ��"�^P���>Ta�T�r�<0O�_�|�uMO��^`�(�r�h�=���'����|J��#�R6[��?E(��D@�f��*��L������Zs����Φδ�?��<�$��~HD�B�3Ų�}@�D&0B�]^�g����dJ�.N�9��f-j~�Q��};�h��\�g��$����Ĕ�y�ra�+n��l6�ҍ?h�!�e
��[��d�[}N�J��7���YP�4��O�r����r�F͒>z���H!��r�0����$J	�M�U�Y��`nXw'������K������-�����%*	�N�Em�Ϸ���n��p���D��4sR}&6�X����Uɚ��5�q@2F��`����H|T�~��E��QK{19�=�)Z�zY׭z؊�w�m�F+"·��5�#6�{^7[i)+����Wh��Ż[�5\'���&P;<rR�����i$���0�L�-���37�=�{�K艁kF�� �v+A�(�Ghi����;��`�\��HXE��K�7�&WM����jRm������꿌�8��o��9K��|~��{����	^2�ሁ�S�]�v�q%+֋��ٛ-h�Zo-|�L����y_�C�F9��j`�xc����/����\�f6o���I�Z8�ޝ e�Zh�׏l�Nd�7®{�򍵷# ��vx�C�$��FlAÝ����R��/�h�7D�N����������N ?��R&$l���@݂͍Jw�R����J��N�N�g�\XM����n@��U5��4
�8�E��Mg�!	\��N�k��O*�1�)%7r���w:%��Y��xw_\۱X���|�Ţ��g#X�-�#�	}\��1:���/yU�W�;����@��t�t -ğq�$Ơ���E�n�0���s�W��a&4�:��OUA��O`��%3�������AHnC���0I�LԾ]�F`ƙ)K0(�]���MB>>PL�N��Hw�m�w���o-OiG�o�=)�d��Sp�+��U���רO5�\��	ͻ.ئ�����,'����q=�����S�u�'مHq��|$��{�LA,�,c�n���L,k��|T>��\+$Ǭ�7C��+ZJV�0��f�3�{�ք�E`#y]�I�d����/Clʕ#�,K���E��a���M 0T����6�1	��1 ���P��;�zA�R��ڧx)��p2����F)�;.K�1�����m*��o�l?"tm�-|�a��n��T$������{���N�/�����E�$�E�4�r=�tA/RL��eQ��J�L4����#�(Ӗ�9�����H\���,���?������x��1/?�՞����������4>�5�A�fnM;��w�T퉡d-Q§�S�@��伟�)���9��-�O3���k-�B����]�1s]Jm��o�ps(�!2���/�5r�B�޿T1̂R �TkH��Ck�"&��ԉ�{.�q%�� Ao��ee攡�ָo`gw�sH���*8꓉��t,S���Jij�{�6HW�lO^��6��U�����+DX)��K'�k��`��W����:a1٧,<?�٧X�oD�n�e�b	;���	h�]���f�>9�ό���^�-=�?7�F�<�N,�<X�,���|A;'�B���A�7f2c�=*��8�c��컥�T�샯g�\�m)Ѯr�Ɔ�R}� uC���_k�V��oVk���1L(�+߅��D5 ���u#�h�3�Ф�>�kR�_q;���(���a\���E�Y��`�5H�gJN��F[\����<M�=\w�"ΤF�Ih��N0o��;e T��h��]��h��R��%7X�I��~������<|�Jv�ϔ��&U�w�ƛ�oj(���S(m����
g��v�����b|�J&Fi����Ґ�Y���v�-�dX#�H�֪ߪԩe��[���T��Y{0*`����R����>��O�L//��N�RR*Ѓ�x���
�٭�P��sr��С!5��PWl�38�<��0��8�ңl)����-�.�M�g?K]+�	���c��2�6��2�gA�i�ꎧY���ߝ�M3L�.�suX��H�� �1J%WG�X��h�m�t�/�9�"G�$��Owt�}	.�Ƹ���,�ܯ�񐕻|��l��F=���{3[4�r���4�K����@��('�[须-��o%�{+L�߼$y&D�~SG�&>Y(&���멵L�pb�#���	=|q$�"Sx�M�.r�uD��2H��ÿ�ZZ��TG�Q��w�ZdS�4��[#{��oֲ�}�E9��/fGnF,��z��^w~�fۭf�&�3�:#ej`Gd3��%���荁�ix�jkF�<�wh4w�H۹�2���n�2��^a�D�˩dr%��o/��A��V��R]�	v	16h6�(�n�]`X��y\�?~�p��@|���K��N)�o��f��e���Q ���i&�t�����]o8�*���&�R��.K�˙{���S�[of�bk[XC���;6I�w�!8˻���~�t�{u�x�U:�����$�� *4�L�A�lGe���'�A<0��.PI�n�0ټ�\�Up�E���?����?T��\�i�(z�V�\�a�d�d�jw�u~x1D��ڀ��̒0o`��A�~IO��_.�!WZ%h~�3.�ff*�����#�p�R`ψ�U
��t��iڙ;V<r)F��j��=-O�Z�LעP-����j9+��7fqlI�8�M��+Y_�y��#�sq�E%�u����(_ut�?��� �J���@WGk�2�9ؕ%΍k�$G[)Ư��>�_�/�F�-5t!�䂭�a�5�6�(��|���\](EԍJx�Y.��,��K\��H�&��D�Ѐ��Vyg�S�tC&�H�d%Z�Y�F���=J�r�EXe�n3�!�~���7��6�2ς�)z1w�X#�t�B�)�w޲��U�w, J��W�_f�s�����υ`���C
pNމZs/qL�����q�se,h_�ʇ�����@ї�@��|.���#c^:qC`�b?�X���6_��#���"�:W�oc��Z)�E���"\��d,~�ݍ~.*5�.)g;�e�n�&Ar�\��2T�OUH�P>�u��{�S�}	S:QxN�^ɳ#��K��&�e�.])�_%k�r�2�ѢW>8���"�ͿO�P�t�5�s`��ht�N �Pm���X��3V�2�`)�J�Y*�K"yԛ�5��V%r���h�M�h��(�Pc̭��#�ۧ3��V��B�E�x�)�E��|�zy�q��//��t.9�
أА)�fWW�w%�2T��6�s�: �rdэvX�K9COTv�����[����>Ӆ��%�?�:��6��O�o~����zL�ߛ@���$M�{����,�% ���
}uG�/���\n%�]���}�p��\�&_�1���.���Rx���jc9@��kk���L3|]�cy�p"��0�/�Y�0R<H�K;��_T��,IC�D9�~�FuBbks뤏�&��.�%�H������՚�o$n�����Eޱu��b<�]ɣY�V��n&:.�H�̩({�ƋKhƣ�I?1Gݓ�S��-��x,d�K	ûSb�(�\(�W� �]vR�����K�W"��vU��?�8h_N�L���.~h��	^뱇J���*g(���j:��[�/�sn�=W�N�eOe�]�0R�ߣ贄���@iE��"����ߕ�k�֕�D>�z�4T���[l�����p�i�&���ߐ�%�w��HW�1}&25VϠ}ݍqk[ޱ�+�����1�$:�o���Wp��)���˂��̈O�>W3����\6m�vP%������(�B�9�z��vB7���ZձC���rQ�.�>�\�/���M��
�e��W�.��K��E��!Q˹� ��jN,������@���4��!4nC�Հ�?a��{j���䲅/�<��g*��eA۞쌝��x�{.��r�tA�U�p����UCvvD3�\s^tb�Ec�o�of0�{�R�w.����1ͪ���}�ג�K��WV%b@Nń��d�;��E��z)hU̖��Hb�c�s��Z�(�`�^۾㤷b���>�C��J�N@n�c�A�bK��Y�RZ�|ʜ�.9N6FW-aB�}i��h�H�{V9���x���Pn��0/mYmսf�<#֖�<4%���=aȝ[Q��bX�x��m�����&����1��+��c�Y����(��iep�b�>hoh\�ȥO�b֣��4���0����!�ٝ]ڶv����5�=e	�fK�I5�I�4^��6��{(�a�g��y(�eA�/�53	���ǽ�����ǥ�Ge���c�|V�Ģ�L ��~�0�e#h��v9=+�������8Щ���Յ�1�x,� Hy���Y00,�{����v��H�w<�Q1��vm�{!��r�3�.�w������f��8����T)���[���������Ug���3hDfAS���� 7������Ҭ����,�e����YW[G}��"#D���j��	8��I{J	�`~!U䌩J.��8IZCU�YE?Xv�"ʪU�~h�4;*ig[�u���.E=���57'Fˀ��w��.��(~�X���9ip�����5��}�'xN�9l33��1�{<"���R�7�����U�pE�U�,γ�C@���,(��G���@K�ͷ�Ӵ���!
�$�n� ��Bs�#�M��[z�������2O��x!=�FY�������\;�߽ɠFQ05L�
s�uSm��!d���IL��^� z����Y�YQ�����ኆy�:��㺌g�:����!İ#��ƍ�|�í�~����9��f�Ǜ��)�Wɑ�+jE�l"���Yt���c�~7)F䄅^�7��ң��)���i[��9������$�]^r���+�?wM���z&d�M��i�[M}^�dy!�Кj05�s�+~�}��0��zv��C��Ӣ�0n�\���A��i^��}������+�~�k]�qvd��,�{����d���B^�fy��:i�ƻ��5O�qUMQ"ώG��gD��٣wud%�[�ÓpW-Oޒ\��5�+�p���u83�t�.o 	 ����m���kh���>����!±9�;c¬"o�-�_\1�tL�W�eޞQ)8�5]e���L@�:$�rY,h���6�E�z����ԟ�����PW��-��H~�&�M��hH��xj�8/Q�h\����ѓ�i��
�!�&��p$w�$Ri@�Vf��@����9adQ��G�P�K�*���@z��M�=9���Jڗ����)|��Y 2�A�6�jF��\�B��������G<.�������>��GV���|\��p7_�0�H���6��a+������ֽ���Z�G^�]�	Vc�>Qu0��S���z?��1PC��������<��]��(�,< �e3[�ˬ}MrVN(��~�5�Z]܀̲ �W}vh?����뙭�H�%���� |�^B���A�g�p�� �����:�;�aS�_�J�Z���(o�,1F	@DHM��椏�h�����g�E����4����Z�,����*\P�%�:��jY��sۥ�R�^���܆k�TK\��!��0�s0��`��D{|K�b ?1j�W��ǣZg�*�sww����Ķ\y}5	K��h�����O\�E���"M�{�L���H)9�����h)������Fn�s<T�K�Sg���W}��]���h!��3�NK	\b�l�(v)���	� ����z�<�.\��n�B`>�xrP$���	�/	%v�v�W�1�l�/#͟.PkZY�y����m��w�6Gj�z���.������(���!Ț�)��G����������2��2�%FZ�����!6�N 3�w�"<꒹�X�V��ykK�C�j��Y>i�릛�G�����J�)=8�<Pt�$2Q%S轂�zSmW`���Oe�x��6'�~��'?� ܭGN+�'�g<�=���l�r�B�9"<����U�h0�e���-�d@x����r����ti_�i��n:k�NP1�:�Ҙ��<e��s*�ߖ������n��w��s_�qk��W�Uj1Ϫa</�,���K�O����ŷ_��=�T��B�44�� �8��t���6C�xkF�n�c���.�j�p�|������|�`�)��\MX�ݴV_���;�p��Bo��h澵�C �E�d�J"�͛�����=Ћ>�C:Lxo�d��#�-�X���7u�R��:|y_�D��;V����������T���W&��_i���Z�Qp��]��r�y�||yi���4zm�	i�j��Hs/qMHȵ�-in�&P�o�G�ؼ�^\�%���F'>;�4#;���+^#���J�=w<��=*9q�N��v���=���gT1R�RMi�*M��ٽ��JH�Ad	˖���F/�5W�Jᔰ���\�2JZM�sK�*�]�b ���OA�-����z�/���#�.&
�n�|-����H�!���K��A��J۴7��{PG�dM�	�����'z�J{��u��f7}�1o=�$q]�TIO�3����I���s/]_�t��[�(�a��	���/�Fxk�X�zj�H�i��]T7���U����J
&Y��+��8!����]�9OS�?���{s]��� �A������?�Ĺvnf�렫��8�]x�!�"	�q�j\����kXȟ�#��ޜ��@
(��d�1Wl��v����L.��@��p���z��'2�C2Q�ͬ�I	��A��Qws$��1"m� �S7A~;�)�W�(<���됺Ii�l��������a�g":���Yh4'XN";3݃.�r�"�-�{�B�1������J����s i�Y	��`�����%y
,Q&�W����q�	5���-�+�K�鶗�5oWF+��q�p:��Z����`)z$�"�I������8{F�˳fwkH��w��RC�g?n�jfNa��B��3���{爽hT;�*tK�E��c(���(�-,X��g�{�ޢN���}�l�{r��P�]{�>&�U�aA�5�^������­@�֍�P�I���˦���
����ц2�U�@�������8��L��V�	�i�]S���M�G�9Xm;�5�(�t��R2�.EC�Q��WM
p/4y�&��	A#���h�$/�8��,Q��)'Mn�ݵ�Y�߮�9�r�i��0���2��L2�ӈ¶vs�T�K� �~]�ȒoU��nHK��W�A8�O[�2�v����H�MP����#>|�P�?��:d�K<�Ҕ:����=Ч���ut�5Ap�Hh?��0~���g�`w/qo��N���$�Kv�?�-/�k���|��+N
Ϸ+a��tJ�!��?��#`�S̕��j�%\��:���6� `q��u(��oC�L��N,�H���3�
����nCh9��޿����pz3�~Z�CH:s4Y#���n���Mɋ4�F�o�E�ʬ�x��	��K)@,�%Ȅ&:7����������y(��u�n��ғ� � /����v���� 7����{N=�_z]��6]��*���H�d2����.Q3D�Ue���7v��h1��b�q�vx���"|p6C�g������~~A���ę�z�By�"�G��������BРm
N��K�l�>_�N0�*�Z��P)!��ᤒ Tޫ���0E�˒�C�G�)����5�|�j7��JL��L�Oe9�%r�����O5��n!I(I��n0�NZ�0DA<.�ʘM5��J�U��3��"��ٚ&"&yQr�,kwf��C|V�>�!g9@sOmu���c��	BJ������ /8�́Z���$ 	9��۰�9��:���d#���>�5�P�2�&�=;|����	Ѿ�}�!1N�9hh R�/l{V���.1���SJ�J�Xe�G�y��~�H�	�|H�H�����k�U~����;8G��2i�x/3>�	�ݧ��AU`����/�)MB$�>�:E�
�K�].��v4Áq�6�^��MȜ 2��+�E.C]�=y�J9���ꔗ(��Lc�� M�Z_�l������z`+%�)�r��)��I).H��k[M�!��k0��%Xql��^���o2vpWkt*iLX>85�P�q����&�,��w[B�_Z�?O��)$�,��M����li���j��I
�������}e����p���Ve4����$9aؼK=�g��6`8�4���Ww�i}e�4�?�m���O5P �w�U6�c�Fv��?ԕ,k=�W���*W^�S���&Ԝ��f!���'w��T�BwX�f;;�,���a�u��T�qgdYeڍ!6e��;�b��c��-��[}��,�ƭ5�PY~�������ƟA])5���]�s�S�^�V�\��Jf�L���ԫ�@�صS����X��e-�Ex�:n��4�A"PgImS���~��H���V�"p��F�!bԂeJ�MT����6����e�<���6y�@H�iP���b\������G�O�a�TCr����Uи!@Y��2kg�C�8��9�!e�Oud���n	��䍆@�p����D�7��?�wq�
I���H�NIE��+2�S*�CC�Y��#0%`fUn�4�P���hH�ƃ�UxwOt��%��vz���H���}N�a�S�1e�b|s�M�e��-	�J}3l|�VЖ nʤ*(8��^2�/�`��O�8�3�H�ٛѩ��$��X�N�#� I��&FX��U/Y��OZW�K�>!��mB��\�C��=��/-����̡�bٷ���ַ诖��=&� �G�Rۨ�@R�U�e瓙f<�@�F��QNm��A�d��K�g�Åcb�Ch�Wf�'��ğmn���4�"7�C��y�ɰQN4��	<M�8C���Ҩf�S�
:�NI�g&6�gM?�X��ţ��t�3JK���`�H�w�Dj-�@<����0���=�[���� �_����H9ׂ*�bL��+r��>�$Cz�y'�vnm囗�t����n��+L��8�Z�ħ���UҬ��m'J�� 5t�����`������ӏ����@M�NZ�9�x�qJ��ߩd|ԥ�F�� M����"�8�㻲��9p��!{Jx�B�d�d���Ӛ��U��#(�8zэ�^Do���ޏ�%����]ud���P�/RP�v��*6p/�-0�H��y�f�+�R%_#6g�Gr��S�`UM���� �+N�ˌA�	I��H�UҲ����UE��?	c6ЍO!сF����5�T�������F�,!K��D}S[��4����3�2�=�*�ʁ��d��a|��*>'��F���d��8��r�8q����T���L�d�>lF���g�d�r�`����F���[z4����yHcʯy�S
=���h2hTW�������B�D���v�)��|���(Y�$�y`���'��L��B�F�4W�U�la�(�[��nF^��V�}Y���?Q�E��O�� y.�X�����zxO7�E @���u��17p�t�-�%�׿��G~n=��3��l��[RdTC�&߇�-�˘S�x<N��]b*���ܗ,��Fx�'��ق������=>��F7O��E-	��s<��ș����m˶]�'T �[�V���ǚ�q+B�v��]�����5�Í����26�ٯ�Ha%���#-{�{�$ټ�'*���S}}�MB"�ʱ�S�`_�z�rʪ��l`Z`�򈾬8 �)3ބX�j�`�m��ȇ�m)����y\b<!xԌ&�>Fd�8I����E,�z��#ê�#�F��9?8|�2Q��������_�r�)!��8}y\����1�h��T��G�]2�^��ɋ3	g+=�}�.C��|V�Σ�$�Q|�L�=�Cp����W4��3�E�A�@��ʾ
�(����RW3i`�Ąf�B� K�������U�1�����?��d��RCp���L���_6rwr��Ed{��C�t#A�Z{3]�4H�=��-��3	�kV�D�\�I�M�XXu'��7�}�j�J�"6xd���Uйٕr�8Xa��Z���m�u5�v����ܻMX�z}ɒ҈:
L�.�A i�#�ғ}�����ZBۯ����k��^m���d��+�/�^B��Р3�����J �Q����+��)�䰑��s�{'?p+Șv���-U��t(���*��ayETr���A�
}�+�����#���""�%���Ͽ$}5����� �3������)*%�Z����t��7�.�?�:>��G5���Y����hsy�F��7���l�S�x;��L~q�|���+;W�91�r[��%����kq��~���w 4>8{��U�� �����r����=��0i�T�E��L��������m��Cր��LK]'�M��'�S�_Ѩ���"�H+8l���,�*���>]��&�O%"��*���"��ݭ�P����-�YMi[�z��}��Q� ��Qo3(�ρ�LY.�\�5���5Z��T��L5_�(�R�6���X^xI�$g>lT9��.nX*p�dty��v@��h;>L��x򿂔�c?�J�cߪ��H�>(���%�δ���Wz�-n��x�`d�����`}�/@����F[������}@K��$��n�����+�G$��,-���{v��P4�����!��0¿��GT~�[�`����H!�K'��GМ�`U]`�i�����y�`ֽ�����?��߻}y�Y'�S�ٯ�'�����]�����F����*�c�E�|`�0�Я ��N!��uFl��j?uf��ݮ ���~�#��Ӗ��x*j_|�騻X���%�5O�I,	���z�҇-�r_W^ߠO-{!�\A���.U�\1��� mH��N��ltҧ�kJ���)��ޭV�
ꊋ�FBj��%�k�-�B��`�=c�+�
u�e���5�Z�[�uz�]&==С���D��fY~�S�N�u:'��z��ț
�Epi�q���D���iO���TO�e4��ͭk�d��Q���x!��1�o���`���L�Hꡤ�B�%	���}�]g�⑮�}��Z�.��|͏}H/�P�/�288�Rb�߮�M�6sg!�i�ؖ�Z����)5�5����s��~��-�S��6�_�G�2���i�d�x�t����]�^�:O{4�Զ��(�`��y<x.���k8����N7Y�8�QgWL�A?�]�f�.}���/'q�6_�G��4��=��~�� gK:����L�,���_ވ61 ��g�?�ڜ�ٿ����{!�����3���O�Ŋ�4��A��'
���B�$��2�W�ȇ	5Yj_b+����#�h�^q�t:wÛ�IK�7�W�|����4�xno�7���>	��5���uC(,|tR�ӣD��@7���������;��+T�i�2�/gÛx�+bPن 	LL���Z��o��l��ʠu��m}�?q�-k�G9��-֚�U�?i���cXդ�1Ȝz��(4Ji�4��L1�)NK���%s|�6���t�� ƗD+��@��q �VX�(\���Z���T����{�Z�&�V)�'��Hp*p1���Yh��7�����y۳�wTj��p�NZC�%�M�UO���&�Z�#	�V�aD�>JGV\��C�N-��*��հ<�>���_�C�A�����y�����{[�8�Ӥh|�����^�g&X��j�r4<s)EF{�����gy��{a�o�2�X8	�.A!+�HG\�$ƾ�
�+M.D��d8�k�8͓�$n�Qg[�L��h��~2����?�ϗ����a�ڎ�+��_�)��ł�������7We���%��+�qe*~�;�����Bd�V$��UUV�ˡ/��Z{K�<�(�x�h�*�!7_h��n�0�T�������@�	>d����l��0�[:�,�N��K}!�XTW�O^��4�O9v�+!x8(8|�ib tfփ�!���g��h��J�f�R��15�����*��z�to��I�p������S�Q�6���}R���d�r��Ɇ�<l2�'�S:�K�I�^��B�)�ٸ6(^I�L�:q��j�ׇ\��R�qx�>�;�£ӏ��6��a*���r���z��L�d(K�ӫ�|\_2��F�6tm�A�A���mhR�*!h+�����[����� �f&r]��#o*nU��5�j~w��3g�+����_:��	�����-ɂ�Q%��?$�����,c=©�EW���R{x�}a}�_v��F�Y6W��FXng��b͆NS�"g��/����\�L�=��Ć�H뮼�YR:��X���K�0�N^�?�:9���.m�TI�rr�ꓡ�	�� �k+L�F��KLԼ��%Л��ף�3�U�/$={mʡǖP�y�
�3��4�DҴ��\�\��޼SH��H�O�ձU���v����r:h1JS�� <���+����45(u�IP�B���I�<i�0HH�~c����ճ��)���,}����>k_br ��~�k6�Uu���.���_Ks(�[']7���Ae��:��L&YeJ�f�~���n�jԇR�گ��0*O����v�ѣK�%<�sK�B��T~�;(���q�%��N�>��n<���E�!��t����T
��;(#ͧ�y$-!���`���A���d���\�J���U��c���g\��r�|�g9܎B�����9����T����n-sj�������
��<O((�k�T�͈�޾��b�d0���U�=
1���{�1��HC�K]��ǆ���Q"��R���<F��N�5X����?1B��~���H�����Ln�c_�a�H�"�$6�]�(�)��pǯa��)֏j�f���'
c��v��/�(�O����e�/L��!�%�ٕ��+��B������:�����<��.�J�q?"A=���������p��Y$�PI�E&���m�9��ޕ���َ�z�[e�
�"����vE>zC"LW]��.�X�;��[e��/�wP��k���������k��2�Bũ3���j�ErE�B���ґ5̑�����>�ݤ="�@�;l��6��_�~�!�k�R�^���s���b����Q�ǩ4Gr66I����/�e�$y�޸�@��s���V�����\� p��y���^�И5��p�����\��pan��s�a�7�_	�����v��-+�Lޔ᪖�s3���-�N�Ʈ����y�}9`��')�_���%t����I9rhFY7��5���t^�&u�|:�_ҁ\���U����v�Z�s"z���w���A�"�y>���z-'�(�Ծ��E���4����h4�\H1��_�?fDŵ�~�z\8?�0�kx�(��P(@��X������r���,n5t�2��e_DG:���"]]P�����Ѩ��&�R��2��4�2�k���P�n�1���/�S�:){&n���.�6{�ي_x��հP��QsgJ ��vK��Yv*�3< kn�*cH����v�d$C�0&2�V^�o���qҗ`u H��a��ot.���;s,ِGC��ۭ�c���_U��ġ���m}@!F�9��x�H����|�D���7�WY�
�7�9�mZ��^Fi��9dE��^SS����^�t r�%��Ô)wB<[w��d�B�@i՝(A�O�V�lo+�����F `G(��&������jP9Ǧ���s�pyvY�� �ޖ�D^��Y����\��Ԑ��q����^�^���iuI���r���'�N�;�w&1d.�M�+`�&�gn�L �{D��/��Gb�<�s ([r:d��V�9K�ǻ��Y"罛�����k5�e�ͬ=��y_�6��:6ҋBJf�ܕN��t5����k
3%�I�و�n��H�-���*(m���������>��R��Z~���`����6�6���\%N�H���{1�uB���B�B����8N���{�٤�]O�]������c���{ZH���S1{�O䒲:M�u��%Ho8:��L�����y�T�v^],�}�7h�ָ�N����� c��r�>�uz����)��~��?%�=}ܵ���e�7(zB�[�a*㮻w��{��ܺQP�B���T�z���G��n/�O��kM9��偯�TS��޿����.k^����#_���V�]9��
����L���{���f�^��ҧ�+c�[�'u��+��2LLC�PK��{�#IT�R��"�-�����ؑ��E�D�mIÏ���sJ���LD%Eab�z�
UY�N�f��E���"%����V�XdK'Ñ��.�gćf��q���`)�������e�8SXv��.t�mJ�q������x�д�����>���Ӭ-F6K,w
����� n�I��؇p����/nOΣM8���2�������g��&c��P���T���ᱯn?5�g�S�j�0-����xl5�aV��R.w!\.�G��8�n��/�,d֑ ��@���;����l����x!��=�sH�������*
C�0���w'o��w�wl�3g�y���j��7��3�x�[dE6O3b(��r�0�i�R�P�\r�Wk2z�JO��Me��ڃ�N;+�B� &��y��8�����d�_��[O9�ݵS�]�� �ιg9�E�e���c��C�(Zo:Ȳ�}��زXj1!2M 5�4Aex��-�Q�k��oSt�����d��p��~/�|O7��S=W��Y�s�NH�u扽��P���!L��)��Z��I1u)�ꞥצ��f3��ʵl/��v�Xޫ�n�^9v�����Ȳ���?�/����N�yi76���'��PF�	X�o��]
)���l+tl`Z��0���p6b5h&��/)��)be�dX�}�f��d��Z��V�����E]�H�"��ߊ�]��v����⤫
�Sb���RK���;����*a��yF,7�A�[����5(�۱��1�8l&�<Y�PZ��O��҂[@�O�aP�8��K�d�9F@N�c�_�� �d��� ���mC��ꬢO �-�j�ֱ wly����fKnY�A�� !X��(Q�Y�<�}@Գ�b� c���8��j�gmǤ��,�ì>�.
̩E�"��8e֖\4�Ī��g��DR߅~�a�ީ�|x\�`���?l"1�/�l&� ��������QSld�� T��;T�A���
E3�a�����.�A�3�R��D��^A4��0|�����t8i!��>����j\[:�'����>�S8���_�^5�׀�	7�p�W.XsT{]lT�4����"�Ψ���&)z�kfg^�����q����$9��|��=9����M�H�?x���X|���9B������W����м摖G:M�M.̘�eN�|䋫ƽ1y_�$w� v�$i���f	J>Ϳ�V,
�JZ�i@�� �J�te�?JS���2��-X˟��X�t�_�7��Y�}1�l(�__�($�r�H��C�Q	A��e
X��6���/�{�GZ�1����[��$�S�ۺ��E�co���"U��SD�:荏�ة��pڵ�(u��	�$E��ƛȐ��W�o�o�3�����R:P�.���,��E��b	UT���¸(���i�]<PS���Uyd�˔��S=CVZ��s�������S�JF$��l9��#��b@���vJ�|� =����$I��
Ydl��l9mi��F�Z;��!�q5�L�H�~�<@���o"���� Gp8u~�m_B4���))����ᚏ�.[����D���L>dz�����9����`}��(�z�ذ����9�:¯a�� �$
^7�0�PD=�?��V!��U������v��r`_7��:�sK찏������0�8g$�-#���ٌE��l�,ܐ�J��cι�ގ�!����,�uj����g�Ԧ묨Y���1_��RMo���5�B�k�z VI�%7��TH���G���oV�v<x� �ۦ���՘�
h���᪢̡�(@�''�B�*�»��7@.~�8��Ոx&.V}��9E��;��i�)���w����Y��58�M��2��]ujU�����'Z�7-W�#p�w���gL��#�6����z������ȿ���r�_������JqKXibD�*����z���ʿ�i�t�����K#�t�U"qU�9��x��Y�R� 'gl��Rv8r/����`��K�D�׷<�>�ɴI��5���4���k6#���eYZ
}�FӦ9�,�O��I�Rh���Y��
@<�ך�T\)oMsfQ�H:�����~ںE�-$��\�J�G�!{��}.��2�������db�gw�Bk0wn��F�LB؏x�My{�]���rl�`�/N������s�FWo��O!�[Bѫ���b�Dx��ޱżfh�sG)'�M=��4\2G@���s�	:��*�������^��K�/,m_F\p�$:��	b�q��g��FQݍ�c�/�ve��ݲ����c��f,Z����� ���∈��T��0���ircV�6�k)6��I���txpjS5�3*ZmB��$0%�i:�މ(�1��,���rnW'"$��A��|7��2�k�_h)4~ ��}�(��.N�G}1�VG�F�Xb��*aφ[Q
��I\h{="74K�YY1��&���k-�z�r9<���%�"���*��T�ݐH�1>`���f�B�1�]B�̪�F�o�إN쵕�z:�T
@�\߀(R� ;�����U�)��)=w�,�;�Ti����;և��o�%��v#�g�hs
��x8Q���54#V�4jd�gp�bİ��^�u�i��ih�k�
'�a�f�n��O�%J�%B|-m��P���7��`ԩQF!kE�a���ݙP��^�?�qOg��]׾�o�b�-jO8��I
C[uS��O���o����'0H����¾�N-�*ǭ�q��m_q��T��,�ã�mr����&\�J
�\R؁q4���s��tt9���'������ݻ&�Fd�}yZrT� �a-�/�r�K��cZ�3V��*�W�Ƚ5K���]a{�@k��㳌��4?�0�Cj���f�# `l���.ч��� ���,��仇�pEv�UI���\P��	��N��e��45s �{��p��-��b�v)�,e�S�ǂ(�yߟ,1�0POظX�Dn7�^)*.G�DSdv&?Y�M�ܱTB�E6�9��G^V��`lNg/ؕn.j�Q�Ԅ/�b�DI[���V�b#M#!�i@��o07�[
�h@T^��9q_<��tc"|�Q��ˀ�q^�4������j>^��f^Mǟ��-p�<	} �O�ǡk������q����J\��̗���ϣ!O�R�}�Ē�aT����t����p��wi˘Z �Nbړ�Ʃ���0��|Hn	���&-=�T��{.�"߭ o�Kټ���qw�����u@V^���ZͽO�)�A$�\��Q.�p��/S�}���\��1D^	���f��2|�Һ�Կ_)�e=��s�Ѽ$p������v��K����v�? z4��.�R�ؐ��2�q<��:.�[��Q�I��4�flU<��6zs �� ��!��U9*~:���E��NhQ��]����&���Gh�� `v��X����	��S��=Y1+��_5��_����,�q��VniZs )����A�ccX�ɷI/!�M���_fx_p?�Ŷ{4%��� ��0����Q�|T�F^.t�{� ڲ�j�;�G�U<�����}$��	�>���CuIl:C۲��|�>nC\g��k@(�����������E�*~�a��d	�E��W�ZE�V���Z2�=������\���W}F���"��5��<I΀���;��(�<�t�C�;"���]��Q��"����}`ox$�P��t� SX�F\q{b��+Z�����_v���{�U�^1u�����T�/�ƥ��{w��䒮�=.z��s�v���EQ�n��"����%Nx9��S=sD�?u��8�-�?��V#h�O,�X������X�p����>�	y�#�C���ӡYD[��?��Ys��i(M}&��µ��z��vve4U��k��-��d�Fr)��~e�{c!ㆸi��h�$�^�f�%9bޢ��8�O,(�Q7t����^�Xs(�[�fF����逈f��(�M�P��X�0�E���fM�����,%����M���� Dq�z���S(��7 �U��4�t��~\��W}k�NN��L�DX��t�h8:I�-����Z�&�4�똬\'�Bu�z(��]�mѽ*�C~�@a�'ճ�����m�*�:��4�<�7(��ϔ]�wϛ�&J��6~���L��5;��`�R�ZR�k��c�Q�e#� hI'��. ���Q������W�}w~��6cZ
�p�>=�
[Z��.ۇL�	��R����U�t�YUtom�y�D���H��3�JtWT0���BD��xJ`6�.�Rj>l$X'<��A� �ЃYH{���MO3�Mǉ7`@�-��*�;Dbf)Ǭ��#(���í�	��΍�� Q;v�3W��(b�� ����*��w�O�n�лX�L-"�&Y%��Ѡ�]�A�����#�dsNn{����(.����M�Ţ�x�߹�7�ó�� F{���>\�8욃���[�>�O�Y�ezh ̔J��Fۂh���)j�4E.��C*���2����Ls~W�*r�ھj�u�����0�t�P�&؞a�*�??��coD�A�ɠ�V`-	�|+ n�U�,ZT��pi���!Z�����f�R������ZILl`��[�Nu-�k��a^��Pr�b�_�T�,��'�{����1Ǟ��"A�~�,��2qs��A�.8��-�kNyN!!�`����U��0����s���pQ�Ԓ�꘱b�1 �t��x��h����_[	��r�鷨8&�B�ؘ\Q"o�7��\�?���Ob}Й�\����?X�fD��Y��j���5�an5$�]��`HOKs�R1��,�W��\�-j��na�zK�[T`����M�YF�Z8�� ��{�2�Ԅ���&�[���~r1���q�E(Q
:�g^���?�:�l�㗮���R2���+$��f�)�EVL��-�}�^��?[,h� yg��	�ta㥌��-�AF7����0ϋ�
�[3�|:7.��_�_#c Di��K,��N8#���(��K�_�`ePL��,Ko�E��	͛�����4��	�ь܆��F�\)�`?qD8��05�~���JR��>����%���KY���yg#J����q�(�`V�$�K����eX�A�"]��GD��¶��~)2`9���m{��L�Ӕ���<�T���D�3�W+ita{�s��ϕ>(l	��)@�"�D�����˳?�8��ϧ����Kc��S3�u��I �e�pK�L'�d�g-�"��:��#\����}���,��&l���}�ocoA�|�n!,�8b�R_�~��ʜWq�1LNYk�?V�N{����n�G����]Q��7��	5.>J�ƞ�N0�_F�r�P�2��/j�
̡}2Jq�.�W�Ѝ�
�G��-�6�5��\DDu�D��N#�&Z�]�m��۔�볰ݤx͘x-"4�6��ų f�p
�S|:�^ަ�I���S���)K\�V����L�t�M�-���}��������?� ۫�� �
!�1V���l��y~��<!�E�O��lQ��W㔔4�{3&;��LN��S:d_���_�@�?�(y2E�������)Ezg��
y���"��p��L**QV�+��(��>�=Ԅ�wdz��a�7/����]�g ��������-_�Zz+M�|���z��U�\=3q=�4�r���ΰ�g�� &�d2}��8u�yYF�f}q��h>�BdⰇ��0m6)6�˷h��5�ܓB.R��=xi����������d����-�6��خ����т��P(:o�����0=tny�˖hɞ����H�j����+j4(��RT��C0�	ͥ:��� ��R� ��#�!��V�M\P)J�¬��0@p���chu��a[;p>�3���ls�n1�L&aB>,��}��^���9���)@��&�|�>�2�
[U�xlj�^I^3o�BOHS��&pM�t�$"��i"����
�[ʇ
_7S�^��(��
�ý�_�7k�]f�f��Zy��Nv�Dn�����V����K�8��Y�C5+�r��n�j��4�8�X�OS�����e�,����� �ண�U%7\���>&�֜^�]�D�q|�6��U&�5���1�
��}���S��M����B4L��� �fo���ǧKC�4^v#}��y2�>�$�;�5�&�W!!�������g���<z\�~��" �j�9&`���%�\�D���&��u�x M��x��[����:G�ִ��Y|�='�?�V��_�}�0�]����Ap�k�;õ�Е�۪%A83�BV���Ԭ�b��$@�=�cH�x�bݯ".���7�}�%���	��RZ~s1q=�ڝ7ҭU�u�nD����!�� C׮`�+�\����Zaʰ��]{M3����4��5�Ϋ��G~��D��V�|i�=�����W�Az�b����f��C�{�ɖ=�u�{"h~��I�;��rI�|6�¹p�r�V1�3/V��`O����Fr�"��)�'����������*sʫ�-0]�v�i8�G 4U��]���֧Iڱ����Ƣ-�y�1�c����6�v���p<����4��V��G�"9
�|�ll�̀���p�O��T�	(���gC��H����n0���X��.3 -a����n*���[�V(�ý[�G`iVTƧ�3�Q�hM��R	֧vȚB�� f�O}��?���ɲ�/Ɣ�O?���5`H2A.��b���O��Ơի���.Ȍ�_Nm,l���'G�s�����d����Ys��C���7�/#�=�+8�摀#����#���/#�;��%#ڨKQq����L&��0q��-0�|f��:�D﷏6�ڎ�!u��Aw��B��'+����ŗYY;����Cᖬ|22���1ױ�I�'�\ѡ�Dm�Bjob�����t\25�=�\���&%���]��*6�P����~�p߯��Q��Q���\lN�bx�!������	I�B��`�˚�����2�͚뗧f�Ԡ�q-+�\�R���m|y�Â�� �yyO��Yo�{���׆��~S�O����K��bo��HL��񃐮�M��I�_�=�QO��?��Tup��R�~u6
�A�:�7I=w	V0��(�D�����^?o?�:j1_�e�����^#�ݏ�Ş�֪�W��H���1�D�b?GGpd.6�M��1����fHo��WﳉC����Y�Oh��g87��+߾���=+S �83�6��G_s��$ѽ�g������9�J晟��
nI�1{&��K��l(��b�pX�w��ж���W��T$�<�O3ήwL��0L���s@��;$���;5]�PY7�*�E<�e�:�}�_#�Z}�4�+����~򼠋?��.�P���!-E���c5&�n����h�t��G��"@�	� ��USƈ�a;�N{=c��fL����������Y+�Ѿ�LE�ff���9�8���Iq��S����"T��'T��~������4�t��I	_[��[�W��|�U!���
�U�~14P~[G�]��똁|��fK(���G?�-G�>�2T)�ӓ�f>z��l�u������V��6|�'J�����#V�z]_zĥ�p��#=g	�̃���n��c������p\�S?Z����ǀO'��n���[Od�)=��)�@z%B���߫�ک�<��=��g��\��U����-���n%�+��Ri�a��m�z73�/�(޽��~(�h$e�nъ�=�0#U��Yt�M�Jp����POV�.�5-s�YznD��H^{��UM�M��d:7i���_f\j������fM�c�;wS�y�t�9�f�X��}UD�{��n����9Zx�u�h�7������i�Ӷ���6�I��oׄe�-_m�����\������<���|��|7��GG�S&[��p�/�ׁpZ�Р��ц�bAc�9{��#si�s���h�)2	�ޘs�8�O�����R�à�ȉ	 [��sl�vE�rN��V�ec��f�#9��Ll?����6>��*9�n����v�n\%ܘ�C!�L���ֺE��M����t�z� $��\~��׿��~�&疘oj�W|�*n��k|�7�����u���Olu����f��vည�eG�pW���j�\�D�캇�>��R������u���l'�u�c[�4�V,d�n�?h���jAH��G@��t�A�ǁ�޿�qGj�\��zb�j�lI���Y�T�����^Ƽd����0q&�.v�r�J�L��k�b���������k�	(��xw0�	�ca�K�},�ܬA����?�;���&�mW����I��DG�b�L��u{Z萓 M�Ht�ȯ�o�C�}ohz�=w-�]��b"~��_�i���q�,��\X���-(_!-��5-��{���3���|1��VF`wӾ+�S�L�/F�>�cAT�����<��n=�����N��Ǿ5վ��r�$Y?�Z���*>�}$+��-�{#��*7�	A�O�G9�z T�r��Y�,g
�����-�Ѱ,&Z2������0_4���`q��Σ��Dy�6Xh�I���!��Xw!ac�:x��>f lGZ���%~M��u��U��y/υ� �n��7��H�0�Nx0+�j5�Ui���2�A���ޡ&A��Z��k��]�1�#`�\�Kܖ\^�/���6٣RQf��1v�@z��:�a�T� i��vg�$�\�s�J��d�n�y��2�d֦9dw#��W�"~^2�.2Jb���^��\��n�6㲗k��$xZ�@E���V>��kf��N���84�q�v�L�&hpF=3��N�w]Z��%\�����5ޜ�%=߭;��F:K�X%{Nn�*-T���[�.�V)-�N]aJ���\t*�yְA�l=i�U��ַ!ˮ�:pkp���,Q�7�M3�ay�5z�����`���^L+T���7� ��(�r��X�t4�.�҇m�OX�(A��A�Y��;��b��d�T����U�֞�P<1�2��r��f��q����o�kcQ_Q�7Ԛ��qt�2�D�'u��u�y_~�Z&LfN�U��t{-�8w_���-ɡ -~cޜB�Z�kY�(E0��=`&��"mD��pC#�T���������bF^X��~�->h��W"�Ђ͔;�c5���01~#B��jx�CK�k$�|H�%�P�������)�;����f��wX��h$����_�O��Km��ԣPҫ�� 8҃m�k�u�\�z�l��5Z�L`D#�΋j��PPMt�:=�<.Vģ�ےH�q����=��wD��KC���b��ۼ3@K��Dv�M��.��S��P��n����|��f%��ȕ^�D
Si����_�9�3)u� 5�/���ؾ@S"Xҡ�u�mo�6�p�'P��3��߆�������F!T`��^�b��ќ3�,x�S��`�B3���������S�:>A��z����'��P�����q�e�tc8Qpf����̞����IU���H�Ԩ��kLɈ��Nm���"�V���

�r,����'�eL_��~�3X��׏���O1��WI�k��ƃ�7�Dܩ7�ݍV�J�W<����@HFM������4g����A� �:��<�C�s��a0u4P�!�<��S�=q蘼|��n;w툉Js���5�^Y���7>|f�KBH�����+��2ʼu��ѥ2��'��@�e��2�Ȧ���}VB_�l0�n�x�ssp�pg�qyZv���dW��Կ�{��q�B8�u��/3�@8bW�V 4�Q�b��3�����WQzhʹ	�����D�ba�i!E�G�Xl�}HC���p�%�w��n9B�ܤ�I��F%$�Ws��2veK����]�r���S�^j_}���ӽ�����o��{������As)dqueNA�)Q��j�y�d~6��4(��ٞc�Ed%�sĵ31�N�C�� ͯ_�l
� �Y���	�0���=�[p��&1���n��2���h)�-���-�8�����y{�U�SpQ<�d�?��s�k���`3�Q9hWk��|3�h&3�j��q�*N8|���&󧷗)���~�OF��.z"�2�I��O��)��M&~;*�C��i��0��A�u�m�	�5�>mZ>��C�؄�Td��gn�I������ErѓV�J�����F�F��,cΕ�X� ��v�t`���8h�^���:0�Ƌ��/p �PZ�W,iG/�<�|�?�
�;O� f��=��l�i78H,J�8�+��&�?�֬�Q��c�.�z6��vu;c��z�u��[��b�B(*�/�]���H��Kp=�7'V{1-
���wk�˻�s�y�c"���uX��N����_<	�(��;̈́5�e��>�p�&����?�]�g�/���x���7��v�L"a��'��:J�OU��i$%h@�G:.��[6>JI�pIs<�u�{2��v�*p�N�!u�/'G�Zr�'���4��d,(�ݎ	ZGks�/|��&�[�]92�S헇v����qĴ�r+����.�~�A8Ӳ2��}7EP�P��8i =[��<�&�H����-L���Wf�|-���-�����"�'�!*ٸ9�l5�?�٘��Ti�%�'�쩼/�h�*�%�p���^ߝ���15ORN�.~��c�ہm�� ��vb]B,�}�|���;s ��ص �&��7Ʋ����p6,�|�x���pj�>�S��~�Ě/���>�����) �R;P�o)m�v ���|�^�C<�z��#Zf�?`<�d9]���kӿO�NrѬ���pb�$���z���gũкJo�4�#Nr��.	h��ޞ�8y7seq�@.�$Ig:������!��"M��F��A������_a�tz�[S��km�j��gJ�N��O�|�	M�J���Ʒ��T{^R,h5�==T>�}�iB�JY'syr�x�+���g�	�ck��4#k;kl��o8J>ߡ=����iNl]*�f�y������_�8��=1+�4k�(C&*�l[[��&`��T^��[���������|�m�����!�'?����=zX��;�2D�P�~�"�~-"e";A�r,!B�� ;DA��%.):5�@Ep��l��cT����#�GJE�8��6�Ob_l]����W��޽� {\��n�o)��(���,�&����J�}"��m��d��E��v޹p�1�	gN��'��h��б�����*�AZ�ko���,c�ZŒ�A��@4���A�<�� L,�,��$b�&�_\�>,�X�k��H���/E��)�!��Y��"���T��me!n?.�yZg�so�sLOx��0x�?���Y/� N%����]�a���̺���� N!r����K������-*1:8��&M�b��c�XD�T���Zr�����M�k��;��1�g� ��AH�s�Gb�4V�t]lٖ�׈�O�f[n�C\h�o��o�k�J^�K]aɢ
�Qlף^�4E���DHu$	X�p�2�D�h/_��sg%J����f��_ �窯π/�}�����t�%�R�MoG�d��R !r>Ւ+(VpR�xw���B��4l�H�j���y?�Z|F�B�|��+�ܥ�����_⛏����5���]"�V
���mm��;{�M������e��^����5�uVjzKTf� �߮�x��[��5z�P�>#�J	�<�#�9�.U�y�'	��_��V�!^t���8�� �R#��Z��A۽����ʀ���3��Z0Lz4䶔Z3/j������oy�V�'��/��iF2lR��>(5�ݺx�ě��C�?��`?���u?�����>�S#�����ea/C��]�:� �E��,�1R�2:����>��mw�ѱ�֘E�h.����u��D'����"�G������B�:u�jw�^8�*H �f����V�ުK�Y_�@_���!$���	���!�����6�"��?����O]���BG'��b���]�`�����m�r 4|���L��L�=:�Ŕ�O��|�#[=Pȉ����'�},�)��2S,�P��M����%�~c�<��?81n \W��Ф�=�1x����݉���V�Z��B�%$W�'e�ujq.P!RZ�nt}n��ꨡR4x�;����S}v'�q~�#_��u=ï�)u�Ʉ��Fs˕V�+�װe�?��m�/���_�*!���uh�ڗ����,u���>Ћ�BDit��6#���n������#��f�­f�&���n���D����v,�a0�M�2|���>�|3ُ��Dvz*����6Y�g~'�Yӑ��Uf��@|A�g���:�U��Z'��$XE��N�����}���e������j��2����Ei:H:�|Yk2n��9��O5��O��V$�dT�y�|�)�Pϻ�p[�/�K�W��7����5b�1�<G�;�Iú����U�O�z�{&�bbl)�$(Qs���$���/�?o ���
� ��/��i��fNw%��w��>���%�f���E�:�y���R�����3~�v!�6��h�ĸ�:V/xr��Ho�7�;1L�愖y�����,��&����'��,���+��9a��c�}/���N��<��������WD���� ���i�O?�F6�kf�/�D�]�2�e��e}K)Iڃ�c���S������rKt�+_쁿hOX���P<�W�O�Ƌ�nl�?���'�]����7T6�M��zq��C7���5�ANVhdc�%�ec%��lfW��D_�Z~��^,�9|��X'~T�����%�~ �:=��!��hb�<;X�D3���J@�����+�z*��<����A�f�Q���g)���*��`#��$�E�J�87 �9WZ�[>���A�������MB�}�pCY`vr��OʁG����g`<�ͅc�(�x�4ao��E�[[��W�_]6��P%��B��4��C�^v���XEP�d��C���(���'���T��/�5C���U|t�:/t�����0��;hj�y N��Sw��&�
��7`&�O���tX_�R����Y;"z9�Ӱ���U�
hO�r���|��^r�Ԣ�F�����	��١��T̢����!v�u���	�H|_�D�>m������AXC�j���6m���ۑd��FW9�=:2ża4e���*�ՁL�9�FJ@�!����4	�P���j @�]@CB9�|k&� �F�����$��A�B!5����o{*���(���Cma��r��*���;����ikJ7�z���ίխ�����T?u�[F�yo��.=t�5i��9M���`T�%� ��ӧ泶�%)���p��D��Ѓ�5	��@v��s#���~9vz0���Bq��l[2�\�<���o0�򧁋�Z�&ą�f��fp�f��K�G�de�"�D5�o�g�c�
��W$��KI��u%}ZmF�ga�@�Te)R�h�� 6-�b����ì��,/����M�������!�3`U0����÷�]�Ͷ��1�q�G�oK
�%�M�A?�z���Fd��p9�����j�u,��f�|��mK	x��x$�eOPR���r@_����J���eyF =�Ax�W
d��y�0��4��)����_b!��'�Y����bΔ4��{�1���+�Q�k���5���.�3�e��~A
G?�T�
�z?�r�$s���
4kPpA�2�u?�54e٬ha��ܪ����+쫨���@�ѻG"���z���ɪB9Q�S+Z`E)�"B��2��3x9}�O�2�R���K\���LɄ=^o�ϤMg�5���Ot0)�F�AH=*�'����zs�N&�e��,�sH_*��,�uX�k).�//���� �5[Oޕ�39ͷP�?g�%�}S-K���rX������	�����c�u�!��ջvs�2�v����P�Bv7��i&�5�)8�*C{Eٻ3֢X
<,��F%m,!�u�Q�л��l�g�!��$<�v�x�O��{��U�i��R��T��p���f�r���[��>d�=]?-������|3�b��@]�2�>�VW��*�^�n����F���:hX^2b��B2>��V��F�h��tո����5	�A{���4�>�	��)k�^|�G��i��G�#("�ng�*�R�!%i �;���.���&�<&J���O�����K)�UGh�^J�s4\��)�����x�?�f�WWf�z)^2�<��ڌ�rΩu.k��)�$��b�4�(��z�,�d�|hp��̰�q����B��\Y�O�k�r���� \j���P�57��͐ݙ	}T��fQ���79����C�3:!U�y���m\�=ڊ	\ޮaG͘XL,w���p�9CE���%����pL����"�9l���L�L$��"���P���sJ-��8i!�}4(��Le��P�@��p"aP�2v��VT@�\s+����Vi�S�S&yo�I&W��|L�
-�����|�
��]cYp[f�M��Q[��;����p���Grs�l���j�W"��j.��V�c%��M"0�nn�
�I� ��NәK=¬A�2}(#SO��վ����x5+L��T���C�v�ڣ ��+����
�1W~cʸ
�-V�m~�0Cr� �+����7��@�7[�T���l�z8to��+����7�żx��er4$gGJ��M�J&���Lr��[��\J�:�"I��2����_*N�c�k�����$�>�qWм��_k�mPIs�*�M�&F��Z�i�A�3�u@F�d��&Fa�eW�i�FV{�J����]B|��SF:��q��=�9������.%ۂ�+y���h�(4�ػ�WX~��B�����V1�H7"^BR[̼���z"m���S���C[E�O�����8�i�$��j�	���9�Vo�F}�b����3�U�G�~�'a��9�@�X"�eI�����p����v_���y���J	e�N�\&$�+��3 ra�7LNz������`r�.Y�Lp<w}�Y�[�[�( �)/=d=�#�$ݢ�xD�{�P�e�Ȳ����T���A��ET�/p��S�)����/t4�d��d����)VTb��S:G�c!y�c1#���?�b���q=�6�8 (j3J-��Ax#�E{@ǩ�ܠw�7�/��7Q���`�E��Ea�_M�!����*��C_��p�S���g88��)���݈`�+�;3�(��+�A<F�'(-��JK�+R)��8�Z�����gqE����x�|��!���Q��0@H�P��R�/�C���I�z'maS�c�6wd�7�7 5.\nxD����Ƹ�����r����;���Ps �f�[9�[�&�\�q�qM�	&P�۳����/
8��K���ŋm/"�Mf@��W�/=X�6�=�=4�&�pj��|���<�>�7��8�2�q6e/紌���P�BzD�?q��-p�V��(���S�@���X��V�Aj[��}�}��x�d���>\Ot��M޾I?�!�� A
�s	i��y�D�(�q,R΁�]'Ԃ*
����6��b2Qm�8/�)��*��!����h�]��(�� �R�`h&����:��Z"��9fI�mfқz ��b^t1�X:kb?o����	���Q[��i���)��q=W�@N��d�4V��V�Ƴ�U �ί�
������:�����k���1q]�ϰ�墬3M��s&4K��amC�?E��z�t:w��	�t��X!]/����L=T��B���m���O�4@��	�M�r�)n�����o8����B�~�:��P�Lo��ͼe8���� ��O�髣��r��O�~Z9ZҰse�t�����R�g�ẏ��xZ����!�\�ıvx@�P1���í"�ba���"X��$x�LX��\H���uWޞ�d�僄,�y�?��=�J�j�h�bJ��b�>*��w���fy��K ��J f:Ի*ǩ��d��<x��1��:7gUdJ���ˮK�b����t���5�P������H���y��Y����pÉ�g�"�@t���(�ދ_�0{4gLb��ǃ��B��^�	"��q�Ek�:Ŝ��Գ�.߫bJ����g-0��R����;�u����KS��,M�����sD�r3a/���Ug�m�GK�^�4�:M�*�u�����Ӗ�;D$�9��8$�5uÛa1�{��~���#��ifI笌i�_O�F��v 
�n���o��~�2H�aӌ:����H��TK��p��8�
.H��ۧ�>;�ۆj�C��1O�h(�,[+[�C@v�"3�p�C@��>��~��bt1n�'�CH���B)�-N��.�Y���e�u�Z#��P�s�aXV����nS�q�u{�B	L�M�l�����n�;_5�ӂu;ˈ��#>�e�(����G��F�d�\���9@�P���*�u5L`�������"�3�=
תb�v��W�S&�2����$���v���y������+��l�W�i`��n w��f��5�C%�F�Vb!�-�š��F�?*uɟPiq-咨SCh��&M#��\5@>.��S��S�;�t$}��4�É'5�vU,�/P�{윲L��p�j���+��M��.��b�9��ōo~�I�C���J�cҏĳ�l
4���M#��&�OFiQ�M.��~p,�=ǃ�?*������}[�)�IG8�I����do����sQ�ST��oV2n!�)�qH�\F�W��@�>y)W��c�|L�P���Hc4��T-�WD��ݕ�����9b�;&@�ᗱ����ȳsL����x��w<�%0��ٰY��r����P��!5���]�W���~F���lOP�e�����w�i�y��Q��tl���:ZI+�w���fĀNU㛞�c18�G��_�����<op�a� g�DH�a��0���y닑��0�3��ܭ�G��9�D�к��U���/��a��g��eZ�a��c,"��2�?��r�� �2�����/ޘ|����IV��!c},^5�������r6��>y/�2�9G�:.��1�'
��lwQ�@)Pvw�ĖGjf���薝�������=e`ۣ=����b�{�K����<��W>Z>�V�>�;�Y�&i����uc��0n�б�u�w�@�M��`����@��j`��T�y��B�*Ƅ������+R՞f<�� Z	|<��iD���6��Y��[��.%�|�!���N�g�g1�q�a��`��J�x�n9-�`_�
�RO�[c���͖���
`�\i��<�r���)}ܣ*��JV[���,��@��m���@��3g�7�LR�8����:E/=\o��N���x��U[��� vb=���VK�FI��=���j��|?�z2�8� s{��Y��eL����_~UX���}_V��]����4��ϞԇY��ڳ��9��z��;M����P���h�'�K������HԊKK����XdU绦�IM:�n��'���G��l�T�%�������Yz�/�`�p���������ÉE���,�c
�X	�۹n���'�@U��b^	��U/�����8t!?�.�� �!B.b���.ۯO�mW6��k�@���b���������A�o����t�N$���%O��xD>�gIL��^��`'v�����S2���T��*����!�M­Ęό�н���e������Ty��z��y������ ���4��l[�� ��^z(-6�Kv��k�2dA_T�S���)m��(��$u��LӮ'�j�B��Z��(ʃ�f��n�,y�"����ER��nW[����)u�]օs����9 Xz��v�˃i�jP��˞`e˞g2�;
��2��-4UQ�=�V�f�̐��I&6���d�J�CQ>�K�*���[�/%mg6(�H�>�]��/i��e��N��ʙ���ؔ С�Q���&�K5��Hƛ�]�^&�s�|;_���Hȸg�0����3���G͈�rl�|�~`vm���O� l�l�$CV<���=33k`��Q�p?Z'4s�r_f��Ds����-v�	�6q��|t����4[?����f�ˮl��EX� jQd�I�(�IQJ���ReH@����Ӣ�|8V|#_�6��R��ƭL����U	~�j��C���le�tx+�����QVt�=1� }�ѫ�Y��^�*}�F_3�V�\I���$�x���^�b?���U�=J�Մ � ӵ���`�t|�Q�q�����/�� �QG���x�Y��M����1������C�yoG�K��[����P�k�B����_]C��/[폵d|��9b3F;�YF�#��sQ��~���e(\I�N@qH�H��kFW�i�5�BvK�f!�ȇ�4*��������)�G `�7��-��aа�l<Y�߆�}$���crъ�!X:VupD��)�H�D��cjc�������I+e	�������
U���<�/|���f�ADә�lEx�|M|05�6�F�s6�ﾞi�]
56���j'Q��2ʟ�͈u:�1��-���H"r`�,�|Y�i�8c��-IY��\�W�e~��cd�C��W� ��%���T`/�О%�x�suϵ�G��p9#��\.�鐹�X�\�Ad֞!/��*�q�-OW��>38�C��*��^��ɺ��}ω(#�~:QK&�鵩��K��	G�R4��!zAB�I ����� R�T��o�l�#�|��#��Da���T�� � gh���L	T�d����T��<?n���R�����Lӛ$�e �$گ5vfx1Un&GC��7���"���� Ƿm�RA�&�#	���4^j{-��'w�2�d[Y��K���DE�e���T�k߂��kzܹ�4бh�,�W6�GUjҵceW�d����/9�
:��(��㪅$5��H�b���C�M&t��	\3$�3���k�4VL��$���RҾѴW&Cg	֢�	��bA���g��Y�Pp"ci$ρq@�R
��'I>��C �T�7�#�#j���}��T�cqU6hB��8�y7��[e�!�#����{Y�@1?���e�?湮�E�n���ut'��]՜⩟��*�@'�fO̺�7`�Z���1����"���7���#^��j�4�nl�����Hg�_ I��1�ԯ���
���SL����J0�N�/l�}�Y��:�2*�����s��h���..��B8/v���`6і��Q�OW�@�~hs��K���a�f�!��q5J`C,Nbo�sE����z�<iT��'��{Xo{���7��
̩�.&�X���Oך���dϳ�إ=��QWVC�q��U��na+ץ�������f2�_�ԟ�������]:�E z���$�䇔�Gq��9��A��ux����M�٘zbG:���"J�\�f�KKTgG��]�� �V�ѐQ���"�sZ����� �VZ�E
���[�(��I\6~�
��r�G�4�E�p��a���%D��p,<l�^P7�,mV�'�&�6h�+谀7SQ������p\�AZ�k_>2�~<"8��%Z����vCf�p�5�KL(�9�*ؘ�BH;��[��,}^;/ �`�X�*o��&5�9��ڔ`� b|K���TJ�	���05�\�ĕ�ɋM���F���fC,-�G�B�k���Ns��|,��Ik-���,���d��g�vprK�bW��"5��QiW7�A��j�?`"�A�fM�L�o|����P%�H@R�&x?� �Æy��ㄘX~Snw�>��ߛ��:�tEM�2�B�J��.��?�W����KX�l/,���z���'��4'��`곡��8Ec.�l��w��� �0�7Df�*����I����wfO�A�Ԏ�l���J�=�e�h4�f$c<^�;wixG�ѻ���k9�X�t�
$�z
�@�56;��d��H�1��r��a�D-�O��R��÷,��#%'ܘX�jإ�id�=�~}�)��A�D���ZV���D�z�N�:��$��v��D�M!������]^Gţ��3m����5���?�A����iH�Te��iB�&*�u��ӳt;+�FH�AA�-z�m�A��@�n��hl\u��A[��w�蔯�L1Z��ʠM��n��?+���`a�B����k�7vH��}��� v�K> ��+�5��"����l��	Fc�C�Y��HdQ]� �<��5y���hk�9@"氚�������k�?�b���9�.��c����/l�Cu��18U�z����|��OL��DK���ٵtU�x!q���@�(�r�QnK�5�𔥈�iQ�3���J��C���Q��%�q�:�J��K��jGMk�lX�������%�rNaQ�I5�w
�?�E2��˪^D�5v���w�[�g�;���l���j�Eʼ9ͼ n�2�i�k��~k��{��dnI$3#M������҇�g/�q#h�5Ox��B�h����6E�`��_�ɇ6Ne2��?��,���ѦAY�JIF�8�L�^߰�!���+эk���U�f[��EX�s�d�~��3����J���%�k���?�J�:Y0���*>���Д).*Q�ʲ�.�k�>�F�uD�6=d�,����ȯ��*���+cISh�:WE���☧'�>��m���rl�D�s���_4u�j�Ój���NJ#QPZAn��~nB�_$�����㍭�+���Q��}R��f�k��6F�����TB���b���]��q2h���L���j4-6K!�Im���nm4'O��{��?"��{E���q`&����6�j�H���0U����jԝ-�=�z�q�	5�-��]���ڛ��ˠY]�+�>���x��}���J9Oj�!�� 4|LE/����/P��� �s!��3$��>��������dҔrk��
z�s�kT`�#�T�l����psN#��^��+-d�7� <��Y�&f���=�ĩ������<+�&��07%j�2������T^����o-�(=��Ж!<�� �SV]��wA�f��Es�in�S���j�{?'��z+o���s����L�Z�γgz,�A��|A�����2l���%�ݽ�dw��F_��a���6N���h�"���*��n�}��y��֘bـ���4�<��a� �F���$[�WP@�Q(y�.J���<~\6���|i��㳀�c2:�
�krx�ߞ�����}3Rq0�x��\����6j���� �xLZ����ik����>�N��d�6��) �TN���ސ��5��vI#��t^��y�Y�xs�b�{��V��B�i8���~�"���Zq����%C9�{��������6p�/T��!�yN��� �ݹl��m�Oa���;@��+[��h��2�)�"�.<Ԏ7d�v����>�ǚ�u�6�*;~)����6߷��s��ӵeX��q T6��F}�Jbe?1[���ؖ��t
���~J)�&-9���H�C���$}��� �v "?��hλ*�&v\7y�h�]tE�͓*9R�����4Dݒt�E�H���C�ԆC��OM]�p�U��� �G/@NB�6�U�Y�I& ���y!o��qMɁs������/�_s�NfAw_@��9�H��ڷ�D3��H�,m�̤�N��t���^�����X�F�XN u?xkf]��+9����ҋ��]�A����r�>�K�.���m�������m��8��i���O����F�<�>��"�jt-�t��>d/�ӘtsK�N;UQ�PR���,j�],���*Ɵ����]GV
�d����u�V`Ԝ]��`�v��R9��h@�qH��/տ=@k#+";�P�ō6m�(o������ �Y5zP��}cUrb����@$�#7b�:u��'���p;N��4Eƃ��B�U����G�@�6!�j�����ɏ<��]ԙAЍ�������/&5s*?.�����!yə:26	'R�F�����PP1ށڍ�� �GܣxZ�kя2�r)�T��,]N���RJ���SŹ�k�2K���%�>���M��U[�0]}:�i��{]�ޫ��`��>�Lu`>����^Q^������O���AUE&V\��T�����\
q|JdS�"@�������`���m��a��K"�0�:P��Gy��+I
He��q�HF��g��KDv|D�J�t��E��.�:}G�X��v�D�+�Ԇ�Ϋ�
��C3��(j$8���5��u_��p��G�\�l����ke cڀf�7��5����0)R�+��-�������P�Z�?�#�^��ȡ���k&����a����~F�I�p��CX��a��bL<�����8����\�B���)K݉�,��<C����-����\� �2�������X��[��/*���<�N񴮈�VF)$f�IUG��lF�;/օ���}R�N���PcE�Р����
�p������:�9��+')N��7�#f�Բ)���C&+zJ�/KkIJ��椧?�V��0�Q�ZŮH������q����Uz�o�%j���Ǫn.3�a�i�~8���Y��dR��!:�ԗ�nh�,V�d��|��D�9'c~.��t���78���ձ�l?"6y�����&d�Mǉ�9�V�	z;eU�.s�0~
��@7s'���TL;��`�r��j�N;"�*`c4��:`�~SH��:8F'	�aVe��;*�8<!�d�(���x.������	�G.[Kjt��������mvb����� ��o���(+���а�?qx/�ƫ�I�Wr��|y��E��x[��^A�ђ�V��!3����;8��q�2��hNb=�|���~�Ý�̰�z�* &������8A6�N���ϖq76&��`�=�o ��O��ބ;+睐cɑ���j�}s��Y�sl�ڛ�n_��ʭ����ZE`4�U)���s 4���i���W�U)��� a�@%��²�ƇC6�軗O��lH��0=�H�0�Al��g�0h��V���6uB��I�Ӎ��ݍMC�m�M@�����g*[����7+[f���x;�_!��nE@☒�1�~H���؊�Wm���p���V)��e��t��=&~���l"�ۈ��UݬG
�=]��)��j�c�۟�Ά®7+3�BmbE�ћ��V���N�J�A��o.����©p;y�q�p3a�{�x���@�!W���:���o�o���/ů���o<N�$g���(V!_єp�fc��^[:ͽ�BcCIqy�����5z�8�����j��c��"�ӏw��.k�9�1U�hu�>7[�H����j$UV$j�,�]t-W��]���d��$�(�*���]4�X�8�g�9;�1pI�Ѵz&!�^�ڼhF���X4g}G,N�y��$���x/[�1O�������6~�k	�Yq.�x�
���<�9e�$W���+�H��i� ԍ)��:���w�E�q`8h�)�y[��`v�L��U�;�X���D{�a�Oo��~G�q/�!���lOS{��x;(�
Q"��k�xq5�Y螚
��r|J�]Ꮝy�M֨����'�+f �]VvH�,
w�^��}6Zj�?�iq�M�A{�i.jނ��O⢹�^�5�JEfK_"
��?�	�TFm�t)^��y-P�`��I%�fg���L�E�}��5���
#;4�l�^%˃��o��~:�hF�]tK��oZ&*���&_���D�p<����8
L�I�],�2D;�h %���=i�#F���9^Z�^����7��]� �-U'���P]`v�&��-����7}�a	p'�i�WҒik00n]��/Tb̒�Y���F�Aޫ>61!񒒀�4�Z�[�u$P}I��9���8B>�$/��Җ�]�'���|�d�2�2�̐E�D��I_�Nj0�;tG�..V�ll5r�{��Y3��	"V�}$ob�p��H%Rx���pE�.��Dؑ���E<�׵Q)�A�ҕ�9g?t�wA���/�>��5�����E�HD[�I�;'l�|r���S�s<�4��ˊ=��љ��]K|�WY�)�JN40��c������&3�"^��zbK7!N������QG+���ozͼ����8��˾��Z���8[�kU�C��B�e��TL;�ׂ}����d����<m��)�s�x��q�g���\y���~���8L��6`�UɬH��Ŭ��~��٭o�?R-�4VǠ�"�g�C��?(>Pðp9eG���s��T�A;l�=��Sb�[���J���1���h�tGPE�(q�W��Y㵇d��#�;�5��~M?��6��r��H/��Bu�
����y�;a�aF�<��|\�^�>��z������g����UkN���_c��<��	��9q2�>��`��'��jue�״9!iKiߥ�w������/�*	��	��+�&�xm�Dt��Q-w5h�FT9�K���&��D(%+���? 5>�P��͏��N�;��p�2�YCh���7�A�.�v�RX�)��?&�`J�̝�*o��xF��&�zon:w�Rd]�,��H��#(�qd�6ÿ��|�a�x �:���/��k�2z�Cn��YFVgى��*Fe�s6�t��s��IH_[x�i�q�phk�K��%a�wB5K(K�cP��.����-2��A�MN��~i�Z��?2��uPN q�Us!Egq������GW��p.��5�IAC��䥌��h��C�d�Xu��sɅ�]'�q�;��[�B�G��c���K8�����*�|k��n/�\"��."�i<z�D��l��.���<�.��>|��S1Ԭ�������8$a)"B�> ����QG�m�ʔ,8��ݐU���O��簸�:T;��q���^�{-\�Oft���o����{jog��ݬS �Dz�m�&�ێd[%��r��g��B.Gt�Ӗ��`A�w�J��΀�]OD��z���#�s��n�/&�E�����qd�œ�z=���=vn������i��v~&��d�Xg^������rE��Կ���
�:��|�0��R��F�X�̭����;6لOS��!Q�Qr���k!)�!����k�`�Gy�MWl=7�x��l�e�鈒bl/B(!��g���Vŋ'�OL�i$\m_�NJ�A!4�`n�
�vO��>c��_~�^�>�`�)�n�i�]4��*���J0�1Fόj? X�;Ǣ0�s�#5�B����)��)7j�[�LK�y��<�����K  �N������V�M.�k�/��L�gQ��!�n���R\��������\?��|�Q��|��Z 6&�,M����3�ˆ�J�Vw����<c����Wf��ʏHh&3+���VQ�Hߣ�8���]t���=�_z~I�Ώ}n�1	P"UA#��t�yv�ıc2�����9���N�5�uP,�z"b��Y*96!iY@��
�g�w��,$��QC]O}���1��Tgj_t(7���@^�
�%��c �$��_&Yp�� ��i܀�ȿ�$z맅6��(#��WzH��M�d3\�����ˏ�P���ep��F%Q�r�ƌ���9�X���<���1���.v*�,�o7З��Y��~k�VuÆ�WwY���Lx��J~�:Jm��G�F����S���ǤY����Lim&��L��ڱ�G��2M�*�6�L�͍d T���}�>%��C9��ө�A=�g�|�%�l��:�{kPnp�݈Au;:��(�e����"tbm0h1�F
��m� �-�~`���hx>����;����ڴ�@�b.�����{ў2�d�
�����0*Z���ְ�v[��N�+9�T���6o[Y�S�@�*|�'QGS�~>�����������N,�9�Z&����a<e&��*�˶a�����E`����{�C��)h��q��0Z�^��%d?�V��Zt��J^��x����@���݃�X��ZT?�'8���M����s
isq��OxꆙĿ����kZL�5	�PJ=��pA��I���
3RW�&l�� �9��n�{Đcn��ښa>D�T����������ݫOj�uߕ��dcYE�<��T�A
��������:�(-D�tZ�i�"����"-���0�����u��Y@��x����.k�`E�լ���(�bȜgm?������U�|��60a$Sk�u37F^k��M��������)�2zb��0�܄��q�zE9�p)�_m��n��D�mZ�[<��'%o�)�I�0���Vp��Br�2X��B��i�VWJVZ�z��Q `���Ͱ\�е�\r��=9�&¬��_��%S^ر]���C��/��p�Ce��ym�1{��V��� ����-�D'�	5�s��}��Fe��t�C%u!��]'Y56�`�N�v�"^
:�^2Y"�F<�C���,�^�N!����tI;�=�}�j�:�t���=�9I�By`���yk�v37q��(��Q	�E����r�[�7�yQå�@)�8���M������3���1�c)r%9���
즻�
v�H)�]����;9��(&}ů�F�[�>����6��D�@��>�f�$��x�w����Z���W��*#��1}�� EC5h"sy%�5���|������s���@����e�
��ή�|�,w�|� -����_g;�aB뽧!Q����f�(`	��߱�Q�9e��w�t��}�+��{�W6�?BN(l�ێu�:P��L�ƛ]Ү{�D�� �5j��b���QHf�m��� {G����FN9�"��:j�|2�`�'�c�|N
R"�)ҾD��ٓ�bt*j#�%�:̗�%HQ��սi>�)H��WM[�J� �m��S�	`��P;)�<�+3X����hj�v#$�[;�oúސr)�#�w8�	d���b��蟇f-vL�>!&��{�zO?�����܀8�O�B!B<���r��D딼*���A��`"�Q�qJY�#I%.��wn"H�h>=I��L�����f�$D~��U���ܷ�M8���6*|�F�PX-HVH�ӥ�R&+)I�-zg2��5��a��#G � m"���t�F8�A��_~���N��x�r{�{��]~�`H(̒.>�(j���V�{2�hz�uRs�<F��?������խ�(2�.煴�����1N��B*~f�rݚ]��ï���FR���P��_��e�7�\�5)�1�ItK�a�a}�;�ߗ(v�T�ɶZ	�����ΐ�D�g�9�qd3WQ'�(���uc��{�ό��,W�HϤ�y��1��ղ<����*G-�A'�@��95vĨi��Cj7�Sk�`pl�r@`��P8k���:M^�#�7�\<95�!�/��a���#NvV��!���P��<�!&x���mO���W�D�OA�(�D4L�kN��{TU��X�P�ų���z���c�j(��# eԏ˧x�\�:)z�����?@<n(�$�p�(/�AJP�z�k8�,�����ғg�S��<�mϞw.491���X�����A)_Z��h/��ЅwQ��`i�]i۵T�ɜ,[B�r}�i��&ȳƦ�<j���������u����ـ�1$5,���!<��.��c<��J1� ��J�g�o#�����P6��}�5��tI� �q�
E��sb��g����S�$�w�_E�V������g���9�=�{�+��;��ZQ	��M����9�t ��FԲ}J���lwr�]Wl���|S�
�M��n���&��8�P��D](i��C���5Hٿqw������!F�o"J'��8��؃@� )�B�����)��un��΋�Q?��.��4��I���L�������FT�V}������K+��&S�\-?���+bjXcӶ=K(�:�V��+`;�:�<��0f Bs�GT����9�*.��a�f�{>ܐ(]�a2�,�ېxr�mY���}�g+TK�P�Yz1�9D\!l �9#e2�H54��O��ߝ�'�o�F�8F��]�����3.>c��q��l`���4\%k ]��^�����2�C�TE.�x��lq⌋���0����O)�(��.+Z�̸;wl�04�5@^��X/$T���k!�;D��fmJH]#&�󙔆��!�՘�s�5
���)_��S����h����fa�]8z�-��Z����%��!��6���a��oY֛�Ŭ(��_����Eׅ��&����_�Iv����NA����i
���T���Of-7bh2�z�{|B,�h�&"
T,������̖��(~$�j��d+"JaN�/q�r^X�&Ƹ�����@���2�OR��n��{��bָ�^7)�.u)��4%B��#� ����~(=�Ϧ����a�(�O��5t��x'_}�b��*	��U/ưq%)�&g���|���Ң���r��U�pg��9��Ȧ�8�X����݊�\kA����_������bC�'&��
"��Pzy�����<�t�Y"�f�z���x�5��V�@Mk<H�%�4m
5򇮄q���Z�	���ڣ����c�׳��L�����grZ��[�1r6̴�1-�)�%��3IZg�o�V���mN�d�*\Ò+kvQ�1�h��J�ZrO��R<���!����A�받�d.�~,#�(��h
��M��^@º(����G(F��[�>�0�j��^%0�c��8Գr|����O9�~)p��IǇX��Y v��hHK���V�%Q(��ڞ��ԅ��oS�M��:J�5aD�Oq/�E��+	��:���.+�f��JĮ�'��T��/�	�波8���DX�I�j}ګ�#��K�i=��<�"�:sH��a���2_��S!�{y�LIu˺%��P �;X@�D� �W�܁I��҇�8��0�7S����P��TM����1G���k'��&��r=rAD�ĻhC�T+A|?�F[�%�,�����I6�MxM�"�o�C����ܥ��<����9&�����Fv*X�ƨ�(���ε.'���w{�Z!C��m��Y�=&+G���ħ��du3�H���؛8��1N��G8��j��P���b〯Ulvֈ!?��'!���q�u2[�+Q!:
{'$��t�3��񨯿M���̷(	�!Yj�-�֔���ˀ �E~��f]�㴬u���������:���&�~f�~;���6~]m7��Yp�W�����_Q3ʫErR��nבK�t�}��$S����8!R�m��5�M�蝃�w[~�-Ƽwej!H���|�l%�qFP���ق��ɻR���羲&]�2i��2���]��3�ԟ���\b|���bq����j�5��m�z�is�&��� /����O[���������&��N�a�u��[etj���Q/]^΀������7K/;˵��b=2R���&̖��� ��;Յc%�o[N�F�4d{u�[0ױ�<~��E�#��	�J� 3Fl1�� ���xT$9�+W^�}.6�����)�6�0�**�����<<���+�Ĕv�L7=��j8�SYߕ}$Y�_�C;�(�҂w��-�����֢(�e�@�*�0V�aCU�շbx[�Z&�Ӊ�~�3B4HX�a^�9:�W8䃵�~��2lkHY�5�)���*}�O��{��g�P^8?
%��s1��z)�(�,R�C��`� �k	���B�TJaq���Z2�d�[�&*�.�����fPӌR��џ�x����7�ؠy�B�Q�0;$�i
�=c4h�߇��2������h�(��^*�#�#C��ȹC*O�+����D��s#I|�N\�Ti�k�a���u/��xh��$w��U�ʨygw�;S��f"NS�U�̵�!r�x���$_J����ew�d���(j�tk�S;u �󶯾�[v)�v�ʣ 3�����7
�AL�a�P��;�Xr($��w���[7�)9����kx��Zp5���x�p^��Ĺ!p�t}�6�(xf��u���6�s��≤���.�p
�. ,�H7J�˟	��6h[�7st�)zw�S��a��\{d�;Eӡ"�B=���P��|
��?�y1�� ��(�O.��������~uC,R��j���*
�3��I{+qN�?�AT��?d��q���so�z6�lz��5[�U�"��a{���}R�)F�4�Ȏp�������q�âԬ�L�����{��@T#V+c7�:Q���*�j� �i��+�s�J��� ��]�6q�=��aA,~���ȳ�-M��WU�S��q��.�C3��}-��v�F��pa�j���x��jA,G��=�}�h Ъ|(�󤃸�f�R�������
W���Q�� �4�Kg���8��d�t2)�? �Ƴ����`g��� �3��vdd-�m�O2������,o:�K�4nP�Ӕ���>/a�RF�!��� 5�y��o�wL�8 Z��p�Jc���P8K� [?45�ak4d(I�P糧3ob��kU�c��h���ѝ����2kzuK�t2�u�p!'�����~VV�k$k�E����]��-�-��xs*�0k�]�Bs���w	KN�B�%��0x�T.�G�߀^Ty�&sP@��dE~tpY�氬9�릋�?�D���slɥN�}�����E>��x�S�8e)?���'��v�B{Ģ1`l��*�����C�\۩Ż�^�Q�'J+��QΩ���X�"U��W�ٛ�؝�0Ob�p<�le��)�%U���|W�w�K�p�f����P�y��0{0]&nvqE��Mju�kδ}A�6q\�h����1�n)F�i/j{��!�{��.Md/�%C�����'9�(,g� ���B�[��n��:�>O�c L��aڸ�X���^kx�����yw�F�DO���5����;�ѣ6�0�G �j�	��}��*Z����\>z������nNU�W13���
M �V�\pKY��7X� ��d�m�$���wn�� "[J�: �$���R���N�D,R��W0�:ɕ(��6�PE�/���P������u����v�m��Eu���hQ8�l1`0���Gz�Դ���c�ߔ�IaS<;�f钇��D�������i��cR��� D���h�C�8V�j��/�S���!R�Y�2ܩ	r�4fϓfæJk� 1N[��W.~ڨ��M�L
�n��m�r-6�=y��\ ��s_�:�%���3�Q:�9^��P���K�O��;��pa>+k��ʋ�3/�C��2(x�80ӛ�!ØÛ������������$���r�� �ǟ���M�&�zD�B��V�>��/GO����P?f�:,r�m����"�X�yK�lFd�B�3]������J���H�.͏
l�y��m��q�% tUaB%�׼��ۢ?I���|mOX�����-�J޷A��'����D9j���v���	@�ŚC�&ڐ��|qEd*�ÿ����-��Ġ顴�Y���WjT;`�P"�ܠ��)<��Y
��qIG���T��Wr�2���Z5���)n�.e3'I,t�0 ~�8voݳ�М1��^1����5��OrW�S�
}�\ϣ"e��𴡄��e,���m�$����|}�yv��xj����1ń��H*��Q�'��`?��8��b���w�?�V~�-]�8b����1�v��0��&���c��Hc�޾Z]�f��Iv�����^��r�}���u
gx-� �����,�ӯ���'����_��W#���I� H��o	}� -��ݠ#�S��z-w�)�
=㌛�cpU�s���Pa�E��)�2t�3��ӧ��LG��9<�+Y$k��0�g�I*�M�d�YW�}��EgJ󢀺oi�2J+m��b?�ޕ�t,k�b��?Oe&��Z�wq"}G���Uǉ���n,����m(�v�o����;[-@1iB�%C)5��6#r{	�)Dm�2��'W��N#�u
 ڏ�s�=���� �m�/xF����i��vƜ���f���q"N�A&��aH��I��yn�0�v)O�N��2*�Lf�'��J��.2�_<�s�ОXOZ��sd���9���ȶ��RhfX�%X��.5Mu����ߓ(����5
ɔX�0�� �j���J��f�Ƈ�.��*֐k�#���֏
�� 5�����=?��ÇX"�d�[���Mţz��by�c�VR��"A��M������*��ў0$��rǧ��O&���>�Cq�����/�S���fZp���H9������ʶk�ç*�N,/f�փ9e�Or-��1�'Y)��p�H�xW L�3�U�j���p?U$A�J|���Ht�Ŷ���j6T�}A׺o�\Ww/�hYr5������7-$��U1ƴ(��R�X�n�H.k�c�D
�/�Xr��h���'.�lF��e��r܂���e�3Lt�u���!�ya�C)�Y�#��H_���X2���guo�����$:�>e{�FY���9�u�p�[�m�t�:3@�a)��VP3�`)���
���w���d��;�dM��\�7'��J`66ñ��	�L�"��ϳ�(�vp>���:�U��KLM�ek��6�Cך�PG#�o=�e�2���vRoqz��鲬A)9�~�cs*؇�����y�_+�ԻClnʥҰ�9J��v�
��w�hK`مm���K�sa��c�@`��r�z�Ϡh��Aӛ��������w���m���C����H�z�x"�vyϼ!��60-e�m���V��ݠ�b��
�#�q0�)�w���h�:[凖������!��l	���˭�R�-9�h������\Ky����8���%�i�	��\_|;�=���za!rW)|{P����|���v'���^��sc2	����U��cxX�n�a�зZ�佚Q������w��&8�8!P
�dQ�[���@���Z�J��#v�-��o�gh�3;k�dI)��Đ}�=��$2���7�`U*�C"���((v2��Ot��|��y�"~����S�߿����R��>dV{�5�� �][FK߆2�)�{��c�AP��&��;�}w
�s�u���;<�x�0zcz�w9�R�%�um��?Cȏ�Rv�Q)�G�N�M=JB�׹�!��-E:W��KZ�Al�����$B��|+L͜]K�Nqx.a�eZI�$f�u0d���3�KT}��$��p\�A �DHPY>�]Io�P�Z���ԉ��>�/�g��Q5�䧼K`��J��H\��fD�|�N,|�2{��:k\���
7�ٮ��'�$��d�?�y����99ZR��_��t�Gv69l��MƏ�7K`��X�B$��$�����i�	M��bE����s:.b/̫���U�̃Ba �C�լ���Bd�IX5��q����\�m�Q�D�Vf���-�
w&"}�{B��)�������屌k��^ٮ���׭H@El+�~��d�w�:0H퇑g������qF��PcU��F2	�eڃx,?�۞ �u�"���-��A�,���Z(KE�q���"s�i%󇔕�Y�h��Ly�ݱ0�-X�*�x"b���5^)��IϞ�^bs�kU�6x�ph��U���H���qEU�������0ۦ��ޢ�(�/�ASX>�۩��a9*��7Yk=\�=�CL �V~�@�Qy��˨
9�s���Je+�����\W��;`T6�����G`�qzʄ89R������I��S&��ςK�wiփ�7ԪfL��H� t��'�c�
�C�"ij���N�g���s0\��d�X_+X��'��b$����y��2;b��m��M������3i-��I����?�NӃ�)��]���`;���W�nv�/����Ԅ`�p
�Ο(�<�Ȉ�>N���?gF�-L+OcS9�������ĠI���@6g*�Ʒ1n�S��������U!�*׃=���`Ⱥn����<�9qd��Bװ��5�������$�|�<rv��}'Y��l>�γD���+3ԫ�&��W{@Aw�?���W�Y9jޖ�<&I8i�Jk�#{S�*�
[�Ɓ�DR�p=�\�Y���e\�H�^fn��l����L�*��}�������B_t�.V�����-�E~���C��*?{��$ڇ�ml�4�P5v�|T	̐;8�]N ,|�9fi�����	���~�����w��`^�ҩ�}�0���@
4�-0�&�'�ȴ!߫;*FL���
���M�	w|����t�CB���,�p���
l��2����ٌ�C��@]���RY�]|:�Z�t�1�sp�X�g>%��Ǝھ��,���@�6XM�����Wcq���g�a���P؛Ļu�i���˥�/��2 ��DţW?�(?--G��v��l!�i��c!=H6�FSN��C�u7W���Y3�I��k�H �7�3�̷d�<v�`X;<��q1}�𐹘�5G*�*��Y�p/�����3��'e�Uy�U��V|(��Qu8�0���CV�H�/��$�p��C3��D�#�5IS*�=N��yߡ��S'";�cp�~x��MqZ\0W���i.�׃��V3H�ܩ��%�&�4��n<e�V�Xནw�\�A$~��\�`�˥+ǹ�y�0�O�0u<������4I�&��\�%�����zt-�2�N�X/P�2>8�i{�sCrI�+4\k`k����t|�s�q��F/i�3�Ȥ��>D���6�h��U���s8�P�0�H��r����䂏� �χ��5�����m)�|gs*+"��;�ߓ6��w怪���aQ#ж,�O�a���\%��h���e~�A;e2��i}j���CG:I!ns=/ޒD�� �	㟠���Ԩf/U�SO�nQ������-2�a
�u]>�tO�D���l?���rv�^ױ���0�1����d�md,#�#�nY��`)Z-��F�V�x���D��Xu%��7����Q�}'��xPi��G��7Y��7�X�By�'��.�DYyXt�>J!�u|w��Uj��sr�(4��{���b"3y�**�ہ/���ψ|�A?*@Ύ�	k5Ұl����3��,/�D!�R1������u����jaf/	DӈvH�^mU��l~���v����XR|�G �f�C��wXR��c0Y�$�.�R��W��Q�ۭۢU�S���h�E<�mmDw���(;�}���k5������;i:��G���4L�^5g��bcZ����ftecb��Z=?�x�EfZ0r�#_� ��<�z��^&1�ڭ������0�p��E�G���
��|�NJ�ƑB����Z����M��^�H�r��tϰ�(��îے�IK��>�.L�W�Bd`���O��6����?�� �m�t�����u����Y�����\�Mx���L���u������x�2dïL��c�v����<��T �F%�� �2���/� ���ػ�B̌�Sj��|A.�4����u1�c��W�.�aK�ԍP�uU����T�zQޗS*�1�h�8�a\��=�bDV�غ�91 t?/ذ�<�ZN��`طh���)�@"Ud@f�\QR�۪Pq�L&s��N¶�#7���4.n�b�D�s�9k�Ү)��9r{L��u��^���H�Q�JKM�s"�n]��ʐ8-���O4|IS�o1�`��+%@���;j����f�:����W�+�o�Z��V8��nlViBP�pds*h��=G^�@4t�]L������iqiP����V0wz�Y7O��e�H�.���G㈒���0��_�9�e�Ib9��(~��K�d4#Y q9J�������8�X�&yҺ*b��W�'���I
�ւ����H�?Cs8/�c�꺞�M���e��m�P��>��aqXk�c��y��\ܘ�a�\8^��8O����#Y�R*^z�E<�N�"�.�I##���#����*� �\���M���
��v6в\s3N�q�euVjN ��������M��mt���	� �X�K���i�L��ӱ��T�?r"���<����(���\��9y���"���i����m6d�%�W��;92t���g��4�0�G��^O�8|N6K 6[*���
�JO0񜼒��o�`���TY#(o"���H�{V�Ԅ<#H:�u?��U����1�O�A��J��⏁�q
�����?k�#Wl 3:�Mq�Č��^W~u���Ƈ��(����Yp�#Y�QW����՜n�.P���T�*�W��׹a�mbH�Gڂ��w����wxSn�f��1VO��/�ͺ��@�7������9�/�B8rH͖x��.G׷�TG^� ]���G��|1��/�fDA��HF\�	�tK�D��!�i�i�Q7]��J(ϡ��<�S�)l���`c��}��S��޷29���(�����������3����MoYH׉����]�C�}5�Rq��Sg2�x8�ik�&W�s^�0��2iU��2.��<>9Of1y�W�RǸ�:"��H�U��<�d�n�k����m���'"�?�=��1�\\�K��0%��J�	��0aI�f7��HK���@� �F�N�	ZĀ%5����,�6.��΢7&VK�sg�R���L���^C���ܳ��������u��a~AO�fp��A�/vf�AA�m]Ɉ�U'�q��l�:z2�F���3�X�B���\*	u�-�nj2���!��Vp�Wo�t\^�֪NR�F������T�=��S5%n�u��q�����͍���v�M�R��,c�	�Z�k[n��,������l��`��N�#���~�F��6��Aa��
w��XW�����oEg]��;z���	�|�y�=cٛ�3�^iDuo��?9d���-C�ַ�0�ӂ�����8ẓ�9NW>w����ؿ�d�6U�w^Jt��^�� ހX#h��PY/������&-8~sr�j��t�1���7�DC���؊��/�uWj�I�襩?������n��^���xi�m��&��!�/*�;�ɿ��vs���_��d���Ws&ư����a4ρD��^G�|vA�T5��uB�����Ot̓����ʌ�*4�-�-+~��7��hfL�&^˔l�~Xx7����?M���3Ĕ�;�N_E�EC8���q�ֲ� �hkt�uW%v24�:V�f���}��Hz��
CԊ�c�v#;b�%��0��>�geN�*�7=��ٺ�-p.-4��h(;^S����(���m(�P�+�<�#`;�@��2gz�nĴy㕢J�<L^rZ?,�C�d�B/z���(=�q�iԴ�.��Kc��DԴ��|��F���ᔉm�!���/�n�ex�hΈD"�8&���� {ɚ��2"{r�~P��ḭV�����_@!�%;�eY���:�e�ғ���Y(t�/V��>��0&�]�}Σ��.������Oa����lߏk��i^��iT��hx\��ԙO��A��q8�<�:�{4�V��7 �%�/ӺfM��{� x)#����&�B��4�a�6⻇{�w��<hX���+bL4no�K��k��{���ߡ4�$]��܈�\EZ7�� ���j��߽'41�I�1�MK�-����H�(�p���k��)�;���&N,^���Hw��R�z<���}t=4��u�H,�C.��=A���8�_��>�_H�b�T6�h��̵̬����k!q6������~�[��;;���#��2�ht��k��qnЄg�#�4�0B�x�hO��W�[;�����@�/����}�xC'�[�R�}�!deS�1 5D��\�N��Nߔ���8����c8 ���6���Ru�?��Mı?|8�K:�S��?|S�@񊯔K����6k�
��������|��4����e1�׎�RL�͚�	�:�
]v�=$��b�۬~������0_;�ɀ��UȧĶW�d�P��v����v9�#1`�,.�`�S���n�,B&.�D|��;Ծ��-����[l���x�dC��o�PH��*ZUh��xTߜ�6�8��/����x�8o�wZT�L<޲ވ��F u�XU�}�\���$$ϚC����	��W��T����Ei�	�Q:Q�>��'s7.�ԯb��kB�
|#a���~���`�ʢU�!�n�,�Jg�8O��ي%��wj(7��E^w���^�EuI l�_�&�q��������lzo��@2o ��[U�[E,��mK^!��U���ц+m�i=��H��"��s��G̵�2��S�'���E+�^�V7��}Դ9,Dg��枸�4�X�T����É����hZ�I����L��)�J��y%d��6"K{��z4��5i6�m�{5�=�K�Z�_)����%�	x%�"J�&zIt�b
��r��ߥl�Ӌ�����ۄ#�ӕR��0��S_Y�!��9s+�Q����E��WEC������[b����VaOwXEɩk��5^�	G!��P���E8\����W�#��u?�-�
�[�g���$k�A�Ϳ��nb�!Վ�l]��+�������8��,^w�_���r&����4K�-ﭺ�Ji�L_O���qb
*#�D�]o��?$H����t�Lr@W�;F@�X���&T���gJr���LM%(i6E�[�W�c�5�Mh��j?H�}x:��#���Z�#鰎[�M��Me��{
@�w��	���d���2��+hv9��l{2m9���P4��N^z;��h^ �[�߽���LW:��a��7.j���pE,��^d�L6�K{5^[,�_X��>��c��� 9�-»��Bi3�7�k"[�QB���.������M5���'�e���ަ�,kݱ�7�,�)�C�o/���i����Ӝ�i욑c��'�/h)nA�Gf���ǳ^u�r����n)4�o-2 �:�
��+_{����J��I�
�#:�ąGOB�il�>���)�>t:8�-��H��E���ܻ��|�����o"��S)�%J�՛�l>�$�,@s�;�'�Y�˅���r�)�ߜ.8����nr�T�o�bܰp&�倕�Ky�24��$n����
���y��ͱߺ��6M/}���۬�}<�_��{{6�<�^C�q����a'ܵLk�ҿ�Մ�` ��oZ�T�I1{��F�c��o���z��7֔t�5���s�̩�J�лYZ�x]�Y��3[eeZR?�T�!a�ƘA;�s��hي/�J25��Hi]ߜz�	�@�M���N����~㬥d ���LL#Ȣ@���j����1��=E��Ӧƃ�K�I������1��"�A��X�;[�z�M��
l��
�^?5��}>���-�i;�y�<�����Ǐ��W$Ʃ�����`�v�=�@iAȇq>_;��p�5~[�M�dEJ��ߖE����F�Gm` mSD�7/J)h`�`�m�uz]��щ��|P�Q�Z^����,���y���t��E�F�~�c�J����^1�+_��_�q�t�*�]�O��U��;<�o�bx����������a�d���P��Uc ��8ɨ>U��?%'���0,=*�xx�^��D(|/z��]��p�7]jv=��g�|Oj��F�:B�k�ׂEپ�/_�U����bݴ<��`�q��{$Q�w`�}i5T��7�j7T�����%�wx��;5�m�0�-%���t����Ah��B�r=ԃ7n_SB���@��`wh�F�_��ڍ6�@gu�{����KG��z������I[˷"JEbV������Y���*r2	n����}�o��BX�<J�=^�F5p�=��y�;t���
�z#��`�
�̊L��  cz�����%��çLH��|�e�Os�B2�s������z��`jX>���u���<���,	�5}y4��e�l5Mhf�Y���IH�^=( �e����^L��BX7,�{[gr ��K��RK�5BA���D��Of���)�u�g��֞��
��@>x�g�H?�%�(S�N�<hc,�N9�v��hg���ۺ
�n�dh8��f��ogfF�|�(b)�[n�*+�yT��#��K)R��H�<�YR9��üFR �Y������뛇p�l/܀ �QK����q�xh?h�B�0&�P4���!��׊�(�@��L��}����,0F�kO�x��.d���T��w����+����R�=�#�_y�ƞ�E��tpx�O���W �y!�k{W	]iR����,��XU2g�1v���%5�!uE�3˧��
�����MI(�ɀ;�໵;�Y �?w6y��w/m��8��6f�[k�G����d��3Q؃�`�u�ϮvZ�&I���.�cr�%�	-��.Km��Z�<3J���󝵀�&=gM,?��.���:�Q5'/f�F�{7� ^�o�d�l�OcD�?���_c���j����\�Rq5�5?�i!Y�]#��9f��a�>Ю�n�H��Jxq��7gN�\{�B����{lO�z�J_#������y=�U �l~��jq� ��-���M.+����,���8D�J�C��AB=�?oR�a�_(z~�'�hW��/Q���9f����]6rl�_:�~Z��I6~�EU��}�
�YY�X�X����!A�\kq�
�JG�g�q���rӋ_%�5��V�S�E�KYZ�3���1�����QHt�� ��Pa,���9�
?#�͈�zu�\ɟ�0��ɏ�7h��J�u�id4{��(u��գ裮#��'*��F�g?/�2 $X9�'���$F��l4�l�,:���yS������\��ݎJtͿ�]�JAι�4vs��;`*hԒ�JVk�
�����w߯�3���:�lLL���Q]=�6GՊ�+r�tN�w/��M����|bu�����6��ֆy�o�I	��;�4���Vz�U�d|�9�4���s���.3"���ܗ�1�A}����K{�~��,�z+<��muv�.R.��E�R:s �qߐwN9�^b�G ��s%�n*�5�M�*_]w�9�V7�u_eﻔ^bH��?�z],��1��^ E��n�2�*������c�k�1�5++�ֽ�)���kew*�5ƕeL���%A9����*�"�z�Y���0w�:�M��ͅ�d-��뱴����D@I����
E�'١1>[2Z�E� ��E4������oƲ/ɻ��(+���@}��݄�e�DOBg̮B��h�!}z+l�
X�{�2���N�5�����D;�ɿ��|���DdJ̔Ձ�ӫ^�jL�kj,U���Ua�ʟY�EDDL��Fz�o����  /<m��ȃWzr6F���=�2��v�8��<z�8�!�S
��Od4{F��d�T�#�����9�Y����C��r�:�16�g�<����/ϷS��B�T4��J�S�	���$6��!����?<���.�	rn4�i��/6����?���U�t���-�3��	�Ϻ��m^�$h�Q�`��	�gQ��sXG���2@�"PT��t���$Et�h�=�A ��Q}@I����ރ�\	]����WV�2�������:�/�%�G6�頪��&X|��|�����.��-��F�뻇��G{�.Y��O5�K��v^��~qRd�5�g�b�I'�B�&f��&!#��Y|67&bǛ��9��U:��R�v4?�"�q�x�6��t�(��G�]Ǖh�1U��8idrQ�tj��p��	I^7��n�sސ[�̳�M1�8:�I	&��H+"f�D����^�����I�-ל���o󴦏�D����F~<W���l�Q�z��j���S҆x�n͋5ۖl�B�f�-PK��q�䭽�.��U���Ibм�j�\�m��G��Gf�Ǉ�S�&B�38�tG�v��|q�O�v(V.]3�ฦ-��FC�ף�B�m�7�o�����8����њ�o��>W��f���hRd�|M��ۆ�C���΋1�k�z���x��� 8a��s���z�L.N���.�
���?8f�L��:��υ�#ƿ�N/�[�9Б���C�ֺe]!��gx�H/��=��U�v{����)U���
zi��K4f[�%M���=4!8���~c-�(-G��~ gY&�-"x��5
��ns���W��T�pB�.�L����d��5Xk�R��X����+�E��-�dT�	YR��i�M���M��a@��	4��ˬ�.���T�Bm������Y9R+kG��a���(΅U��9&���J �9q0{��P��Cq8c��?Vʰ$�?X�?�U�xsL��v�f��ު����.���f���B��IG�ҺܠD���h�ޅ�#���,��9B)��]�h��3�JȻ[�q������2���aw秛��ޮ�u�O��d���,$f�N�r�B�%�ŻZ_�;�G}V}���׺��Kp��j2���ɭ��c+�ԙ�d���<���X�y���W]�D�Z~�eF�N���_�<7�H��-��}�ߙ݇q�F��*������8���j6�/��c*����M/��j�6�������yn�h�=FK�૽����̛��G)�� O{�Zq2ܫ��A�?M��m9�r�>#���d`[�	�\�_B�8�<���FYB��mN�f�N��ܢ���z�8s��.�1�t�M��z�,�� V9�V�����p�F���؊����֮�	^�k~�l���zpbv5���ֽ�P�p+�5��ǌy046w��I��A��IdBp/n����CL9��K�v��Ή��:Eo�[�V�Ek�%@O����K�g�;W3�K7�\'39�Rj^;>�fc}T��,�R�㋿��Uw���FCrk�h�a��\�ϼ۔j�d1��o�=:'	�@p�T����'�1t�'�/������I��N�o����q+yd��H s):$Ȃ�v��d-U	��%��u\��ik3�F��v�t�D-@Ϋ���L��fk������1����X6ó11����,N��_bZ��@o�+�`�氐œ����3깄��\G�UoR�P��R-0�8jFG�&Y�<������p|M���R��_Ti&��W���)�s2�Z��M��@�3�A\��v�M��0���r��(w*u���]	�N���a�ю��h�9=.�d\T���f�:��v������& ��(Y�}���vLj}��kʦ�'�=����'��Ύ�5�P�O|�ؿ#b�� FH́W��	���UwA��c�[�nU��3�t���6jw�y�2^��y>i�M�m�:l4��gf{�@�S�{�n���u�k�)*����'�TzP�m���X-��1���C ���UN�P��v�S��X���9j����-q⢶������92E7��y㌠��g��Jj�g���4��@��K�4�����R�[��I�m�A<�I�krR�w�x�^�D�x�!9kU�k�ۑ$^�%Tk�����G��N��ufipҔy8�OՇfejo��tQ qr��`�z�%�㢸�{߾�G���?�2�lR&�v~\��b)���7?���$�ځ�g,U���$nn�j�'��|FQ�����	a�>GF���h�К��BG���%��<�'�?}k⤟9���e޸�ܕlg�s_��T��E��	6A��9��I��ɯ/��*�^�������ƪ �(��ˀ���Q4���%�cӸhT�tu��Sm=R�Z�b�諜�8�G/
��Ӻb5��QքU��>�[���*���J�0$x1'��"O�O�����a���\n��a(�JV���3Y`�	<� 9J����yeP���9:��X�V��HUԁ��9H�����$'�!�״Cu���H���4(�'���I��C��i;��q���%u�:Q #g3��+�3���ƞ�B�,Jm���L������@�q�rI�٠�о�p+��ڠ�K��f����s���
�lc2#�*�&٘�x�&������SX�u��}��U4����F�8`�U8@��ZƋNǜ>�jo_�j<��wۯ��`�´�@6R̓԰F+��x#�d]��<^<��*�KV���a���w��m�l�_��eG1*�׿~�g��=����|��q�fm5�L*�$��ilӑjWwĳQ��LH���Pz��Mg�C���q'a��5j�'MЕgO�d�d��P#tį���,�z�(T.Da�xQ��$�!�a��3(.����b$���!1o��G�nT:�&���Sk�;0o���q;�=G=p���Pf�TeD����ɿH���:�㠓^��@ 0PED;e���
= ұ�|�)Lnz�1�9���a���t?
��\aD�?j-�G���i�"b��7^����Ku�j�<���U���z���X�Q{�j�u(�y_�nT��qT��n�}X)ʪ�����"og]N��f�I�%�P3[��w�+U���Byl77)�/[��Ɏ���������� ���z�ԛ�&�c�f�Զ�'��ֵV&�H��J�h.��xU�+�J�
%����L�-Oq[���L$m��!U}��(�@���#�_/y��wR�_��י}�ؾޙ/��L��0ؖa�-%Y�u���9��ue 'MMJ���(��&hB�٩��!���<m�9��T��2�����,��hd�X$�#nYY_�:'Q���:�V�ߚ���E�d2���NZ���h5�w�LrO�y����(�kR��c���,�Bk�X��)i���&a��d��ON���t5�7�F��L�Yg�����=�v^
ӧ�㽏��_%.�3����'	r�k��j�M~���t
f��wJ=�ū���
� �%�+��[н��<��ٽ���� ny�F�NE�`�����;�i�N�A�h����FL�>�{L�S�w"��Ӛ,�뭋*�mi](č^O:�3�;Ŵ�]c/���~y��u߇P \�B����H]TZ1#y9��E	8d�M�#�m	&��R�[>i���bxwU���a������t�%��`�D�n�R�'���FaؘN��xP�ʂ��w�h�œ=�{�����$�G_�xZ�=7]Һ3���$�+2���֨���|#)^��q`X'B)�u�4i�,�J����_��A!��(p�"?��<=^Rطv�#���!Fɾra�+���p%O�m甿z��	���TP��{���� �)��h���G�cj�t5���V�5{��񉷰(���A=!�+�P-}&�)wKc����.�7	�$�9���t�V5~�*kHώ�}d�˴��a���
��Y?�w/kC�ǦӴL�~�@�\+`˫찪���a�Z7�j����1�kD�b
)pw�.d�_��k�Xsk}�Fō���c��}�������F�`��D[_?�XW����X�`�7��O��Ӈ4 á�-!��} J�b���9r��\gG���םQP��2��H����p��� �O�f���L�k��R,*��h����u�������)&��rLb���ˎ��B`l5��;.2wW?J�81
9����LE�_k�q�/9{��7o)���C������pN��#�uHZROh"�ˉ�ع�0��-�Rn��f=p�6���e��l������82a�dd���m�`���A���Kb�M�y 7DC�$z7�
@`f�z*7P洢.3�;�h�3�1�����x�x�h��<�yS���ݝY��Ru�mjd�Xc��}���p���ǐj�'u�������T�"�P�X�����1_DI�*�����7���&7I1e�dT/ýC��k�C#p����K*0���tA{�s�J�|+�a������F����!�_��0��D�p����n�⌐�5fǞ�v��	vCi<iy=y!��$f(��ש^P��}��ܭ��3���;��\,y+�h�b՘8f+K�`C
����h��E�ntc̃�+r��V:�s~'~B��5��S� ]�v<Ճ�A����8nL�к��P�]��^��!3��$�N�a��c�)�ҠkjQ�׊��ޏ�z�гO���i�Ő�]�����eB���'��OS�Ɔ���g�0�%1�~�9~h��%[$s7�YFyH͢���	�w��s����W��<�o�O��'�%F�1P0 tȿ'H�<'�8�,�� �_p��<�*a��~�F.V�b�=pa�L����V��8	^B�T�pg$l
�q�c(&6C�W<�i��RWf$*�E�ګg`��0a2T�U3T����ewX�m���17+�;z��r��dƙ� ��t'Z��� ��;±>4h��Y;��^�o��V�gc�	���y��#�j������h`�ը?%�	��ց��;"+���4o�a)�5W���L�p�&����,����.�!�0�d����4�b��L���J;��R���ܳ��s��A�l˞%j��K��E�^>Q�<m�u+9&��U�%v�g��'׹)�岫M�ްZ��� _�{�4p���<!�]�`y����'�D�h�*�72�]�3t�<����JQ�j�HID�`5-)oͤ�ŵZ\�4N��yoqq��d��v�J&���w���n�v�5�ȯmA����2���г>�C7M����I��龩T;:ny�/��h�\���k4�0�	)�G9�� �#R��Y�_�~/<��S�A��0��74	�[�m�������b�o	9i�y�}��m���ݍ-`��vlȮw"5I�BH(j*mK�u�{����*�U*�XW'E��ΐ��'j�u�����1�oES�.K���f�	��;��KA�e^�)�́�y��H�.�h����p�0ooˎ���Py�� 8�E��0j�ǔo��;rF9��"RD�yƼ +c�~̼�A��>)�&�'3+��5�'l�I$`�����	i|f��A3]T�~ ��)i����Cs�L"�%��5ː��6̪J�8�lz@|/�����b��q��$���%�����_�6K�̐��y���o^�Ϸ��65m�4�<�=�T�����M���T�0�������^�|�.�Z�r띨�_��|���7H3�w�uv�s��zy��{*�ה��'�o$,��#�78!P�kRל�r��\e����:��*U��?HN��Qz[�+���c�C���¶$qg��z@'��C�x���%"<���I�ᠨz�a�1-�/�T������XFI0vЊJPOy�Y�*	�I���������\2I�$ВAXDJf�{nU������D��s����/F�O��ȭ�0r-쏜�H^Ղ���;f�������B۩NV=^��:�3e�Sx��')�6��N;�p.�Udx����[������b��<�F	�֝w2OK�Ԋ�R�.��&���;�#�{�b$�(ǟ�8�6B��~��Ug��aq����:ϒg��:	�uQn��9���#y��G���� ~���%�:aRԉḌR����th���QV�}��2���#��!8�OQ����F���a%@�o.� �w,GTQA����guH�����'�tҽ'`q��ڛ�K��Y�7Q�2�ab�G�W����+��0�o>�+x�t�bL���`��x��	8�B�B����H�%�)��*�+G�o-}zc�~����A*��2N���`�K�.�?�.�W.���N͑���։uHǫ-\��G�'.5'�� ^�L�تH,ğ�_���dyT��j��m�1�s�m$�g6��ޣ�*��"����=/-��wP���&�Z&�.a8gM�$P�%Gs��QP�NxN�Pe���fax��\%�~up̿v�E=�8(�yЍ�� %md�쭸��K����x�L��z�F�9��y�oH��v��X�O��ǜ^ͦ�q��υ�[�J-c��s{�P��!P$���~Tk���/}!����~�zXn{�t�YO��d��C��e�QeOl?��G�̟�9��y��`Yᩡ[�+�,�2���i5]k�mWe�Rb�0��/�,o�=?{��VӨ�K�Bu�C����!S<Z��)����`1��qg����`��u&���`y�C��)YU[�K���"HfT�����g �0����r�Q��,�f/�
3��vY�\�͢u����ߤ�CX��� i첣 �8*"*����4#�2l����eͰ6�KT�FjW���2�?�E��6�����X}q(e���8G.!lR��C=�V1Ck��:	ͅM����8�xч��j4�Y���?ԗ���*��
%����K�$6���D����H�f>��U���Y�"�*��դR�U�{� �Q^G`���~�>�{�m>����_uU4jp���4:f�w�wЊ;G���)F^v����!#�A������$EO�B3��j��'O�����6!nQz�� __~O�3�f <u�ե�~�7��|�W�=����?��W�'��g'�(�f3$~��2{2�È�b�gq
c 2�"���\^��D���򑽅0�N�2�li����	l�2�jg��0PJg�\��bN�(����7��
� ]��.�O���{ح��i�*��ђ�̢
!�-��UF�5�Z�H s��Vb�c�T,��_�5��YU�
��`U6�e�q�= ����=�7�`��>�t��j�9K7�[����KC���|g�W�˶ M��օr�Oǣ�XT��)�\��zjߒ�����Z�HV�w���5���%��uj��dD�;������S �2Ml�T����	��!����B�=b[XLߙ�d¸�Ү�o�;b�U�қ
F�5�@�S��-�tNmb�T[?J�dI�{��.�g�6����"�\A��4[�Yl��G�a��:��/x�\�HC�*�w�ř�+�w�7��(
1;�����4U)�hƯ��5�g�U�ߨ���3�I>�cJ��k�] H:����+l�x��*cu�����.�r��po�a"��]�tq��H>�]�q
-&�
�7�b��ͦ'��r��I�y�JP��RÉnӥf� ��"�!�ʍwi�\	|v��v�����&�4�}*C\U���� <!�6�뙂l�G2��D�Z[,� � H�JY�q'D��v���D�9���7>�I�y����;��%�2Ͼ�6�腓�����J��n�<��?�ؚ;
��BI7X5 ��A�����m/����p���癥�a��0�0�jЛ�*%,��d��<�:x-mT�8�r%�lM#����/��M��Ax&�	W�e��2T�G��)�<�����P���/����X�3��_c��vB�l�縋�VO��n����#�I�Cؓzx��d�u�����;������/�f�eyj�Uܟ3����R�B����Ua��j���B�g�ڑ1�ړ'3QG{-�ĕ�"���i�Ԣ��83�+ly��>��vȖ�6ή��p����πN8M}Xؓ��{?�"�s�Y��4�h�EI+;���P����m����$�C� �q"O+E�l����{�}��dy�C�W��m�e=p�5�#��/{���
�;��㴸C����y�$H3��[X��~(������3��wk����l��p�\̪���Uȗ�i�����J�*62�f)J����.���H�c�&{���{���4�9�:t,(�Q&I���v�_�A�y`�PB~V@�G_����;���U�U
�NT��c�,)�a�F�p�;�N&�"����P��PD�f�*�y��h2������ :�XT��5W��ٶrOI� ��e��Ҭ�nm{2I^i*~�Q��XGUG�`�z�K�Pd��9� m�R��A��(��cY�()��e�����M#���ʇ�ho�{1��L[�w]�uY��HUp^������ڲ��=��w�?�q�t쬒�2�xC�BΝ3��<�ib�νs+]F���^���ݺ�r������)�K4d��N�3W�Ɇ��|˿�l�!�bCJ<�|���ʝ�g��2��]��GU�ټl33�W	_�A3�yM�x>T�ӬƷ�����Xdmw[p�-x�~*u3�e�Yt��?1��Yp��-��ٍ)�2�lIe+|_�>�cA�������EM����
܁��#Ԑ�b���9dQ1#lm����J%�<z�������!���Ym]���߮U����6�+&��T�-��Y+�w!5Йģ�v&�t,��X�+^��
!ۅ~���z(��=�[�3;��]F��r��g4�T�!N��6Ŧ�u5�	�x��U���jW�1�H������P���a�1�g��Hp��Ґ��M
3p(������o!��Z���p
F����V^��^��Y����`ޠa-�� %W<Yi�.�OOC^쾾���=CN'D��1�Q�v��U�MgFu��J���O_���W���4��D~-�����@����g��O�nH��w󹢉�N����A��#6X�>4:k~�Fr��-�H�a�禵1�
<EL�j����^%'b��H���T�D����5�Ԏ3�[M�d/1,P�C>M��j�;��9�scԦ��!�1%�]&����	[Qz{����B_�%��ϡ��7 �
 ���c�S�s��1hF����ӱ�>�P����7�$�����Ѣ"��6�9�����\�v-+���8
a1�O��q���q����}c��/��n묠tKT�j�)6��/�����E&�R������h�G�K?���O�}��}X�d���s2>�}����p �N�����$�"r�|@Q�UK�㥩�_��Ro�T��>Dp�&MA���Nx��u��K�;�)�^,˯���~�R:%�,1]�Ӕ\뷈����ZO���c���Mr�RBtV%ܔ��cD9��Pd�ZL$\��B3R�I�Jx�َx�r
/@�j���?9Ʋ��M��6�Dx���xo8��c\g��~�T(���S�OgSs��3fD��L�-�x��K{��:�3�$.S���#�\��*%I6�������s8�h���|��<bӀ�n��f�`���y��$v��g�c@�)���/�qB�h�4};@�3��](�'V\�mypk;0[*��Ǵ hs���/��]/}e ﺸ#���X�w�qkf�{&X�fQ�S0�8Ih�B��W���1BL0�#�JuF��"i�̧��ΌF��%��~�[�5�0������ ���p�u%.���җ=��YEh<�	�{�y�_	�!NRa5���?��g�2n+X8��� �)���]�?E��A�C�� �����4���Y*SY�l�s�{ס- ��&�/U�������nV� ��`�a�U`x< ��c?��v�0����T�79���V>�s`���h���}&ύ^e�2���x�O���M�K�9�Tۈ*p~�HcT�V3Uc�QD�l�):
�5�h�M��_4|5£t�٨S�K�����z�E��;�s�LY�>������KV.�
GK�}]���n�r��\Y'�5Z��~C�(�٧k�=!��-�1��-{$
?�I5���5���ф6�Z�¨ ��L�W_��Z��� Չ��},��������8��8G�LTR>�0i4N�S|�+��^|�O!,����>A��^��S3Y�f�$�𴃋ܙ��-ǯԋ�Si��g��m6+ � �4~in�rI�����x+(L/���������3�91��M&H��.J�<3��U%v���ws��r����I��xPCP�]I���H��Q�,^��fe���Q�6�>���h��(*�
����1V�Y�B��jXgX���.$(@ɊЄ��\g@	�C.
9YJ�=b��A�4�0�@���2��߆��c\T��/�$ȋ�������1d(��收�s%w�H����'�g��P"u�DݝLp"�.J�?)�$[L�CH5��6�n�t���j�ˤȑ��M%D[�������	���إMG�m��r�oz�p=�7�p�A"J�k�T[��%�䏠��?A���A�v����|sr�k<��7��֑�6�(��b��Hi��>Qn�!v��g�e���D�ZBq<���LVoJ��Hű����lp�/��G]kb]L�T[�ʧ|⛎���������_��N?9nC�v�Q'��\8�썂�">�b.45��_��MR��,4<�nϡA��.�z����2q�:�:ː�
P�e�K?Nrا�	�*����_<�	�EF1aF��揗<��c�=|�մ�p6�E+����|@?��:KG���]�>����eꅃ��<������/)QQ�����{u��+��bf�h� �y��չ_�x]���������˨t4��N�bΟx���,�ȥ�1V���:�Iw���oT���?��š/�"4@���~o���Z��C�S6*�U� �X9������]�C�"@?�i3��ręyw��O���:6@�	W���,�ֈ< ����h���̫S>J�;TG6�89�*�u�)ye�a[��d�]���g'�����,`qq|���,-=�!B�������	*~��$���/"��&،"�j�!KIx�;�p�ڠ=GXe��g�.,�d8�����*�Vhk�>�mt��^�2�g�B�� K��(]m��:}����E�!.�L��r.�����_�*f=p����ە�V:S����sT��%��s_���]�F@���?��<�������v�/��>o,Бk^ͽ�8�5�9�}�����ɺ@��m��j7eh���c�K��VG��=���� �X5SM�"P���i"J$ ���,���>�����O��7h���T��T���<��I�V���b^����V`a���t�(v)B �����c�(w�_o&Ϯ�Gv�FU��I�`��8"�H��ڡ�(c04�티�:�HM2b�f�zsfs��ӭ�^/T�-]ںI�ioS�+�Me��],�vBy��0��6�:�y�0�r�х#�m[:����F.�v �hg@·��Ea'��5����^=Uƃ .\Di�V�pgcG����mI#��T���ӹs�(�'��YSĦ�(i���/�m�*6�#�a
�Mq84�=ԍ)Τ�O��ށK`�W�	�p��F���.�x��sNK�I��^o�BKW�Wƙ�����`� cQ2��߰�o���ERZ��\�C}\M�o���Ouҁ��ry�֢]����;wy�(��l1#� �=:6^��a�*������xd���ۜ�0����8tB�RM9@E�&�]���4�|.	����\��E�ә���R#���ٛ����P�g�S�^�sv�kiY|sD
�`B�����V1�"���}��;���7(9���/c��[�����Ź7ۃ�40|�ϸ2/ݝ���d#�0>=Էz9ƴ�ޒ�qQ�;�� ԡ�9��q��y���q< ��s�޷�Ԫ�:`rW�dG׆0��v$����@{C�b�kkI���q�v��T�"h ̵��*�gK���0��v�}�o5�K74��̃O������ɏ������d쏸 �X�2��u��ʒ�t̨�V���e�/S7�L��d�s	*�����vU��36&���G�*�TMf%� �*�ЅN�U�3Բ�[�t0�(�G�h�4�mX�Ѻ��s�٦ݰRBGqp�o��4���İ���6�U����Z���3�����@0|�����<�3Q)��K|�8�2�P�&��=g�Ij{3ۉ�,i��۩<�Z�RĜʑT���j���<�,��J=�2�����C0�e��C��QA�7�i�x8��o$�oq)��p���\{������x��e�u%�Z�ge�8u��Q�Q���)�E}k͠wk�Z���mX/ͣ�d��a8���Y��"	p��x&q\�\��������W��� �o̱�߯��k�x8�����{�%n�_~�50��ꮢ�c-ح�%B�a�+�҆�/@��3�P�T�2p}�ލ����ne��4�Cꮭ	��	��x*�_�m�N d�w�<$=x���ּ�@�&�U���MF4�v=���Q�cZ�zƭ�x4
�|V�+�RL�~���/ez���Sj���w:��G ������^h.����έ�����c��"ؑ�y����ۧY��y��Ŝ�3��)r�m6���;�U�PI�`}NL��.2AիQ��}���^�Nܞ֫�i��3a��k�NɔrK�N�p!鐀�o�I���,o1 ;0�T�f��Ǧٹ�&�[������Oj��Z���bj����ֺ�u��wӶ��qRj�d�6� ���.(���>*�����S���2+����;�P@��ڽxPic1#�P4k���tV�r���3��0�7ʻ^,�)�L��k	h��v%W���=��U�'�G������-HJե�,����M�� 
y�(0