��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\���V�fnvx��ÍG_;�ȅe�~�>���9�>��Y;�0G+��X�LPIj�'���}�����Ʌj(U�
|g��?S��S��=�_�m�_�b����?��4̕��֢"	1�W��p*tg>�Bl/�Fm{I����c���,W����!.�;e�����G�G��լ���UV�6$�:�)��v�jc�����#c&H+ k�ސ�V ��2���R�W;�}~=�-v/tH�Mq��$�/��~��[K�#�A��~Q(���U����tz4�"�N�^�փ,���"�G8�z3՜�^v�i��3�<����s2�;��G�Y�MK�e	8��&\я��"�en�v��A����h������"�sW�yG���e��� ��͜��L?!�{:�&~�)�J� �(@m��E)ٻ�g�W��������/I2����L^؋`�8��F�/Mv��bftģfA%���7Z ��!�shy9~Y�K�$�E���9ظ�]���
��>�+����5it�Xc��24���ڏ]�� g��r�%���Dѽ�V�^>DF �g��7&bM�l���!�2r�� O���j��j#�$�%��<�����}�cv���,ͿCG�٬�	�|%h�B"@��Zsꆮ�B�	�ba8�½�<�Z�˟�}�%��r���8u3�8 4|M����R����L�C�>T���˺$%A]��m��`�@l�K��»���7�P�s��G��B��8�� ��a���7�Gd�
ݱ�u����M�?k�,�{�L�?��-�m��,�rD)��eCtck��F�y��`�oć�n%�Φ�j '(�)O�@ �d#�G��%�P����L<焪�#����$�Q���T��E� ���h+���!fu�R�Z�^ן��6c,�t�c��КP�V��a�h�����H��^�(�%���'{'JB�4�)�G���hb��V�^�R��M$'��':�:͎v󸈟������{��0V̩�`7 ;G,V�fÍ.��cbx��/��T��|�O�0�0TB��ޓ�`o3� J����.9N}�sH]]��¿��^��Dw&|�C��J���ov�4��{�������>���"JZ5����j��
�r\� /�V�Oח�'*W�<Ďq�bA"�XWT�a�Eƈux /&n�`$�}�0_��s���$�����<zq���5�Je��8��T0�:�{p�GX��m��K�HD�HZ�����d��R#ѐ�t�<�]����yH!]/��X1�մ媱�acHѧYX�z|���9�I~�=�:w�����������1ÞA~�Zi�+�7x��b^)x�¥Cv�ӪMO"�v���ǐ�8}Q�t>=n%���P�9Ѩ�vJq�����bl��& E0�>���m�I����(a.��)|���X���0?�FM��PH���V���Z?jQ����1�/��p��9�_%B}l�T��]���>��^!Wղ�p)��G�|�����]�	�4~��FS�j}B�pp���q���/��^ı��bPE�cr_6������ӿ_Y�� N�\�7��$�|�����Pu7{��،O��K��rT�$p̼f�p���q/w[���b���b�h�0�<���c�ۚ��ۮs��O�T:C^?��9�2��*h�Kz)���*�J[IP�����%�3�R+<��p�Vv�_�5B�����鉱$��S*���*OS�z&�/����p�3.6�d�9�&���l�׮[J���$R:uƝ$\��hO����PK@W�ʩ�A�ߖ$>I��h�B��0�+xNb[F�L��=y�p�=�MO��)���߼<)�	r�_
'���z0�X'Nu�b�l�� �� Lj=��\q б_��]�G�[Sq|h0�ݹ?]�;f��r���s�4�~B[��P�p�t.�͕�^���rAߦ��a�S�}p{���H���q���j���#VO^*"��$��Q�s���=�&��+=8;dd�I��?���GE��i)���*k�<\ҐѼ{3���� M��oç����S�dhMl�
�0஫\|v^M�Dw��+�E�%�Q!C���y�����uh�8�����+e��`��w �C-_KeW.S�l3Y��/��	�8��X��6�~��ԣIT�j���5��0��3�&���5�s�
B'��Uѫ� פS�m}=ݙ�'\�j{ Z7��ve�����Q��=.�1��ρ\J�Q������lh=h2u�r;��ل����	<�p�j�.�9ʲ��v��>������%{��j(��548����V+�{��<k��TE�2S�3��/@%�Sx}eT�c/� �U�{����J��}������j�ө��������J_O&g�](!p���^��(,��T�[���bƍ�� _�o�A�|��C*-T���8z7ɝ���S��4��
�UELw�{��~л�Ɏ�߽֯��-����b�_�F�Ϙ��4hs(t9���1/:�.�¸G�r 59h��W���|�"�P�_��zo�W����Qݟ�ѫ6�p�3�����������:��9%���-����:�z���i"?5�8J8�dU���&���v�c^�R��в�M? 
�t�����Lg�����[v��)�ًd*,�~QZ��|X�Cj�ur��>�@Џ��OAa�3�H��Y��=Fqt�����	SB,�\}%�	�!9�O�X�=E�����=���s��EYi�A��Z�Wj�QRws	�f�o��y:5Ơk�����Jx���L�fPm0��pe.�����&T��c8�lpE��1YC����>p�%�.-9���LH4Lb%�HR��=ѭ�Ec<�P��@���sg���$�G���Z*��rX���,@AtU��eT�_�z
}>�a}�%�ro��}b.-%c��{1OL
gZ&�g�������ۦ���u��,������֘"�Vl�C�5�z�kR��$p��X���_
�PNDNX^n�b6Ip+Vr��<�3�^js��� �����"a����)Y&csp�6�p}Q����Z��kH��3��P=�;�y�m֞z �Ք�j�X���a�li�\F��X����9�P��}f��t�.��=V«I�喟���WS��^{G�[hż���@|P��l��`K�P�HX�b���:@^��A�8Qo֣>u�p�#B�J�كq()����� QM?�(�di�ﳱ�w+f���8uuΛ�+����B�Hd�Z�(p��~El��=��)ڷ��q� �,�}2z��#Ye�Y=΍
e��:E�]�19���aa�m����'m�V���%�q�E�[e�1������KWi�L�| ����2�_���a�"J6g7#o��m��O��WX8�h��`1ۡD�Cva�>	�6�o J�jd���J�����g��z�����n�$�.O�� S�$�<f� ���wj�TBѥ,����t:F�x�`^�m^�l������c����zZ�[��SV�0��'�"�}KQ�s@*ͱʳ��!��B����WW�a�w�(��e,�/�\!��v�[�G�*{�����Ώ:t,�.�R�b��Z��Y�p#��W�
�uP������R�[�D�6�Z����e�sw��	�T�,��?F�KJ)_�	V�14�h=BW�h�_/���*F9����/���5�O.И��~ l��p`�mD)�V.�X���/�'�N�S��C���˗g'T�^�Ne�*�����d�8"�^�s�0���ͅa鐈���?��@r|��F������Q �\��^�T&�0��Z�s��4�^',36�5߼+�#��}�%Q9��w ���X��Vэ|��ޱ���,`(7�>��ډ�	�C�!�J!����@��"g!J
���
��K�G�d�vȯv���f������gE-\ti�.��n�sڙvr�sfP�,Vdc'�O{<ᴖ����Ⱥ\i�1��G���L:����N�"i)"w�L����
���Ca�B�(J�wY����]�W<���ً��pL�B���5����K�3V"k(��r�&���N�Bn('x �͏�HaK��@a���{I�i��8�~#�x�,�9x���>��JE:'È�2����<_~6���� �D�**���y��H�-��͞�u��)E,�UE6��␲�?y�3^4�>�l�u�ѳ�C��9�q����sI鑰�W�*���Hw>1�%���m��u�܄���>'3�������N�$݌�&��p$^	V�_�{LT�ީ��ڣz�ti�HF-�6[���j��D���%�Wr�~�@�z���,/�R^W2���C���lG�X�,��h��ǆ���*�{ѡs*��fZʦ�ҞE<�z�'l�G��h�NFS����?(6{�I:VU�m«�4�`d�.��B<�q��8ulJ����1����
]�(+�/�"h��m�_ZY
כ�Л>�OÚ�FA�����hDU
�ND�m��g6�㻺ev��>��^-]X?�-I4�i�D8�(�~z���̺i�M��rv��])a'�x3ܼ�+�&>A~�83�
9�LB&���?Sf=G�.omr�=�Ĵ>Sơ.@�G�GR����e ����|��i&�ߕ/��+h����w���#'^�Q
��ڥ��[�N{�\|���d��2��7j���{��c{���4϶Pƿ�_��(���A^l�����w.�ã���A�2Z��k�� ř�~V�p:9�f�Ѹ�-2{F���׭�jj��a%43@hE���t]OSpO�^H\4�9ͱ��6�g)�L�}s%�*��NR���{��މlԻN}u��
���e��߄>,Kk�,�4P�4��G,2�}H������z]�L)c9�i/r�Znx�in���o�ޛ��Dw��8��2���Toq�y�8�E��&F���Hm=.���QV��Vq�U6�f�d�%9���t���\�4�䂎���%g��p��olj6	�+�~t�>��e�%S�+���J7�̩|X|����^� �*E��1P��NUZqeHa��]K���0��ry��e���%�s��I֒�-r�MBG�PZ���Dʖ嚟�)$ɧx���
�2�f� �M9E�w:�nSk&r˻0�WD8��~��N�nǌ�I�V&$�9��R��Q^	�;�X�(���}� :&?ףe�����a��*+p���mV��Յ3��7*�p�hY�+��(8�X�X)��ԗCS�%XG��A���d�%�S�dZ'xAщ3�'���{�N�Ӯ-��YuL���&m]�A���P$O�S{sV�O��}����v܈3
L�y JD�v�������D���_�M5�j��{2U�B�E>[��@�@a�x�Aܠ!-�o?�ly���%I����^���R(R#��{��=��wZ���H��2rh�#~��q�@kߗ\��ZaX���Hd�S��Ȳ:��`�>���&J}�t����Ffa����K�?Cl��3��m�!I�"�R����̊5!�"�R1^��F��vG��DQ=�ў�=%��֚��n���Z�v�΃.̻2��<I�)��:	�����zi=s3�ͧ>� �|��V9�������/"G��ԦK��߭��a�Z�pQ+�Km�i���<z�U�G|��>��~�Z�ݻ6E �y�(��Q�"7� ��)�l��lM���R�cִ�+Ϧ>�T"C*_��j�;C$��V��NM�H�m�������X[X�*�s���s���l^�;>\��d�1	6#�<�<�*Fyj��1��,��X�����!��M��Q��TM��]���7�KH��P�ng�p}�䈲+�� YP�w��}F|�U@�;l����%/�W\һĦΐ������g�;z��h��0�Q�+n,�W�rM�Rg
��_�Mo?��R���f���XUoD<a�Fe
��v�U�M%��'���7ǻ6̣��f�F>�孀��o*]��t�Wy�[!Dvj6�<��l�7���'\�k���q�SHUaP���ίv�"���Pz
pn �}���em�O�����i��mʗdF��_bpZpQ	�v/
~����q��`�GLl�w��2�*
-+�ՙ�y���R�yΗ���lgh5�3��j��~�����I"���j�y+�:����۵m���̽
+Q�WJ�CSo��ߥO���i���(�C��qk�q��������B� ���n�o�
w������F� If��A�3��D���
-�4�tI�`�b(���Kk,+�n�
������X���(�H� �v���n��g}��R�5����R��g��>zbT�nM����ǎ�D�F��8��у9�aU��3�(�W'(u����]���T�B��3�Βbv��Ve06=��W`o�H��ɀ"4#�BS����ls��7;�����+��㵅j(D#{1;��iE-�fp43�F�^#�Ӫ$��j����b��]hw�U��"�[^���4!�ĿLG!�t��pt�y�D�0��o�QFoQ�`�l#��;;��ʫT��^!��9D�4>
��R���R�mǏ���6��ië7�S�ࣰ�3�N}�(�p����j.q92�;�Eys�a�w�q|�e%�g��F�� |y� "n�����D�3�1j�fi7�"����OU��Jx���LEҹ�I��r��}CCz~ٚ�ȿg�P�����n�X��m{����k���y9%��}�G4  ��L�����^lMn��8&��(Fx�D�-����W��u�@������[0�v'b}Ń��]N�ɘ�'�ߠ��$V�