��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\���V�fnvx��ÍG_;�ȅe�~�>���9�>��Y;�0G+��{�����Ś!�\��K��5$�̏�ٿ{K��	L���i��ݪ��ߔh5�^���m���p*���Ѹ�h���=�׀y�:H�{U��d�Q�ﬠ��fr�"��W��d����*�H��|�����F�^<^6`g��Nm��5O�g�6�fLj8g	<�H�_d��q�^͡	�v�]��A���U	y8�-r���/!��/}���wM�$k�"%+@+"��v�S<s&'�Y '�[��jN�
�᤻��b8B^>���פl�i�>Y��Ȧ�|1
�S�j`��k�L�銼1H�*UD$�/]eRO��d�x��t�̡���H����a��MZm!�ǭ"���|�42�hcfRFzC��jg̝�ܔ�G���˙��]�~&xUf�>L��pϕ�X��!�\�t�γD�=D�w3�o����2�|��f�-*�h��ef�-�F�C�䬆�\^xÓQ���7(�yǘ�ϒĝ�vB�;J4��G.���˭S�`�� H>N۽!KY:��2�'k���6 �p�j�$�\n���}��m_w��*(�2ZPCsG�Q��V8��0�>��s�5�F$V3,M5�6��D����������uYx�(�w��z�M|������Ս�Zh?�M�t��������4)zZ4�yn�����|=5�t��O9�<��ODyo�I��қ�q#�<]���r�'O�f.ZiiV�1jf�� ��6y�n	��Y�]�����^�Q�~=S�� �u*��4~ϛl@M���CPtZ��C�{��̿�R���˽��Ӳ�/%�0�s�8��q�2�����P����$�$��;z���K�����}�@p�=W*T@��
�&��Ҩv�T|�
h�o��{�}�r%�ٳ8��	)�� l:V��Mpl�7�k-.�N�}�2���q��j� ;���KC�7�4VQ��K"��C���⯫��������R���P��S����RZ�X�ƚ��FO$=Uj6�
L�%r���f�|ג�a^��il�%����j,:����6�yd��2ى��ٯ���k��Vt���.L,�ل�Y��ռJ�"�,X��5��!��,@�01Ut�Z���C��x�ȹ�	T��s�4�ˤ�f���+C{��Dvg�y��K`���ķs���[h��%�U�u+��4f� L2�2�̳���6u���c5u�I���X��ǿ��Ѿ���!Uy3�c�>Mm�ݼ�����5͢�FbK�e�n7�Ͽ�׎�`������*8DZ�=a[&.MxSA�C��E�);^@i�C��ք}�<��]�H�'kC�ޚ~�3�E��(�+��{ݍ]{�{���A�7����_V�ʨ ����9�I�Q���-����=�0~Ņ�k��¦�Vs��xm
tĠ�h���\��q���¶���Q9vR��a��,�z��5@V�h�7�����4��R		bW��,<�����d�B�l�����O|Ҍ��	��p; �E30t"[A5��i�n�;�C��#�Y�N�G�?n�I�$�?�����lMr2��qadRȂ��1�����Ki��