��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�i��a
Α1S%� �uj?�L�3��TLei-3^5]E�$�ԑ�����o�h&=8-�t���?,���9n�8��kl��E�%l��ȶX�G5�=g��,���s��٦�΅^؝�xx�$VZ�Q��j�?#y^
)��|ՃW?Y�
�=�vZ�{�FLm�E0̶ɀ���1���L�X%!J]e^�vr]��7Gz�_�ŅԚmD�<�ٓG_�T��E��n�J�f��nw�2a��SТЋ5��$u��h�=��<6�q0�J�p�>���6M���i� ���r�F3ֈ��IJ�yC=z�"/�Vl�O|�E;�Ѝ�Kxf�;9>&���r�3.�6�Y�xKַPj�q�*BUs�5�J+����m�g�
<��8��'�R�a�72��L���<-�����/�]2��oB�0n���_�8�p"K��7řЌ��Ӡ���q��3� ���r��'�I+p
ڸ�M�}��{��xb&c�;���'W꿶Q�5�wJ��*KQؗݚJ`2I�k�^[|&���ޯ���{g����q�3[%��L��3�5�?q�b���a4NB	<O]���i<�ЎM�nP$�O��2�+ ����V�Om؟[6�8�-s�6��r�	���lQ*'�у¥]ܪ���o~�T�hܨ�rz��lQX�O���v9]���_����G��PK�xt�2y@%�2ލ�z���i�=q6������!��%��kK�9�:o�/J����6ZT� ��'7����e<�Dfj����@�[��_B�B�~�i�� o����ԭ�g,�)|�h���`_a\�4�����v~!c'��l��8�3���x��*�H!�'�/�GG�]e���i���\y�e�R�ja�t,��Rcuʭ�J�����PRf�A�6��vîKuWc�ֻ`��I@�����)�,1D�+�O? %���$��୅�m�ٯc�e�����>@1�N+7�]��C���ʺk	��|���~H1E!:��I��8c�L	ʰ2�M��s����un�Q�j�x�A�5<j3d����JPet�M� v�������mA��n�ΝE��>�m%��6�^ӫ��D��T�(�g�R���p@���[ׯ~bK&�+J�������M��1��{���Ifw�	�����d@�Ddgn�d*���#�=�1�̡vN�g�A�Eԛ�ZЊ]�
�9�C!�8vy��v�7�^7>ݹ�/Y���:����_-��>�R�����>�/��IָA�I
�mT��MU0(�N@?4���5ꪑ�Ч")��s�ӳ�NR��w^�����AՈ�����\#9���w4��CZ���iA�������i#�1?�{�k��g��X�D�5ζ�kAZVI+n���:�K7��H<�vVoW�P�H��;�x���:����Yk���	״���b������Ub��o`�3T�N|wK��J�C�U�矐����S����2ʮtx����&r%�Q� ���UQ] z*@��'yp0�y��!��m�69=�uB)-u�Ͳ#�ކ�<[!�/�xm7#}$�a��C�Ď[��=� (�u�O�zŧ�7Un�א�ӎ�]:�L �:�l�ɺT$�����Q�ዂ%�S=ŗϭl����v���7i�$8"�M��o'�vĸi������ej~;������&Eܫ=�V9vj|x�ȫ~�Kl;�Ko���\d��%Z������~����˳@Q�"9�wCxx��#z��X�5��D/��ЅS�s�s�+N�]bi*�[�Y�`Qt��?�2$��H����˜�i�}�ϱ0X�L	�*��q}�(q�v���f�{�?�ȩ#w	��O��Kob���i�9p��4�D�$A�^�\p�Q~a{�� ��l�a!��%J�T��h��tlIE� ]�����0�,���I{��T0�qb[ສI����F�Ջkn�Z{�;'��A"6O�h����l֤�5�v���1�����l����(^5B�Սud[G\��p�,���yK|3g���Jq��ƾw�(�[x^�'#��8q�#��޿V����Y��.�.aV&e��
��eX[��F��̃u�Ѥ6=c�p����v���۴����d ��^��'@"�\	�6�?����>���0Z����r�}J@T�_�\�Uov�.�g�n}->���@�*Ɋ�X/�5�_��1�����Y�N�q�ARQ��5�Po�P���N�yq����a[ں!����/2u]!1����th+z�#���ʼ��`��h�5B����Hv5��#�[�����~ۿ�����E��a����ݢ�m���ϻҨ\��w�7|��'D��z�gɂ�I�Sl�=a�'4B�͉�6]�[J�^�Ϭ�I�?�F&wN��uJ��9�TQ.&����XKy�[�����@
���8*�eF؜,���]�Cf`-5���8-g{�/�E&߬"����Ȋ�Y�纷�>������_��3�oGI�[ ���
�Y1�@�p���!ЕqP#ۗ��S�L�:�9�zt���*�1��1X`9���NkNrOh�#
%r���?I�������=;Z�t^͟h]˱��.��Wܧ6�W9����g��V1����U�}i��B� ���b4/a�� �\#H~aW�{�̩m�
k�����{�ì��6���=��*�J��Y����ݥP=s��gpH�q,���c �[!�&�uh��X�m�?�+]G��dg}ʔfo&���ޝ^�rgK*����esӡ��i��G���zq�������AV_wt��t��q���0~��H�xtZ��?E�����)glȍ���oe���N$�N�Ä�D ��&���VC��1]Dee��P��F�x�0c��6��US0�c�*�/���ʍ�i�ߎ��آ��ZI�*���e�j���t���i-�E&<Eko�C�7�[�	����2nS�%��S�7�y鵩�Mt�m��(w��tO☈�$o��Z\����&��b��/'�� 6C����)!�����d��� !��|�������TA��ѩ�mO��'��xof�P�bqB��ӄ8dk�$�y�z�-vl�o��-�s9�f��Z�\��l�>0���A�7�6�v�,&j���uÉ�tsA���Z��ЧT~K�ۼJ�"�*�����+J�o�I���4�v�j��P%/�+u�[�c��W�A/;��:M���4%e%u���5���s�6bN�(�~�{}�k��dd���"�	F�N~G͛r	�;��he!)��#�4���N�r0[S��8q�b�	x?��&O���IN�a�h��6��8�����؝ ��ܯ���!�ȴ3�9�!/�\���=07����Eg�d@�� Ok�>�����PF��l=�0���'�2�6M�ﯧ�2��S��P��Xa%�	.���}Qv�Y�<R���t!a|Gn#pTPx���T�iF�k-k�ˣ�i〗����M�k���lB�V� �g��t���ij�@�ש)���_��5~q�#��8�UքO�HA������`���0�O�B3c�rؑ$ �#�3���7y4��h���.�΃�v|:v�����~�y��U�Fϧ"���;?8k�0|�-�E�O���赊�C�I1=��xr*2	���2 z����j`� ���`�l�Z�<PQI�+�,Q{�+>ni�D���D}碀īQ�2�b������F@\��]-��yЕh�����\�:�	'VxKxY���r	���J�p#e�A ��*PZ����I���;�&G�NO7�'�̞�@?��Y�l�|� 3�����C��n�HQ����6��l_�I���?�������:в�z�XX�|S��^������mh��19)����e4��sTр7�b�� 9�s��9�%UO�#.`�3�twi��O�V�ې��*W��6Ǆ�(�u�^'���d�Y�~�M�%>��ޮ��%�oߗ�A�Z��!C��h��pD��Z*x���k������-
�%���m��y�������UB�ұ��k*�m%����NB����>��[İ����}n�¹����jLW�+��(��ԙ5���JY���!*ix~�.��e�Xj�O$�z���t	� Û�uy�Wєށ:4U��+���g~ꭙoQl,��u�T��L�T�|�Y乐zk��a��)~��M����hT|,��*?yaƆ�n��1��W�;��S<�뉥���%vt�r�`vƎ[i�AeT���{�����c?x���=��v6BH�}Ϧ���]cd��~� ��>�ߤ�d�5v}��pTȂoU;�JG�#���A�2O3���7��.[tu��z\�*S� �p,:�ZS�W�%mi�2X�D�#ay��C$F\B4Q@Ų��>J�g����~Z]�՞�a��O��4W欟�9��)�z���Ph�H��<�70 ���M0fd��@��Y�4��ğ*'F��Rŗyf�蟓��_=�B�Z\ɋ�ힽ���$��,y�$�ҁej��
�@Xy����=<����n��7?ܿ0�t�pK��3# �����/<{*G]�vg�%����چca{��.���;��a>�蕴<
>5�	tF0T3S��{�wZ�pI7��e^��J���'ҟef#�f�!z����u-Eq�M�tI�s�az%��4r}O��; ��ㄮ�e���eE׾�a�R1p�ab9���1b�d}�����8�JW����YMw�>���<U��4-*Uq" B��pL3I�0�����̅9���:Ҿ�ڌuB���9���3z��2�h��;�����'hs�!���1P$�.{q�\�T#�?ObR�~ �o���1_��H�P�r���'�V���Y5!Zin�_�n��w��ְ;��.d��0¨K��]Dj�8&rnK^#�s�����T����txj��y�I�dH�cZ��Gq���2���N��{I���,���[G�"U��ON�Ƃ;b>G笏*U�	i���nZ�E�a��=-�p\CW}7,�9{�p�L���V䑦/J�`���j= {z��\ڑ�!�zܗE�O�*��l��1��k)>�t5ӫ���� [�g�(Q� n�zfY�@&ʄ�{�Z� z_�Xԡ��S@�T�e�R�+�^kUb�ԏ�3��?�e`O������!a�-G�瑻�y�9\��`F�w�%b���K��/y'������5�C�8P��ǻ�ϟ��z��4Kg����!���cB��xtC��b��t��V�
l^BǺ���7�����9O���p/�K"�"[|U�jL���܇���m�,�0��!�r�,���A��_�On�����f��1��:v�|ݞ�ᛗ���CúB�-���r�6���<0�Z5<�/#����%8��KKAh4�s٦�=Ѩ�m�C�A�j4�9<̮=�����BN�N��zy����Xel^*��P�?�P�FQ��<L�$E+�z~��Mш�6����Ӏ켫���c�]�fZ��{��,c�`�����7���"���$O1ך�tM�4���z��va/�O-���e6����v��G#4��K9���N�036�8tX�9��
�uH���)v�Vo��N�9\tx!MS<8f�:ac���WH�C�'����諒�
ϛ55�l��O%���V>���j*�.�g�N��y�Ĭ5kA�2s��F˂�}��/��XZ_l�����!*AE���6�)���hk�������Ge͋�{��:B�y�ilzf)K��lk`�\����8Şr~5k�`+C>@M��0���k�4!0��/Tb��F�^o !���h�Zs���<��;6��n����4.�}��S/�8�8�t�j�Vuy��! 7A
����a@��������1����H�7Ro��RZ�by��>D$X���>��}ȕ��=��#+�~�'��U�g<��LB�34���Ka<�g���C�k�#O̅ǯ+e�G\ em���Q,߈�����#1;��������R7����Έ|v��x�d�:�z�r� թ�x�����@�����B3V�QF\<>焜ۍ�O�����T��`WT1� �E�7��]DDS/�ɇ�OѬ��O�����{�>@N����s�h�6�d}6��������e՛+m:V��	�q��͜h�|�l�}�GTU�A\q��ź�}?4�aS���M�Ղ]�r��!�%tH\��>ȼ���2�?��o��iFվ��S1�����	�8,�I�,�?��M�ܲڇ�
.{�_3� �Oh�_:��7#x��t��֠M�el�^�4��/����	,�J�Eg9~��dwBs)��ҘvY�|��T;�'ݘ�0�;� �U����U��Q3��A��E=�y��kU���6������
mA E<~[�Wi��/E沾|f�_�0�C�����[���4S��y�{3~�O�fl�'�-�jTs��*r�� HC$	@��t�6��LV�������Þ�~�n���n��!X\��tT���?/��Db� ԛ��:8��aKT��&�l$���4�&K��s`� X$A���P�1J�2�F�F�\������6w�&́�# ���g��^�/�,�s�E[���0D	���3��e@!%;�i�sE�`�K+�5��rf6��讨A�:��ᵅ=���ƿhs�zY�S�#��ro��f�t�z��tǉ�;P��h�^�G�W�!����.�����r��p��I����e��ʕ��{�QB��\�*�ܛ��'����J��L��sw��U�S��Ͱ�"��UKh�lKY`�lNw*��y7ƕ#� �|Cଫ,Y�#I>��T��t���6�t�Z|����߬W�M�*���O�3D3e*��{�h����\{��I2VRA��g=K/rO\,�C��C9�;�M���fHBq���9I�!�W^C��d�P�	��R$���PC�q�8�t���О��HH7&�$�g�rּ�y�I����\�8UD��E��
�46�?�B�n�:�Ƿ�%$�~Z���G��������D��eic#"v���P�Q�8����������xO\1t��IS��l�� ��E���p��ם�%z5��8T������-�U����1a�,򶴗Ŕ��:��"?#���1�F:Z�{��^ut�,����g��<�Hb���$�'�}����L������O���O��	y�H�hm�Th���9yO@�S����ی�������8ִ�D�9b `v�=�i �g�K��}�B0�$���i����_E
bN,����������F�,�L���6'�>�-����/�%�s��uɛ�$(�-1�hQ�����9D��Sc(!Dp��n3辔~���J{fT�Y]���Ii���5'�����k�*�B!�%�1�-����q��1��p�y�KIu�����q*�o��&�C��v*����&i4R��4S�1�ȎX�0K�� Sia�6�Eap��:ϵ�N��I�)'}
�2{�|�%\%��
��|Z%���ع�9�a��¿�Iـo,^��i���J����ʧu�6`�i�L�^��'<f�ūS��*C���\��\����n�8WI�>�oҿ�!��ʬF�B�/ſEi�W�Y���遮n�h�pJ�����K��F�_׷�X�=��T��+	��C{�Sp�d���n�S�V��"kk'o��4ԩ�ŢE�{f���_�愡1�5A��b��׆�����uύAw�"e)ŗ'�Y|OC�쟬���K9x��Rx��'(9�<	�xt�k%����K�h�9�n��#������6H�"p������0W�>1��Ţ��x���K�+F��]c,��4�c��OX�".=�K�)M�I�p���8�4�
���c������OL�M�=�%(�@q���s��A�z�/sRy
n?g!�c-�o'� ��H�ծS X�/���1~��R\u�(1�}$]��ɧE�x�� �?�:��ݤ��x��l�n�/���!������)�s�9u��+���Zv��}I���X`OV�u�1����4�uU�丯z��A���6%��?b��4
N�u����B46U}�C�S��Mj��S�c `RܢF���J��@��>i �BZ�R���'[�ɰ�x�40W2�F+�`��_��˩-��Ӯ}�*�~�hd�?� �
M���|{��lU[��?�����G���'M]Wʏ��g>�_Y7�d�����=����i���ƃz٘W���#�4ٰ5�Z�"�@S�r�
�Dy<���%ig `�\�${�����S��_U��O���?*��k�	�>z���:= �BP#�Q����J�.C�Q�`��v��"zB'���Ϩ�Ĵ�&�(jPr�dM���g#��f���m�^oB����妓��꒫�_��y�n��w$ߵ_�U��B��Ŀ��I1��U����B&y�.8��R����RL���^K�ļ��ޡ�����s�첄KR7B�9 ˷4!W�BS�����A�#��'��'���x�����Ad�,����pLͧꝮ��:#�IvT��Ǩ�*ɶB��R����;k���5���_X�7�0ҭ�X�B7S7V��#��CK�ݾ�)4��\��02G�(8����W%�Xs�~�8�ve� ~׮�~����*�;V���J���--6��j�Ǝ��#m�Ytn��y��3���C^M��m��a�EQ��?��j��1��� �Z�l-G�;2sR��w�Z��F:qp#���͔�~���yY�U�����d f�\f�����.�s>�8� _��5��4^��t�OV�k*�k#֊��#��4a�9��!OMJ{'Sܼq�`�t��l�{1�1-�_!���4�2���/6tET�S�"�dȤ���(�wx�� ����j8%�X�i��<#��;{x5<��sz��h�@�[9�����jt/�O�ɇ.+�hQ�7X�����eH�Qz�8���ѻQ�@@/I�{��֋#0�S�j���Km��ʴ�zX7E;�(��.�d{l�Ρ:O=�m�����Od,2 �=5�{�BB�?A�Q���q�:�ƭ�����BR��1!�#;�h�Ҫ��mka�n\d#�����Σ��Zj�(6������+�Ii@����ES��d�8��L���q��W�����E�����M$���3Fh��G2������O/���-���W��w�A]�?��_�Cr/T���)��.u{��a�:���N9k�~͹�u����G�X�H��:Km��"�}���t��̿���~X�ڟ��	�ga.��*%g����^yFY�[��9�
���c��!sun�3N����7$6���,S�ĝ6H䂖��!�@6�W�g@,`Ð��`�J4�1�+�B�ЯO۞�v5���� e��9�6Ҝ��$<,=0Zǁ�=�bw���=?�X%��f�g譈��n_�J�#j��)����1���6�cR���%,_�>�\����5
>n_ĖTA�3K4=���>L�5���iύk4,�$�D�,bv����[���{�v��94��_�X����Qq�Mx8��]�{���H��
;�����RD��!���Kf���J�w�@[�Z�;������9E8YO�s/�+`�����G�Y����
�Q�S�_�bZɞ�UdQw�eD.�y���s��61@�v+�������M���0s���#�C�k	�E��>=��럲��5���,�5mO���b���?e����=Ʊס���M�İ�":�ŬB��%:���m�ZB��⩾n�v��ti�%��Uv\�ʼLV)�CRl�;�@�FԾ�u���A0��=����$�n�!<^��IP�sL+�p��ә�A��j2�'�d����֟S
A����8�g99�7k^8"������Z=i\Wٿ�p�o�"�4�$��3��J���6���j�}����t8��֥��!ZÜkoi*P��?o��.I�]�l��6����`�*D��#f�WuN'����]��$�/�Rе�:�}�uh2Dm�"��T�Tʰ�f��dz�7A�dc��g���^(I�������[w��h�HTd�'���������G��Jj�j�i�Yao�{Ā{1��WMC޹��9�d8'���`N�'W�UK�13�~A)dG�A����b��Fn�T��*����A���^��hep��� sQ��c�f@��h�W��1%p-ocܝ�*1��hB�H�Uh������E�#�_�g�l���{�Q�����8��̙�lq�Nu��5�*ǭ�7�!��#�8�ݰ���Z̥c7�e���|;�ν!tOc�_5ܻ��^*�)f5�'����gtJ�6�����m�'��u�D���Pa�;��h���Q!�����hFޔs��>����|�[}�-9��&��&��$���qv�nw��I�e��X�p�I���X;!����b7����|ଢ଼O���ЏWr÷v@@ɝ�9�����ed:A+�sg,|MQ{	`��)�:)~���ƏY�k��^�h��r��2vUa����}	��)Q�;�H��r�nJ���z�S��� �g��Iv��ɏ͢�L萆�~ٿ!!V��W�됝V�CqYh_����_�L� ��BwIZ�M���F~A,�%���N��p=�[����k���	�c4�-�g7]�s��P7�m�MJD����^g}LJ�k��d
����c�8J4�?ۊQ�\E�f`w����l}��\��3q�����ĥ���K/���ųU��"k�C�����-�$q{�w ���|�z�C�����n���m��y�����P��+�7�yO���cW$��:��FY���>�U�Ç���7+H}����\�hF�D!�X�s��s��2����¤^F�~�w�(_<KWK�F�@$ym<�҃E����cx6,X���v�c'T� SK��)5z�������p8"~��ر�r�u�R6B�/ͯ}���]��Cŷ«��i]&8��|D�䂐#x�#˛�Um�4P�R(�=��T@Ϊz��"��s�zm�vQ��)/��σ��2M������<&����+�{�������z�.&ԥ��{��~*p&����
��;�g��{Nl�^��k�ۑ�+�)-�p�_������9hG�*`⸊��8����c���C�s�B�+����hi����2���Q��l�&�p����y��(H=�����[��������j�jg��a9� =SدVm�-�m����g���+����J[��6�U��3`V���JC7��l���!�<��P��X��}�n
�-_r����n�����VZA\V�������H$b�iAD�ε��u���
��hxn�fܘ��YЮB�8u��;{g�ڙk!n~��1H/�e��d�+��n�޳ߖ�P��|�s?\�%��z:�?|�0x�-�޵9���'�*���*,b��0/'�c�DyKwY�Pq[DpA���c.��S�޸��Q��*����cN�k�͜߶s�KN]����53e��7=|����*�N�O�oVy��[3#����.��=�xL]���K��d+j(ˡ%2��]���4�@��`m�7Д���@b�;J�����;�������._f|cר �<����5��Vvar�>�r�e�>�Ez�w�߳=~+ޮE��6��/�!'���7.�k��yFS�)�`a���+u�����d���W���� ����Z�q�$|�;D6wϼ;�tQҩ�ף��J��$ďܕY@O�$���TA�k�z?��}Z���$�M�.����i���^����bW�c�Z���-!����S6:�����\������~��f�0�1U'SLv����gTٯf�;F D@�O��X�X��:g3��U�=dq����0�޾���F� �p����v N�f8:8eJ���Z��0F��k�S�YTLRN4�b+-i��u��E����[;�v���kd����Q��X����_8�	����Z�J��m�@���V4�f�3�CyEME9�qQg���&���nt�ڳ�y߅|ͭ��J�Ԕs���	X2E�.$`rN- ��.t�G�&&7����7Ё��J��-��fۍ�@���Z�����]J:��ތn�])j�j���}^X��L��b Lp�KS#�IBFb�7����Ul۫Ĉ;n�܈~3��i��5�$spC�#�$N.K�Ħ,�s�I݁]���جd�at"���T�G�����w��$*�sn�4����'�J�aѵ����8b7+$*�2`�O.ϼ�b��E�`�"g��1��� �U;��KD)Ǧ�8tO�̶)���)��t����2L�	z�Q,z�(� 7��E���Q
$Cv���9���@�N3h��܈0h�<�<W?n�a�֒��@6014��O��0�8>��Rm�*q�§[%��W:$��>]+��51s*[��q�h�!D� %�����l*':��N����"Iy�ȭ�F��F=��������"H@�@.��==���t��s��R�98Y/8y��/7_�0��ds��Y�@W����M��8I����K������o��6ycxX�5���+�o���Z#D��N��z�D�̇�:Ӯ׫
	��0RD`��;��1Wh�ӮlY~#�эf#z�t�=]�ۘ�����f�L��~�<e%d�ۆ����65ּ�B��ئ����1�$����S��,�\>"���`���̂P��R�%�	O��јDp�4��2�����	7-IȆ9�՘(�eO��n���\�F����?�n|�ͦ��{����g��M�w�TfA1�zk㢘�J��Ivj�c��ڒ(=?6F7���Tb��?y`��)�M��@�ʹYL)%���L>��$W�ā�Y��x�c��n@����2���ɞkh[�[����(�=S\s��r�KtD���Y�o�5�(�a�q��-��=��ɷ�p���[���?5�*�5�3_�Ү����@�m_��kGᬮf�/�q�_����%Җ=Y��a`]�\�����ChJX���Q
���]�#캽��#�A��vg�	�J��A��r6�CZ�@:��?�pp�-���5G��r7��<lE&R/Q��z�LN!7/�]��@����Zp����dؐ�aзq����!�#M.VU�{��OH!q
���G5x/���&��R�g�>�#V��Dk�nL�2���;�m��)���:J��Et#��1Xs�p,x4ׅ.�����S��8H���������T�D>kj�Y��-��$u�����n�|U ���,nۻF@xt:��mӯ��H�%�߂|��W���l�i�G՗��W6-�$t�"�����\�J�>���IES���ᄿ�O���&8� ��lt箩�V��-x��L�h�bH�
?���Fj��O��tQ���k|�g�[�4L�'�����:�O�h�%�ڝ�o�ee�,�I�H��2oK�آhv���υ�[ �n+4�.;�5�b9�"�F�
��ť���ny���t�H*B���� �B6��Gi�k�1Z�u�	ͫf��V�?�V��wY�<2�p��_��=�!D�i]�g�\�y����^z�e��;�ـ@���)]�c7��$���4��^�IOj�4]� �NEa�!�^n �r}�ˍ(Z߂�p��D�����p#��t�l_G�D�������E�6H~�mM��[�{U�s��+v��A�����*T��X-uxf�$5�o����Ap�&^�	R/p��2�uJ�a�zt�y���}Z��&��F�hG���m cu��{D�A��<M
�ϴ�~e�60;&�x�h�a�O���t����:�z[���p�4��_��%פ�ds�,>@E��:t��< �)�^�Ȕ��aVp{"@~�F2u�~�f�o�<��e�߶�HѰ �PqP��?�k�V�N'd��,����;(e��5�qO�ˁ���l����:�V����u�U�\���������D�l��1��Z1��FXJT��^��u��]Qw�5(fZņ��;	�M�~��,K�!�����������ݻ�d�j�!R�)�O�`�d�����w��j�;�9����#���)����b�l	�s�f�̋���!�Rf�Ȍ����S���Χٜ�`:���l�a5\��U8VPo�d�=#(/���j��5#W�iZ��?G�=g%�R�=n�[���^�F.ӇB�IJ�P[�9�}���o�n���q|]�8��s:٨����}�����k���n��<�¨��?9���Ԗ! �i�;����5�
	>��Y��L�;w�V�&�|�b[�M�O�Ey7|���$ �0�#��u��2�܊y0Lwg���f�������] ¶��M����~Z����'�xpa�w���F�V��52�]ad��C��R�G0�$�prO@�::\���E�od�iy�m�b�j+���'��ϋP�.��M,G�?�v���~����.�nsNk��F�/��#���H�������og(��['ar_�>7�ž�Yn6i��Qf�-�r�#���dK�c�#�EЬ�A�d�'�m�\q�1H��ʄ��#��?�\E�ew����et�r��#�d�#*��bWb�nD&� �G�AO����!t�o-�<��i�ڔ��0,t�o���#�����~�wv!fw]��K/��R�ǳ�Kx�1Y��n�LB�A�¼cW֘�D1^G:� =?S�Σ�����j!�+�V�����o�Ƕ�����)�����DrUM�ig�L�3mQ�Cb�;��JT/�͒>m�U���1�
��/��T��j��*��İsG},�Lm���{U|ڿ��[\yc��bs�)�V��lK[0,
h�5e�f�X���d���>���wa���1vkp�`���D	?f�[�8{J�e�3f��H��DD�;��zw*���L������肤 ��A�ڪ��3<` � urN-��
R���=��	��(�������9��U��b�9�v��d7��T���۔]�~`7���i0��^�(�5g�l@͏���3�a�ܪAx]xyQ�˭��|'K%�l�ϩ��/�B����f�Vh%<���,-q�gV��T�:)��fC$��6cLX��g��]�慭����Nm�	��rݙL��L�tپ���@.�����/�M2@���oSt����X��1<~+
����r	V����I�[���VYk���+SL��@-e �GI �A���0$t�X1t�4(����?
����L���_$M���\`�2�YU���nh#ޑ]���B�2Y�ٯ5$�)1�vb�&���V��>��U��:(�r�z�,����x֡p�m P�$�������v�'��f��a�n�`~	���,�?n����Gf��X����<� 	�\�Bn aǞYq6k�6pV��L�%D^�Wę�)	��T�}��hy$�B��g��1 ���
j]yh���&�R�e��3O,���؃w8����6���B�\3'U�c۹��R�Z��G>7Y�-�ʑ$QH/�+w\�Uy��rZ�}S�/9�����hd H��V�%��;�`@s�	��p6���|��W�g_H\����v��ݩm���xZ��[O��su��IC&��	+r�0�U�ɏ`d`d?�+�ĸVpQg��%�}W�-e�0ˀ���B:�+r��Bz�I�Ri]a��ЌU7�OD2�ag�z��LɥD��ݔػY�?WO�A��Дƕ2ީ<�r4�s�b�?l�ڝ�OrUmX�/L���B��&ok����՝r��	9:*��a���Zǩ����}����m�� �%L�
'���1�*-e��Ա:1���F�=^�Qj�6�N��47��LR���k_^'��"Cɨ*	�MU*�|�&M���`�>�i@6��|�xLf� q�~|����k���Δ��R�� ��{�Y59`M��Xߘ`�}^����Ȳ���D��m(<iG�lN�D�"E�/������CޙB�q��dŮ�`���r����W�uu�k"�*���7__N�L��<Fss��"Rw�q$�
 gx��D?2��1� oR�ͬA��b.��j�mb 3��7������w�������e�)�l�]q���������r��f�-@V�.�M������۝%�}��A0ͱ��*'�k���!��_�d�pR��	M��6F�T���T���\��s�?k3�i�/������54��������9�09Պ�4�sg^�H(�nM���.2��Te��\,m�ID�Ф�i�7� �[V�&׵����P���E�6.�i����,�wV��5*5J�Z�G4�pc\�6+�d�v��ct�/u���=����2�R)˽6b,�;F�O��0��2���X��#��(q��D�E�R�S�('�N��=��V�g��@�.z.Bc�S�P�˵�9V�o�����4����Aw�$���:�������=�8�A�6�N�o�Uv�o�NV ����vT��S|�0�W����p�)�U�����:���r�kfk�E�7Y�Ԍ���Z��>է�S��k��H�twK��hO��܆LΧ�?b�b��%;C��*���n׸*��Vaz#M0Mp��	q?�en��(O'���!����sL��ŝ�N�]����X�+4 6�v���d��Od�v�/�Ӊ=��szkAb��j�Ġ�L����GV����d%�A��氿Pޡ\r�	]V��&�	�G�A����v[�M�2����e$ś�'寧�C�d���>�T#5�)�V�tۊt�S����+�O�Pi|�˨��;+�Q�R�lc��nj��
Z`j=)g�Z���!c���3�tm��h�-�6+v��o0�J�5C�Bȕ�֎T"�X�"��*��f�$�:H|�)[��訉�W��My�0�A��+.�Ͼ
������x%�w�W��ndnnL��R�ʟG��q�C~Uyޞ���P�� 9����k J�j��Pߨ��y4�7�ş��d�"`p��x�]<����$JjM�d���dӚ>�����5lf��C���:�K���a��B�$�%��!��q��5Y?�|��I�	�&�6L�ʔ�mk1�i�^�ف��qr� 	����=\����}���xn���\�zVeHo{D<4zj����h?� �_��5�
�|&�c���Xjgd���/l�����;!��>��*���֔ZAv�Q�� �5��qG!��� uWVl�����cI{<	y�x
+Mj����&�^	�"�����'7_��κ��S�
e%��{9!@��,��uY�.��=^%��7���f[H�Zd�
��U�*Z���MO�e�u2{4xf��� ҙ��B�ph@:�kA���
��Q�ʮn���E.���'+�0�e˳j����%?�u����\<�Yb诟1@P�hT�/����E��!�<�>�JZ�G�/7�5>�V��%�M�(�+��앵a�NC��*��:��V&��_(��<1�:��,�$��F�Ɠ]��{Y�q�fB	h��g���$�%�H�'Ź嫛��,�|�����'���x�pT(��0�)�ZWt��j4�V�ٕRe����D�nRԙ����(����6t��zl�0[�ZNr	��4�L���u}_�%�Lj����\��gA���� N|l�I���6w�_)鍇�9u+<��[h@±{�\!��4�*$��%�	���{��M&Ƕ�ߞ���]�p���s.U����]��m�b�pn��3�L�
�Tȫ}�"ﲺ8�1:W�T��({���'����va�l��
�ݻao�|��y6� �/=�X+w'Xn#vt����*_ϛ�4�S�"��_�U��:7>�~/vG+�q�x~+1��!֔`{���'v�azZ��Q��8
��n��n�p�G�P/���*�ҩ�<>aO&�Q�֜���=	�o�&�ݢ0�/1��@�y�٠�l���4cM�w[�\l?`�c�t:�fiV��lmy�ӚԮ��bh���+�Y:�Ej�l��u]�_���X;�|��z�)���tm*�[���#�H��IƧ��5s�Ȍ ��3`�T�:= n����	
c�_����r	��{#t����/Ck�߂�I���g���A��q����ݰ쵌^��-T1-��B��	Gн�apZ��Z��y�H�.���0�j�8Ϙw,�L�����bT*�|&G�o�R.N�����o_�m�?K�̨#���Й[�x���_��;{�������m�`�9����3Vo������i�������.l�XWD�R�}z��2a���Z��dW��DS�9��bY2�F�&���&�ݣGĉ�D]xp��s���c��`��&-�E�L����I�7���u0�>E��G����J����˜�]D�pO�Q�#����f���@�R4�"��?�)�I%E��X�ʻWj�f��{�2�(�=�ޱ�r���.���U�������%��\ſ����!l��P���u	>S]m]=�	��V�ƀk��NO��B� �-��{��_&�9�d)��a�F����%N�8��5��rH�Q�SRt������q�:�)L&x�	�Z�R~���vZTw;fÊh�褜�I2.��y��*��G���z�.�E��o>��p��dé��f�E�ׅc&1R�A5�����-��C|6%adIז���r8t��j�?����Q�;��Vr�Ri��t�ʿ�w��X9k���MښLKM�x�xՍ�I�=-��b���iL�U\a߮18dz����]�y�n�:4�s��Ӌo\��`O�r@Ϥf��?���]}�� ���bg�|$f_�����w(�}-�,h��)}`��m���+҉��7ߘ;l�9eb�u�N(��sa��Q�жX2 ��#�m
� ���� <[���.w��w��i�t��yEU')�^��z%��^�t�&Ǝ]F��ck���*���۵�[��:V!p�`2T��������zQ�2k�� Z3&�y�03�]S4A4�yI��a �%���z�d{
3^����P,K��6d<�]WrEm�v���&s� ���2ճ�|j�����z��5��yt�n�4@3q��kѺ�f�`�5o�����/FX��N5o�����=w��2�(~�^�7�ۚ���z����)�J��� ���ѧc:{*� �j��Q��m�� r� 4I!��\���~�m���*�[����Ua���!�B, u����%ȯX�y��� ;ʭ8O�����$����5��Y�LYh�z\}��E4�*���D�+�Y�PEv��|"�eɥ�;���w �-�M-�y%�?�+&R�d:��_��b�E�+ݥ��F;���
�};$lCUB�¼�P�U�ӣ�(d�&FmN�.w��\v����};�e�9"�����  ~RB�Y	*\3��d��!ά}�|��C�^dW��u�ba���\宝�De�p�-��"=��ig��g�l���^!�,9S}�>��K���YU��3��g*��חQ���aW����F��~$oᡧ�%6�	4��#ً&?,3D�⦜#��k��e���X^I�es0���Q/A#@� ��O痪�M��5�p3��xB�J�0�s���c��z�w\�����u�u�B�������ur���f��V+�x��k��y��3���bֳ,�t�������B�0�Iةt��\�s��.`C�	;���(��x{���H!�(ܣ7��g�D�����ֱd[�xn������[�(�Z�uU\�ŷ�7�f���VS]� ��YW�WkXW.��/Ym�l����Z�Y�Bwm$����
�l��e�Lټ�4K5.�\/��,ϕ_A�]�8�^)�BeL�G�5bE噆�tr#J����?q�Ӌ�Ս�N:CYr��ͮ�q�+!�|L� ��r����^M�3s|�SL���\���'�Е��M�W��}�f=W�m�"�]Q��'�>���l.��~1֟w��2�+�=����^�y5q����O{�>bL�.��sjk�������5��Ɗ�QDFӆZn}ڽJ�=OKVA�6�y��Ч�镎��?�R�J�M���e�
�z�:;���h:iUdL���sm�A�T����&�2��4���ǢB0涣� Č4�:������h�D%mۜlԜg*xɓm�0n�T�0�f_o/�[����f٧��!�a���h��8� �b</7�(���o"O���}R��{���d#�19�&�h�?0F�G`����ۿ�m�f)�y��6��pg_�pV%�K	R!Bd��b4�"{$�rw:K;2e�*����������إ�tA�k���[���q{K���� �����_� c<Ƨ�H������l`�ԥlǇ2�=��R|�}.g3�S��"{u��9Ԍ��gYB\M6@�Xs�v�FƗ��wC�NO{�r��u��T�kxJZ�R=�6�x��B8`f�a�����*V�҃�?<�X�f�H1?{l�Y��Qʏ�HV�=�F� u!�)%il�����Yں�u��������t��F�$C�	�:������yƷj����x~��|�+�Z��-�ucS3�AB����Ft������0`���cB!PFC�=d��|w��
b� 1U�kϕ��qU��6\��≡�' ����Q)%|��5�?��0�nH��;�2h�3��=�\a��h��	(�=�HcGx��G)� �K�?�����0��NM����a�����'7<�T
z:��ws���?�E�=Q&=^��jB�P�a���ҙ�7N\���ܒ)X�+E�]�W鯱����WB1g �X0�u�(ٖ�[��A�X�\4��^B�ql�yI��tX��%[\����w�uCL�-�2<�{�E�: e��۾�''�r��X�3{q�SJ�T���:������-x^��ӿn����We��� �wd�tD�=�A{�MTq��HW���y�'b[��� ~R����h#c�� �q�x��]ҫǺ�p���>�u&�3�*��4�T�b�vO-��d��,*gT ��sh+��ߓ����m���%�<.�P~�����M�Ú������úd�Si�:�B�����T�Yfx�ZUishқCR�9v���9`?� �D*F�2f
ћKa5i�9n�ד��rg���Ɇ�Ԇ-l{Z����K;�K������I	���b�����%{Vf�'_������C���N<�-�7�3Z��O�����ӂb^�V3&���j���<��Ld��=^z��뒻3k`a����ԱW�9@\��s�&�
NAd�>ז�tP�a�+���/%�w�K�eG�X�yc}V`�(5��Y�,֏�r��J�/2Q��=I�M��"��~S��r�S���c	a�z��adVJ�O)�����"&RC^����:;v�.@4����r����W�$
	���7�t5c0n�-�g=�����̕w�Q:&w �w�R���~���Z���|���� w�1p_fr�ݖ&�XF���^�u�n�# �VT+U�W�`}�������\���l(�4�¿;V�r���OS+�����:xI��*�ߠ�|�=�1 
]b�6i�`>�A1q(KX����!1<(������$T�<'�	�	� &�������VJT`�VE��`Fk�0����av@Q\v�U��X��H�0�eF�i���@�Y=���!�� .�c+F�2��=������������L٠ͫ�p	C8GQT?��oþ�#pVٲͳ33W ׊32�����\N"�۪��H����5��S5������yΝ8�����D��a].~�,&���,�	�䶭�{P2~8y?���^�ߨ�|�4	o�&̐�S#/�����n5N1u��n�=�0�v��'[�L��:9i:N-f�1�nO#,,ȐP[Ad6��"@��U�o����ɭ�(�#�(��������6�h�,h`��rW��s{���Q�v����� J�T�	W\P�~�;b���6t�~�
q���(�s����[���2��x�r�̣�\r��T���ʝ�-��i�%��K��1
li^�3�3�]�zO�l�Me��_f�뇟3�T��!���m �o���}�����LB2�GJ����M<f�45W�����'� ��Td�e:){�vo!�~��4�\5�� 8*N���5VU�����x�-�C�x{��[���?`��];�����w<�ߗ��Bn��2f���`�x��ϟ,V �N����UyҰ��F���)u�6�E��Rp�^��9��D�K�L�ǀ�
nAo4�Ir�[�4aF��}�c�'���b�?t�����:N�%�a٦���EZ(^����X A��D\_)O��5=���duUW�ݘ��SaK�e��2#�O�1,x��O,q5�й#rl�a`Y�%Er<"��E����F�4�)���}�(u@�	���vw�iՏ%@n�q�	�Mau��o?��:R��q��4y�ɔ�n|K_ƹ��}������̧{������ *�;�yo��|\�2�q�lЗ�	<дBJ@�f/1�|�eat� ŋ���e(�Ә��P���+ '��-�,`34_���*�8��D�H��aY]�$qi�Nkɓ���,l(*h����cB\J���5O��jUW��Q�b�|�5}ȇ�9ѫ�&���(Lς��6Yxp�-b;P5�K����fz3�Q� ,�mO��;#��W�2@&��GEj-uf��OlQ��^�ԙ�4d�x+�&���ؽ��\f;���|U�I���$��n�;�\�����Pp#���%u��I�EJ�S(0(ޘ�����������Kk~&�L�t�p�V�M����b S��\�K$- ��x�IY�M��{Tɹ"���-��̚<:j���x-&��
1����cE5K�o8��h�C���K��ވ�}��*�k�.G��|�kX�OSg��9��F��dāF�o�IY��7l㙵����m�	�M;�l?&�@xX 3�l�<�jY�ʳ���xP�<���.{�dZ�pt��&�WM ������?��K�zS%o�ڤ�����C����F_�<��3��};����=@�E7`ӛ��5e��n��x%&�F�K�)dt|��0�j��``[a�:z����z�7�х�+�vr���y�(��V�^X�C�T��3b��9��##����
�7����;����a�����E��{$H/��R���'�U4��o�jΑ_�IΐZ�5]�[ӡm��c�7��] �����׮�}��BR�c�1j�7�ܛiH9�@Z�?�W$O��' �m$��<W?;���:tϬ�S{�,�kn9���Й�����Y暋4����^�cq�UJI�t�݇M����&U��0�����`��a3��ӿ	���-�
k;)yK&�!-H�x-�}�FB��������i����C�I�ɘ���c;��>���!�A۞�#�W��k<0�O�:6�c�X>6� ��7�p� �q�j}L�L2ӽ�TA%�OU�5+���g���a4G��*�j�����?����j�pڇ;}gq�
�^�x���:g��/�B���j4{�0�5���U��gK���T)X�K��ğ�-ܮ,eR����*���X�O�o*�Ҿ'��"3w���m~{*�u�^�.%T����Յ䦞�@����%�'�'��7n�(�.�LӜ��(ճ3va8��d9��↻����`TB7�ywX�L-%�k����ُ��VҢ��roAjfZ�~�;u��Aٺo�,+�m:(k��,*�eìl�KA�x�N����@�%н��:�<���I�~P�8����UqUt4D�f�‐
證�T�j`KT
�x��Ԍ��	9�fy�&����2g�A;r�p�3���c�-7����;)ҁ1�R��7�����8t�*�����ΦQ�YX�.�&\u5����@��ÀwW9�7A��f��6d��t	l<%J������4��XIixk��Q0.!3���[��(�%�uӲ�ͧ��$�^�n�}0����w�Mi�,��ق�w�i-!������nq'ֳ;y�,�#+�؏_Ԝ��L4Q��x7E �\!ʡƄA�=Jhu-��~���:���x0U9K���w4m����Ե��y
Ȁ�1�X���ӻ�,f=��2@0�"�rW<G0�Иt��m\!�~�� �%I>�%�)���5H�TСە�t0��B'��d��̤$�c�	����	���4��:�Y�ѭ�զ6�`�vBθО!	m�F՛���'ڻ��1�|�=2V������5R\y��A��Jͻr��T��5�Q�d+����_;��i�^�(Y��c��C%���e�S�� �"���ݽ|ҵ��F�!O�|���V�~���%r���)Prl)tå����*�]�T<m*���l�9��96�� �_��%r�:sC�V,����!���&�{$O$t/��.���Rk��]޶PӅ���g:Xj��dl�����Fq&=�A��ᒶ��v�Ԩ���nI�aYw����z��{��*�8��)�{��N�G��DH`Rj���3~���O%�n�oi1��+@Ӈ���=,��w6#�c����K�<2y�g��_@��:���d�M[>�p<���K��A#̲�Y?�����١/�_>۞��#U��+|�8�}�_�+)J J3W��A{��?�%E^|�)�w����x�FY��爉��7�JC)S�&H�C��	�7%c-ޚ�@��XH���J�U��L��wO߫O���uX2����v�V"��9.'�X�_��5��2 w���hj�y�{>��8���O3�8��n]�S/!d�`ڈǀF6���tVҾ���ֱO�x���ٻˮ�@�vc����\~�=��ݖ��j?��܏-���o`�[��{	�9�h%v4$�F�T�~׶��^n^�DT�u��yNx"|�P��T/�B�:.޲JÊ�	](m+����ü����;��䕺/rr�+���o<�{+���t��uMl��ٸxQ*�n�/
U�WV&J���p�|>^ݺ,�%<�r#hZ��F��u���2���b���+����~9�o][�w�n�췇3��dk�k8W5k�*J�6\���\�v����b��46����t��b݈3���.�A�:��T�8o�zK 2���?BJ�ލ�U�1�t@��Q��vף�7�[��Hc�R��o�����D����=��s�҂�^^T�M�N�|�Ә^����2�/E�o&zKAxR�8
¢H� ��i�����x���4s���h��{�w���6DXwc�g���ɬ�)�%t��%�	r���B ߱����]\@�.k1�t�`��{����7�{��Ϳ��uEY�}�Uq�C�d�z����7'��fçib�j�����1�E�u��W�_�L�-��_þ��w߆���	1�Zne�۲�Wt%�>�F�����p������D\f��K&�[�l~��C�2Ҵ��3�/b��qQ�:���\����:|P]�F.ݑH�j�
'��׾�Z��ހ���ֶ�߱qn� c��}���$ފH�̪���%tq�}���@���!�%}`��e@��i��χ��q���YoW4��ȣc��^J�;�:V��l�B$iPH2�%�D	���Qt�@!}g�&Axv|3M?�^~bNʫ#n�r
�\����D���}�2�������mu��&����匷F ҿ���>f�A��^���+�m��L���Ӯ��R@��껲����H=܋��lq!=*|�V ,9�G+��`���%,��U�Ӫ�]�d�����nX��6�p��#d��	ȚP6������{�|�͚م([�c�ц�>3.0�Z/�?�2�ƽ�����b���})���=v}���Fx&�(�܃:E�/����AdbgԲ��5*H)��g��lw��js��ofJ���׋�T093a�;�rP�wu���T�t��f�s�e�>�`�!c$����߉5��*	��Kd^Đꧩَ�점�^�%mML�Х�*mx�)?� ����&�٩��QRS��C��5�
LO���A���7Qn�7�U�Uf`zJ�����γ���Ό'`�Q��T���Q�\۟u�}.�ump,�a�̈́�gÉ�A⢼t(�0�IS\<^�V�����!d'�.�n�ɏ�����~�d��2K��1�p��:�ւ�+f�<��Ė6���*�699���@+>*r�7.	O��P��D��aא~S��	���~�mop2D�����?@{�;%f��6?λ���K�E��1�{鋓�a~'��6�S`�x�0z
.C���ɿ���͋�$�`v'1�� f�8�(n�H!��݃�Y� 6�J��l=W��^���QX$�fЃJ!�G�9H�j,P�M�b�:�D&��W��YU�� �JcƝ>0�w�@s�|E�Źq�e���[�
N�,��k�/w��'>���ĳq�Z��X�����%��a��?�:+.�"��'³P�d&=מ�Z�<V���9zc;�pe�_�"�]5/���)
*������)�g�6�Ћ���+��c��ͷ|�F]x�b��XT�=	 �
[r�*\`Zq:^^��x���^ +�wZ{:ΑAJ@6�������]	W��V����B�m�_��a���	^���
ך4`�Q����mM>vs9j E�y'w�G0<��GǶ�ŊQ���P|�p��'m��s��bO[-e'���%��֤ƪ@�Y�rv
9� ��<!�y�REdq�QJ���nEzס�H2f	�W�{��ϊ	�=ȉf�Db~|׀0������<�����5
{k�W��F��J�`�=Y2�k(.��X���Y���!f�l��e��N.S,�PAGhx&�����M�|�_6��顟�55�ou��T#���-~U�}Ħ��L�� ��=��t��J����}� �-��\;��F��������꬧]OM.��P�J؇�)�ڝ��	_�4w��/!���smپ��Ѣ�j`�G�1�B�P�[�ٴ�į�+��w�M]���E�vM��nL���[��Ն��QEJѷ��ue}\p�zu>�~�k��iH�N�}T�ez���YS�_���m�̍t��Z!)�X�xԦ��F݂���8�����*;6�%�f�G�<�pGO��sդ��,>�T���ǲ�!�>8�:1:0�g_PpdZ�S(kb�_t�����_����
��Ϸ�[��#����r�djL�O|��ŋ��K	������>?�-�m8ܪʀ�:��7��o�\G�?�}I�Q� i��u�,qZb�Qm'�=�F��L�P[2>���; �z/��3�c��1MԐy��:�:ǎ[-N����h)2����ݗ�?���1� �5"�����)�эP��|_��Xx��O� "';�܎��yg�QUx��sf1)�u���Yh^��t6����ѝ��aC���qm�Ro�D�M�_l�� �A6�� ��N��W��E�1��2�*�`U^)�Z�>xxŎC�3	��!W�〄�׸�a+L�OB/P�����<+����o;a28����B�cr밐L��z��h�.��"��E.��8]/�˜<�|Q3��[��L��Sh"�g����D���z(�kި(d�ǹO
7YD�k5��ڶ:
�T)���Ȕ'T�� �R�-���5,zh��g	�PN�IP�4>�Ҝ$̸����'b�!Z���̳SZH�g�`MqU6�χ���4V		Q,�󇓥Na	)�V;���4�\,z��ԏ(`����y��&" i3�f���z�I��)��0�8H6/
i�h�x�}s����lDR��Xu��5���(��~��?�O)����a[�W���2k�7��K&G�3g���'�e�b$q��E��&?
c�������Z=��t����9�V4����A��Y,/Mȟ�U[u��׌{�ʾ�G�Kj ��
�X����=0~ly6X@�����_���K���o���Y�����Ms��fe��ĕin#k�^XZV�5��� 8��]�8�[�\Ѕ4=�BA�Z���'-�i�r��S����+�^^`���Al��o-�<��\]�iL�H��T�B��S�4,�{�d��?@&�^qÈ_CwT�:��|�X7(�<�������x�V�Ne��Ԋ8Я�¥��6��^���Vo��H���I�6�F���K�1#sF�_�~� Ӳh|�Xښ�S�G��ӧ�:?y��LO����ɾ|�`�!	�R�}G���f�<GH8R��!K�0�5�&�#�_5V��� �:��io�15m�>�,c|;~
cYoA[e��k�a��s����[�Ҭ�L�/5fL퉡3�_.��{S��ˊ�	�\�G�� !�[��eQ�ٸdB`�Nr�J�2�sJ�<uU�G��Z���L�Nq6��8�,�K�OZ(5*�
���+��$�A �TE���RL˰�,22�v=�lO�!�0q�P��W��b�R��8.;���'&�ٛ����-�|�c��ȹ�.��0>LТtl +�0S���u{�r�?OH�@�!5��#m!|Ky6���÷/�_7��̜��pV�)e�gƜ���̀��A�o�B~�^�<դԹ��fG���]Q)M���p�5P��nC�2�4E���M�aDa�t���8�G�`W��B��n��:�?�R�����S��+�C�Kyb� ��U��\�.o�ґ->�]b�~18��+��TѾϟ�v��^c.��C�@�M	-w��#��1�rTa�\A����+� �q�ݻ{�Iu���7���X�ND4;���)ߊ��Y��s�`�Ԙ&,�r�� ��������}�i�YZ�k�W@��K�'+��Gi1��,Q�
��h�W�S��� �D�%$"`��*��?�iܱ5��zS�9_���7Q�fOj R��`>�<�ʫh�c���u���(Rp��L�rD�׿�a���)���  ��<A���s����KM�� �d�7&��}�Y��1���)���Иm��Y�}5���B��9�g�Zب&h��6 ����KW8�,�s��j��>7^V���C�P� �s�v_3:���!Ը/v"��z�����>��]g����g9�Y�e@E���we9���%�|�D�ͦ�%���t�V��VN�kpf�f�e"�S{0q^�(D4pN��c1��˧��-��{�T��oܠ��&���Z�-�
�/�Ă��y��)~r��ͭ�ظ,*Y�L3���$:���ˎ���*B.����ۓ^�,��oPS�� K����,�s�N�O����=U7�����	�L_�]
��	��ϑ��gKD*���&�SU�̭�]�D�^�l?�5`Q����]�u���ݘ\� @��O:^�wS��F���SrG?�9-��x���Q�a%�'l��8�|W�9����AHN��đ�"���?t��HL��Q�'��d.ͥ����0�ݴ�9y���=m%$��8*T�+
�K���d��hV�(E&K���lR�l�n���iw�G�'��&��%�yx��Rx���ۗ���i��G�!�ڭ~�p���>�ڬ�({ʠ�q|���T��*1W6����Do�0���켆�GH�/p�ub����L#�$_�J�(~��/��o؃��8:Nw��S�^a.]3p8+�w�ݤ�}pyOY[R�c��+��wrN8_4���۸��+��(,q���y�� �}�	[�U��=�4�� [rGN�=�xF�;��MS���sZIɦ�
r�so��6�0�Yh,��A;�~2�!7���[=yZ�cC�5�T�����J-� ��>p+�p��wu�˛<��q��l��4���F���|@��HLR���������e���(ٗD;bm?x�Yui؊X�?�GŨ*�W�H���[�\��w�}�;f�׺��1��*�KS�-��~j�/���,�8yĳ��X�b$��ܙ��ˉN�xP��>3�� ���е�N�����3�����( &�h��1�a�}
��<7��5d'y�nu�9�,\��%;5!���A���:$p!d^q)��,�Z"�_��hb�Yءm��y�tfP+���7"9}G��qN��+=���b��jI͑��=/	K>�{8��R%J�t�:�g�e����t�1!���F��f�X�����WFV-�V��b^��]��E:��;g�r���'�*� 8��)�������C��d�tb��9_'��������2Z8_aj�%~��"��TFe�w��)hMB2�^R���]�0��2�2�~�,��Z���H��'�5F�犩+K�R�l_$"2\;�T� 9�>�͂�W�G#�ʾ�ߪc���[Tn���)2[���&�2�4)�%���F>z�k��}��9�$�����)��mW<_����� ��Z�<)�11}������l���o&�h/�	sa���F6Ez)fjx��������^�~�?hq�*�h�&��gw~���h�'�K�ս:Z� ~D����)��lU�N����!T�TlD�K4O4�p�����J�9�j����?��4�Ύ����t�)O{� v��~�����S6�xs���6f�U��զyt�.@�2���<�9�~��wډ�%�0Im������{��ބ��g. ����N0��,�v:���4��8LV����U"��"��^�L% ��<�B*W��������3���z��=_?z3�� 
|%f�L��g���Fų�����`�"L��}j�Ux'SRR�7������%#ng������[)8�2�H�}�<�D���א� %���u��$lݎQٶ2���x�X�Gy�M%�}k����jRF�uCrC�⬴�S�iٶS�7�
�1�t�ϭ��y��A���W�;�U�hM�eV�j��f2����k-)vI�����S6��
FOv}��IjoW�6�"4��RR��BR�:a�9��|��i��3R�n��I��6�b�R��2�":�(fn���O*"G�r��9��&X�:�s���ck�rz���Sw���R�w����֔ݯ̤�^C3h����q��z솿���e�]�<0e�C�Ʋb�wQnG���cy�tB�5�!� �T�#���'��@�IN�C�|h�QY<o����%'��QkT�ZC7=yvB������S2��/1T�|㑎�ץ_�n4�/�jî����V���^���7:���`�ǚM:>%��?! )d*��`������̀�& 2��{�9���o�k���9N�D#Zo\JXD=	����chU��#�y���Ӗ��ŷ]� ��H������c��{��N�z�E��M`�����?�.M�s����,=F��Q`n"�f��e#��8 �X��J�5�x9�۲��K��h�U]W�H���/Э ��\�6KF�{���a4+N�.I�EsJ�k[u�$��|�5��-�q%�xZJ�Z���<�>���K|��lUM�yd�Ƒ�e&6ұ��
db�l�v=�|�~������*1�f���a�K���c<헋U6'U���A���Y����\�5����.W��	''�>���<��D��\S��A�z�.t�<)��� �g`��S�4T���m�^��Vmk$r�k6(-�2j)��yFS�2T��a�4��a�:y�Ć�wD�&9�A;� FڨP��Mi�)��E0�ƀ�I�U���J]Kk_�٠'3���q�8�����B���ʓS���5�K�jP
�� ��?#��= �����JA�(���ӏ�O�%�&?,`<��I� �)���9�8Ue6�
�+p��+Z+")��
����t4�2z��_��/e�r�|�A9���B��� ��Da�J%,���W�k� �=˨9�r�e��Q@��2��|5�	�s,��On,L>a�İ�C���o�u�qɝ+͑8
����X� ʍ{�,!C�Ґql�K�aP��r�ZV�O����@i����@ �%�IS�JtZK���� �R�l�䍩r�k ���}[��Y�`��\�(�kX��<~V�lFB����)��<H�CǊ�PN|�'^�GԾ���%�Hۮ�.Ҩ�aFX[�?
��D	��[���ڋ��-Mo�%�|=c��;�{>(<�IG<�.د�u��ݟ�"�x+�sr,H/��Fe��N�) �Gn.�����x�8�1�M��mèk�ڝ2ct���'�����/�z<����� o��*�8#�F/r]?OL�Z2�z+����S��HJQy����̵N`A���B����ꐥ[9���sƚ=���� _qV�|>��BU���?�����w=����� -�$�ด��DW�&�V�� 9���P]�x��^�B��S)�_-�h2����9z��k�	SiB���<1w�0l\;��N����Q��t��P%؟"���u�CVl���a����iP\fZ�1}`R7�v^քdK������&��F��h��|�1!�#Q`����֭�v��<���(BhܼS[�#�L<�:!�Cx D2}�a�G�kQyH�s��l��PV�xqd(���m���@zYY�a�Qy�|�i�OUC��������b�j�z�e
8l<{�-]�yi�_�� �U/��j-�����;�z��"8��a��$G�����c0�V�J�1c�}{+�퉒���0�	���kT�����;]�9Jk�&�Pz�ş��\u ���QSA���KJ�!(�_IT�)m��W����V� ۮ��Xu�Cv�$l|4��B3��n�S���w���
4�XtC	/��,q:CO�|n���e������`Cn5���ў�["���w/�X��Sw�8�i�r��#W�N����q�-sR9��b�����Ɓ�%�f@b��w���u�⬼4��Nb-E��H&a�i���>z����{n�c�>�����0��Z���F�n��*�~��x�)^e[9�t�D�Y	�P�<����?ŗ�)\���Iu�_��4�j9�+>4�Ś��>�Z�<d�~ٓ��C�r`�pL�T�u(���Շ��k��`ޭ[���ʘ��"̹$o`�޴}0K�Q���a�6<��b��=~*t�v�+���$�g�#a_�d6Gz>t:��of�oQ�<��m�헴��ŝ����	�*���חr�?\�%�G�Q�-o��̬�s^U�of��yH.�P��[1�M��������H�����N��| �W�ևu~C0�wG��]WM�נ�@,��;�H��Z�f�!t�߂4<�Q7�|�-n�?Y����I~K���!�L��"qc��Fʣ1��)�r��5x�;�]a��b}Ȯ�-sd[z�ǉ�so^Y�t ;�Z�U^�?�<�(J�����w�<���UZd���Q!x��9���f�s\�T���I4o�Aک(�����ˁ+7�?T1C���4��/�{�jw���CYQ�{�^l�Љ*�w��(e�I?VE��k�Uo�&������wZb�E�/(|J���cBY��S�ŕ�H�5a�"�>�G +k����G��A��o�W�����3{��=z�,Ӛ�]�K�od���c�_�H�N�q�x����hH�"H��jE5��sa�n�?�Ť�#��/��p*,z���zԡ7qc,����Xlܖ���5o��`<�u �!�����&%@�z�]zTW��-�U�Ε�}�@H6� Sbɪ�����-��R>���C�]�P���w�5;��VZ�ȕ�D��6$�Ez\����-�� �|�O����o�пUU��!�F��21��|�5��w�~��QAEŘ�K�U�DTe�6C�A#4�� c�l�J��eW�\%�P|�sMc�Fto^?]�:GVu�E�e�D�>�?H�ū	~9
?ׅ�����?'\�*8sF���uK��I�wJ3������@�F�%����4�����������q�
�5�8�چ�� �ɞ��Zz�u�z��j[&��w��7
a0��{��?N	�C��������\]�@�P�O���}���Y�q�j��b ���E�~
���B)+�ҿH�z`Jx��Q,�K@,�-K�S�g>����֫����">Wb�vr�-C?p�t[�#@>�&��E|�ܻ.�9`����=����O_�+ǵ�g��-�)-ޠs3�N��./������@O�t{V����rB+w�=� 6Ȕ%�f�uxc�,~
�RFbv{��k���1]��-�K�_q�c�į��ϼi��^���:�9Z�!�~ᴾŻt� 5`U`:w�&w�3�ZR`[�zD>-�݆�}�襅7�+p )��}�}�R��'bΌ\<{+k���w�H x��C_�4֗E�O���`TZ�b856M��!<;4EkG��So��N�©�:�9�︭�kSA���N}��!�ڞ��6����{o��6C�G�ٺ�B�����eK�����8E����E�g�h�q��&�z���e+��Q-;���?�L�MĒ���xDsz'7?+�RP������#��ƈ+�	P�a&i~Ƞg��p�=94��������*�f
~�;�N!3:e�Ń�Z���9�Ӿ��	��H�-�C�kN�N� SL�B�~e�H��	��L�%�il�\��J;x!��1�$� V�JWRhg���՛����ӂ�R�z�;5�虳����x^Z0?5G�s��(�?t�yVoiN�i/;y�a4L�c����py�������o�p@�=[��0�	3�LNX;<�1��L�	�	�g{���+CL:5������L��`��H4kj.�wK:@�@��`T�B'�~w�X�TW�j.��$Y5Q@|3�'/��b��S-i)�N�
�Y����t�~����i�� �5�^ڭ�T-��Pńq�3RQ1���A�aj��R!Ʃh�˩��w�נΆ4�.@2��\��n�P_�ru'��ɂ!Qn��]���:�_G��7I���V����������X;hev!�S�&����tW��~�k��M	I�7��z��L&��0�8��,#hd��5�&	�
TE�|�=��~�_�f�T�3Kd�BŒ'տ�%��gzbؐ��3z�9=E,�\ɴ�E���,��g��}=�[�9H^Z��Ͽw�Nȫ���<�K����#"�F���:��?��Ԓ�G�C�!�q[Ӥ�a���� ��[�T��#4X����}�=5bb6��V�X�~S���Qk��(�8�8�W��n�n���Qy.m�S���%Z@��ϣp�CW�n@.�1�	]@�5�>�u���0'�����3}vh(2/��R�U���{�m�'@���q���6�]?��Nx}ν��M[�Щ����A� F���ƖJ���f��	ٓ�J��"h���=	d6�(��G����͑#ٛ��-�C�堳���Sd�E�C8
�%SlgNV��d����|��k%18s�z�5ؘ�&α���X���w�G�OFf��Y�!�^����հ�^�H��ɷ����0�����},��p����וc�e��!S_\��Y�y<V�T6<�8l���.��p���]�E�f��
S��A@5Q7|{���*��5�*m��x�mxM�i��6K��crg��]��8���-{P�隊`e63o@���ٲ0�E�3��}Caö�Q÷��d�iɫ��D�K)�����F�	ghC�.�����`�� ��h��鎙X��
u�o^i��PʈQ3���{���d,簸�S�ށ��}�rT��v����?�ٶu�G���x>��􌄫>H��y����?tV�ͽ�k3t�*ǡ|�W����m�V�>f��"��6V�˗�B�b����T^�^ejc��t&�24�^G�_XKr)�EЁ�PTn`��hl��;��`i���Dѥ��\��j{0��dn��-�J|ś�˛�@*�5�aο[V'n�43�����6��rL>�"�"
U��F��_^v��G�u������ĕ^������Z�@�˝"�	�-�p7��:��������>�)���g��w��07h�Z�PW�� �б��RC�q��砙E�
%�g��:)�hFJꭴ�M��P�5�ø�"��e�\� Ƽ^��wz��_*(��/e��:xȭ[�J�9�5�'Ms�E%������TC|��zUyǕ�q;�n¢غ,K���Y�+�~}"5N{Y��Ah��|�F��~-3@+���UT�b���-{����{+��=*�o��>�������5�wv�fCq%j��p֫F�03k UZ�b���ѨwG���Q����\�p�aPDv˚��������5V�g�\^M0��QG� ����5��s��j������]+��V-:���L��R�Kw��H�KMz���N"h���<XCf/����3fd&���X�}�����L ����!�h9%Z��{�dav�T}�.C+�W�])�y���"�1��/֞u�D�L<�y V���9c���}�R�R1�.� �A8�Gvк1>	X�b�ݘ�H�SBU�o}m,͡�`-0cUT�X� ���,�C����j��u8X�d5"�o��ٯN�\���.���Di�
SQ�$�=fN
����x;IK�#"����|���j���2%�|q�y�˪"����Z&jS�'g�_q��(-�h�>7*���l'�D�3��"kdf���j+jL�
��9�7!KP�&`����E�J�8�tc]ϚQ�W� ��+�!���=u:�V'Sd��mitDj��p=����0���v]�������=�#���T��?7S�9��K� cR�
�te�����b6Xu�İ�cB����_d�˺"I���p�=6�W�4(�9���[e����^2���S�t���B�(z}�-���$�� YVT{�)Ҧ'�R2�/�}j�K����T����Y�>��o��`�g���"��������	BC*����S�m{�Ű���:<u+�0�rV��	�����r4�ĉ���)p���-�F�}tʭn�:�b#�k�oB�}q�.��`C��QdkF/���M��s���0�f�\�4&G�����{.X$k��dm�C���k9��ZJ�SW�t����������	d��
X�:<���	�@�|@�������=�����\*���	�K+�K��Uß �*���hg��_S��=9�Q���3\��z����.���Ǔ�Q(Fi�Y_c,�S^4�l�Лu�BRhF5km�c댄��hc؂2����;`(�1u�@�C��������Y�Hh�U����]�#�d���?�+�S��t�fM���u̓oϬ��#w�F;�ه���K��Q�%�l�=z?�ꏕ�쮮�'��v����nT���S����^@=C�y��֝��,N3&����f�oV�"�|�a�;k�慡��nf�ԷH��V�s�>�K8p8�ܝm1����1��<�;�!�MNH/����b ���U�i0��Z�	�n���NLe5�h~��e��L�<��E�'��HM
D�o�n�U����y��Z�7�]�&o�e7.o�%e�B?�4�?+�Լ�C7�#���Z�}�5�������I�����69�
�k���K�Or����y4�
.:����*��ߨ���ix�S������9X)����f�B�o�-���vx�[��_17��KF� ��@��k�3xn-@ɇ�=|ɰ�G�^�4V[�/�>(q�:�����	F���KR��!�U�p1J�ϫq��Y���3�jQ":�ӯxw͘)X;9V���i�����x��Nao�^�Ҳ�
�)�OC4��� ߋ�q��i��r�U�@S�z1ؕ�㤟���sQ����y�ن��+\�yŨ�<6��1�꺐5R��F\a����Ln��ɋ57XV������0;�F��Ɣ�������1h�����ݲ������`��p������>��0F�w��z/0E�u9��@�}�R���0ެyp=X�ci�� �C�]_�Ǖ4�ߏ �!9��"����p	\�8���Ǿ��76�T���p$�#����jؕ+�b����	��l���5�\���W�	&�!��>� 9cs5���5�@� �V��d9��Yh�x<�1{҂�-�Y��#2����T�H.����$P�b�Ⅹ��� )3�Ϫ��<��\'����^O|1���D~K�N��X�XK�pwi�wg_�����I��?.����u�[̉&y˰&�$�ƒ�f��i�f,1���2r���?Wӽ�ބ_����Z ���3��n+�د�<~������+��	RK�x�o���|���T2p�e��9�������?a��b=�Itk9ݤ��'
���n� �I{�N�_`��U:��]x$rE��P��
��X6�>��j�N�٢GwO�ܨ�vh��mWL�~��3@���������K�,�8���#��]M俹5n����m�E�~�d�T����}��/�z�Ѽ�>���G�gx�y�����|f��g�5��K�R���/�4%�>l��5�t�;�.��/������}�ڐ��I������ݍԋ9�pA�<E��
˟(�
�"@/75_�cL�X���:5f�2�B���� ������4Z��ĸ��!�6��b�2�	�}w����0]Hv���=8��}����Y�gu�%�"_yZߐ���^��OU��tV��f	��f��@�>{*�x�BKƔ||��L����`syw�����
�{�/����:f��s���ҡ�o�����1#U0�e�C�b�V�8��5m`Gy��E����0|:�\��u�Ym� >����q�f��oJ��`�Ab{E�T)�6����ow�>�K�}��� X$��z�֏8EL�I�֯��xuTr��k�NYa��Wt�,�>�T5;=�k^���u��)��i�iw�zA�w�&js����k�9�Ү�EyF���-��oF����&o5+
�t�0P���7_��9��*鰦Yߜ�^�K,��u4^(�}jN��(@H>Y��J��:�ؚ���Hl�QW��J�}RNO�� �[�T@|udB��iD�8d�܍���#����!�ӏg �A�*j��57i⒇^ҵ؅��߬��W^��{��䫢rN1�d�3��&�0�� K!����-`�QB�e�����?�G�yz�\-�n+*;cC��]�Bw���o���U�jrE�E�©$w&L�K?��sݩv�	N7��`��d�*�Xr�9�C/��uX7]s>���������H^����_˫�����nIѱ*�4���M�%^�q�b��P��Y9g�1�-�n�!�5�a^��ԗe�y�G_����t���v��p`r��H�$�O
+�Ơ��|q�X̕�\yC�}޽�t�������m�;�R�W���Z%����4?��:He�m�.���"��%�k�Rײ�H�^�������[
)9��ϚB��9�����k���R=�L����Z�.lpOU=���iI覗&�̷'r꬛����Ȇj�Ey�}��e�8�W����MS7��G�n�$CZ8jXRE�*ݟ�'j�S������W�:E<�l�uc6�ܱ-y`8h�|�]��Ra��?3U	.��UL�e=3tp�j_���5bL����%w'~�9� ɰ$~fp ��P���/�N��Y#���w�Ҫh�^�t�&�(;����>q���-i����|���8Ȋ�4��%|z�����xJ{�T����OL��Tx�,��&:QR����z����)����5s��ڦ�P��2z=f��Qu�KI-��M�a��Q���%C�P��DiɄ���il��{l���n�6L:^���@�X�Q	'c�=�g�!DN����	�����r�㎽���ε_7R���&f��eSh��`���t)̸G2%��sp��nN��	uȹ�r6~V��۲��\mKN:���zP�Fz��A1��I�G�;��w������j�@�}�G�V����0f�c�s���R������� �p5y(\��*+х�C�OX����(�b�����o���P[\j�",�vh%�ʚ��2pKK����3W*Ef:�B��=R�9E���_"̧���h��l7���' ��|��wf�b���u�u.а����I�F�<o;SWD���m�E<0�Srx�ޣ�����YJ/�Х��5:��\��\O=���i�9������[���z�s�b�v��@�xs� ǂD%7�+'H�j+k)<
�UE(>dM�O�n�NA/ߨIT�a8�s�|g�Yaÿ��)���ʈx�4f����Oz���\O���C��޸�l���H�V;�/�3��(,�+�ނX��p����F�B���-����\�Ьc�Ym��mOr��O�@m
�����E���"4��+����]�djg��'��
{Ӧ2����&c��c�~s��`�����y���Oܼ�3T������ș�jL��8(�q0�<�h�d���ro�ol9�"�>�?����LZ9H�?w[)��!ٚ��A�ܹ�3��oB��%h��f	~<	�"J�?(�3�6����5�s��|�9�������Uښ��@�8sDq���q���M<D����t����L�Ӆ;Ȼ�b}e
2��PL?
��)��N�̝��˗�'��%=R� 2/\W<�=�b���x�;��cP񥅶��� h��9C�1/TXX�����!��jx�@ �����
���ձ�6�"p_{�����틷�Ʃo�������Cm�� ��`+@Ζvr�����XF� �ݙ�ͣ���*�Ӏ�R�׻�kuE0[z��+�k������-c��1-�������u��P�u���!ΤP�`�&�_��X!��s�C2��k�}u��P��!���%�^����J%�d��f�|T\R��7���@XVʲ�FCʥ�� ���͢���B�S�̓�b����{:g%�;
I,��1~A�z!|���	�<�3~��`�(�N����.Χ��PE��G�N�0���O���R��/f"_�a�3���k�y1�wSc����2�A�ܻ	��A�O�?a�(x����@N}Wi�<q�������n�߄N����"�ԶE�q��b�'�l8sW2/��ޠ�ej���B�K�
9�F @�s���H�ɗd$溶Z6נc/��B��N��ņ���9+�L��'&� S���]�) �� T>��Z�z����P���K�5:x��y��>n^ن*IC�kʼÁ;��+�'����ߨ��H�Y���`bd�g����`��|tĠN��L6G�K<z���\V�<mR��#){��͉�Y��rKг�ke����+�� �Ҋ��q8Z�NE��
0�VF>%��Nd�7�����osND��\Ca�����#�Ocoσ�_)�9�@�s�"]�g�ȐG�V��V��kV��u�m�R?�^����"�IZ�W|%W���gJ,��ܺ?(�;oG %�l�p���'��N)������ E�<M���2�Q��0J��Ґ3ז{
^V���7m�=�t-�T�dz��C,��X��hy��L��r[�2���)�"�ٯ����<.q��
9>i�g�a�Y�.��?�Ux4����LIe㠾E��䤍#�?'�/�"����/Y!⋬�sr4rN��ǎ��^ <���@���-��/��	1M?�����XDSKޒU��J��`^�o.��R�g�{���6/:^��K��;`�X��o^-�
�H�5����������߿s8f�E|�a���lsh��"ą�F:n���n(*���Z��yX�Y\ܥ��9������|�P�#�(F���_�����$��ԁ�ȥ�y{����2�Z=y�Pn�pJ���'�1�A075��#aJ����'���IL=	 W<ݟ��/;\�=�Rn�z/��>���?4�i�Q��LU��`lT  �Ylt�*�ٜG����\+�4�i�����9%/���v�I�;��DV�5�J%����	-�6+�!;��{��K_	F;[�n)�s��}M�\{�]���+�tE�v����Ws��M`3�#S�$�~���_�~طD��փ����'�����^��~�R��#?[Ljij���O�֒��hH��44���!c)1�w&j��8����\��.�%0c�V
Ȧ�؍p\�G�����.��qG�C�������Z��l�����A�o]�5�6RN���^9lY�XK�f?�G���̖�1��<��-U��?�]p"f�O�^�<S����^���|g����ʕ`��__�ѳ���|�	�<�;����-Pi��C��0[�G�у	�P�/�S�� M\��
�Wa�����Õb.�B)��6�
�EOoh���������"���G!%h��%X���L�K��#N�}�y��x���o�趟�܉�>�2&����#fPu]�g��b7ڱ������Jl��>�b;�A�e�hw�!�&���ӡ��� ���(���=m�����iT��8U� 花i"�8	���c�����H��:��9�� tn�M8��bS���Gd��}Z���P�k��O.
��ri*�p%��GB����5�`V����pH𓄭h��[B�zLȦ�"������6P��5?�zg�����=���8��_�O����!�|!��X��SO�ޮ%��������
1�{!-�73��uyo�v��!�CY������BrC�V�:���<��l_\fi�lk 9A[rX�iQ9�ㄿ�J�j��5!�ւճ��&�쮫*�>��5ڙw/�f�pw�߷t��3�����:+!>e�iY�ϐ�v��_���>�T{���#|�����m�O�K
H��_e�(��HRx�p��_Њw�O�tMV�o5=�)�5}�~��E��#�.t�_i33t8ö��Aǽ���R/e��܄_q+�o��*�AXF��löم��{�UK�K`+3��ު��r��(�E���'�)��E;�'��q"݄GX�Rk�j��G���Y%�|d��՞2���XD��6��՘�4�Z"��k� 
�6�F4k��d����0Bv��2��O�۟3K[�8���I�VF�%:e+�ńJ���tC{��
�=�\~�C��;�*��O3ù�K�kj���P���AU��dA��#d�}��*{ǵ�5:{<�5�B_=�ױ�|H�����㤳lM����� L�nH�U&�,���$�am?��x3c4��tUC&���l"�tNRb#�G>v�q���
�,䴌�zJqm��&�i�T�VZ8���UL1=Di1Z��n�͒��T�^��
���[Iyz��8�Dt ���r�+R�������Df�G�͉=�t�3-~�oV�m��]f�%�L����˝�r��x���J��A��IW{`�K�!.���J�&�2��X�F�O�����-�����3}!�)\�E�܏���YN��u�T�!�0��ͥ�΂6��5�jr��PF�ۈ�d�0��X�-	�?��}L�]Q7��|-��{������e��]9�8oM�ѐ�����&��t�=cm�"Y�-�� @���BRz{;λc�5o����o�C�(��%ϋ^��몜�W6�Pu�Tf���r����q��n����tҰzzQ��r�� ��oT�M��K˸����<)RORG;��o��?�W�������!�IP�	����.�B�Ϳta��h(���x[��G��ttDK~i�ّg0�&l�k�T Z�uXҰ��8�{�@��3x=<�#�.i���'������)�؉)��y6�+;�;��J�ܨE�����9���-7�d�p��I��n�zjӮ��:��
��	�楪��k{���a�7)�������Xs��ҙ�W��[�Ӕ��IX��-ׇ�=d���f)N~@QU�v2� `�*fS ͺ�/k�Vr"�0,E��.�/��xQu��"i#Hy_�]�,�dqۅ�E:iGhA�w���g	
�d5��P��z}L�Iٛ\
ң�;ȪV��wT���N҄,%-)=%|�P�g����a�+�����ײ�Dj�s��,���u�����-F$�܄EH��W������M�A����iD-ǿ%)FT{���ނ8�����>D4T�|&k}�0έ��B�w�}?�kה�s����~7�{63����ɝ�I���f�Ś62Տ6j�y������L�O������2��M�J�?�J�0��7�s.1�{=v��KuC`q���<���֫{b�þ��`��Ow�:w���|f	���%�$�J�"F�4�r�8�2Q8�����m➷	� u�$��Y6�̬V-f�V"x��4��R�[Y����}��TZ�F�x��OX�
��:1]���lP�����(���第�l~�#vAc���IO´%$4���y�s$gk@CN�vj�y�8A�4���$��tR�0��ߢ�#������H4��5�M�R8�
u����Zlg�ѝM�,��w,�� Q���=��,��T��w��r����P�����-�xE|k�f���xM��������:OY#��Rq���A�� ؊t��"�;Sp��=B-aN��M�����|��Ǐl�!{lm�D}!�����<A��>WA�eS4"�J>JJ1v��Ά�0�b�v�8��}h�L&�kDcn�dd-���Y�3+��wFy�4呝]O�7i�?���h;G����T鬪�(���A��B/��v���:O�6I�߁ b�g�u�S۽�����ea��.
e���6Z	�}������$�"�:�f+)��p�f�N ��v�����h�}j�h���(�S�9�pm�ǞXy��h��!�I��H*���RԸk0��2i<9�0m��Q.F��&b��dw��ئI�����D�wp_<ا�e�o�����
e�
���Wa'��C�����������n�cF��!ʣU@��oOqb Qkt�.��]eNPF
�$�d���b~&���֩,D�o�0z8��$���'��T�ެ�)�a�eۊb0��35���~J&N�.��ꘃ$l/`9���߳��MZ^U�d�����#� �BT�vy�Pڴ��He��O_wq��]�U��eVH�����i_�{.d�W|[��0_l{�.eU'�#^.�?�"�u�c���&p���O�`q��5�ڸ3��|nE���A~����w!��5oh��x�!qib���qb��������,�� ��Ni����0{�hx-�^�ռ@�D��oj#�A?U
S�Z�*��@�>S���^5:/\z����ڭ���Y�$ �k��o�=��ڀ�����;�|GH��-$_� ����-k\��R�Xt��mzM��n6�����0��_���bƮw�
�2��&��̅��	�X��Xv�v�ݟqHv�����&g�������.-О��':(�`�F'E��4�]"�"π�Ф]�
I�Q���;[���Xa'�M�=V������e��6��r	S��	����:8��8P"'T���(�J�����s���(��ِ���N����'LA쥃���*9���?�;�R�k��I�������jHP�"�W4�)`�g8�hXn]ü�^��6}�� ]5!�w���iԓZ�;�nas9P<З `�r9Y"$)�9c�f�ޡ=$�<p��	��.Ў��&�9]����L=���B�>��.f臽Gmc��mh̐�V&��T7�|j��p?)I�E��r{���� )�h����<��H�R�.��G{N�+����b@g�9Wt$ulݠP=��X����Q�"�\t�jP�R��m�Q���7��N�*1�&�2�;�f��k/�g&�zo�A�Ik�!��hTg���m�9���m�Bt����C�:鱢��N��1�_���I���b㏻�?�F� ls�B�Re�8���Y�"�y���_��F����d6Xcּ��\ �Ҹj��@-'��佦vٚ8�1���J
�����)��9�<���:��~�����t���`�"��}�~������V�A�Q�S]�X"mGW�����wx���IIH��\��� �D�_P���^�{Gl�$�J�^֥��!��N��)|�B��*B]+	�?~��
�h��=~�
������ݐ]���zn��-d�6.Z͵M!X/z����	g���)砕��c����7[|�����p��@�~����4�?���@�v��des��-&n�U�Xp���W茛���^�h�3QظB.�A%� I����ۺ$�J�U#��6��_�,m�^�Z����:+�mf���VFZo��f���43���H���s�c�P��s�Ӌ��'a��
CD�N�zIҝ�cK����[��x�����}
�q.Ucu8���;t-3;|�K~X����>��ja��zP��i�-��w�w�f㪋r����k�3͓AT i3s�s���6T�f7k���Uc����7��NM��M~z���`��rEj'� ]���K�f"�Q�m;e���@��8��oeX�5�{�3�'��ݖ�.��p8�u
R���yP��&��NmGwo��8�����.�J+�6b*g���7��x|Ɵ�����8|<]�wc�nM���)^�4�g�#tHD�Ny6(y[m�%�Zy��Nmu-\e�M�W��^ H�l�P�<�C'�z�ݕ�+L����;�jX�;�Y�~��aK��l�ǡ�ќ<�}��#6��8�D�=8�[Eu��x!�짇q�s4�btr��=���{p�NԂ��p������-'�������
n�"�k|Jb���R��������6���-�O�D�=��!��<������\Ě���]�ǁ�؜6�"���AqW)h���|7�`xĞ�#-(��~����)58q3���5��]�d������
k� �)&��e�<%*ޅDd���D�M���
��@�C�;�vY �u6���*V��U�}����uvb�F��y>5�o9wD�Y�:uX��y�K�2I���|�娨)�W��V�(~߶.���̯�Qz�|�� ��S�� o[쌪�fsK�H��P9)~J�J�^�K`E����>^��i���sOsN%}��m���g|��/���B|�j�:8>����#ϸ\�ʜ�vN㹞��;��^T�⸘�bp"x}ַ�+�	�IU@�_�0u�>lO"H �@���r޽��Y����I�!>�2`�
Rt���O��*��/�����i�0#LII��:�!'�1�v���&"�~k�T��h֎�+�e�TH�x�(���_#��V�&�d{���9�T���.�	�lY�K�'�n0��n����Bs~LxAvy_&�w}'�R^��^1Ś�+6�ޓ�����V1BA�a"���n
#���oT8m"R��jD����\�K�̈́r�&^C�+'b-3�]gd�+��,���WQ�پ1q,�x�,��˙�R\���͡.�j��?
�V�;�B�n}�}
��n�UHXtgy� To�lOT�X^�����z�u<\�i��ׄ���gZ�l� �~���R*KΥ��\X��"�v.����@�=�nN�!���%��h'*q��� u�*��WW
dĺmU��?l��[����ފ��D�۠�{�LtLk�)O�.�Q7iF�|(��h������]c,
Z�+:R��Ϝs��%�0+E~��H��A��ޖOD���R�f�T�OƟB�h�Wy�52^'�WW\�"H�6̿{��:]�"MU�0ፌea1�q`��Y[VZ�-?v�Ӥ�5��Zm`ᕖK�5ulVc���c���}X�Mh="�[fh�`�(ￍ(N.Fȏr�o��6���-*�	��tˏ���G9�BG1[�L"�{-q���V~�E>�E=f��3�7�v�;\�ҧ�E*\Ñ?+oF�"JV��/t�j3
�`�� �N<� U���/�D�1��Ï�}������"u$���*c�*N���~3����"���<��H"O�Y�W0W0��+��]ណ�/=
�N;�-���4Ý�k�� ~�9��;G:a�i�hz%ed��+�cx��gy�։�k����M!&oB�ȤטIo����OW���
��{��>�f[�����1�@x�g͡f
����R�%���n��/x�d�5��-����TM�z���U��昊C�_{W=�'�f`�ł��ܴ�˞j�U�7��l�)��Ự�c�D���z��&v�9��G��B�x`@7c�ޯ]�R���s���B���;b�
�t�᧖�|y�tt+��g���{s����'�N�f���L28u+r���_��.�b�_��!�8fH�Vy�8o��k�#��K|?��w-g�FP�i<������wR��6x����5�0~�Җ�%ߤH�@��|&�Y�-��N|�5 ?�w�	���K���8X:� 4�\"�`���8�LՋ�.��CG��E�Es����"g�O#nƝv�J�`U�>�s��
��-Ȋ-�S]Ϸs~_1�/kqFr[݄%�}��%�-�%C�x�O|l�C���y
��>��̭Ņ61; �ᛒg�O�hɔ�<�f��W��j��BB*�7����u��WI)����ۃej�hq�s�J�
�f��t?֨X",�)!�����b���3=g{�۴H�&���\��@	���0���V�(W�5У�(,�6r�m38��m@(Axt�!/����}h���ƽ��A|����&k�_v�5�κ��9֠�N�c�{z��VӲ6ͅJ�}������6��U5�4�^�AF�;�L�`^ּ���D�J�ґ<ܽ$Z��)k��*�d(���M�@'�UvEz�O�V7�f=�� �΅P=�&ʿ���*uq?��".'�1%T�4߬�Xz'O����#�����!� �~�2�1{����Fs�w9�w�1����X�l-�(��sƽ\��g��ɭ�@z���+����Q|޵�A�����#V h@�"��D���u7��U-t���A�;6��qH�}s�Ӫ�&Rcq��-�R�oaHp��h1�Ay��X��*#��h�i��c��H���v����xv�Jr�^L�Q�Lg;���B.Z���4��w���#�:Z���K�+��\�6�����qQBa��B�	2ԕ}ux�5�>�p��[C��S|м���^��{�#l~����5��[&� A�F�:�4�|g�����9�P���C��T9:�t�����;	$��r8{Z:ul�p��������q���W���O�Ph�p}��l�p��(;�<�@��W��li���s��7T�U�lb
����0�n�r�A�H#�+��Z2�DX�x��)`[_��~�*=و���������V?��ҏ4-��_��zi
������&� �[�'*�}në|�o����Mw=��g���` ��2�r(�w)�U_���h�1���-x����P��V��-o���xc����>�Ʈ���~���ߘQ�&ֻ�*_П���O�������H�����U'�G��u�´Q�y��;�Y0��w��P�d�?Tv�D?U�������:׆viʃ]A��e."s	K~��6ˎ���������fv��$�RD1+P OE�BK?+/���U�-j�o�p�ay�������m�5q����b��������~�5�o�����`H�y]����n5��#�P%ѯaSl�i��>K&D[�'��v�b�&���A=�}I��r$B3@.7������8X�'�Z��EeP�:=��8�I��>S3���0x� w�~��VO�0��Vc�����kz�U��Ælm���K��F���t�7'�fp� �� ){�E�H}	���j�kI	OA���2��L8\S�@O
8ǰ�uE���#�!<(�&˭7n����~���"qq?/�o� 4�I��'�I^��l�����f糭�A����A*����=/¼���]�qH�Jh���/l�=�x�n��;�����0������z&ǻם[|WIwG,�碉��Y��[P)�E�6/vr�(4W�ʊ��$��@?q���o�2io47BEX�c�}�&F�i���I"}�4������p����D��@��ة�PBp��h^SS��+<r�Ok�C�V到z7Iy�Y����+�ZGG�����-t$R��>�G:�z�(��,8>��g�ثbL�[I��"t�i�u؂C�^3�<Q�We?�W�ɿ��O��u.y��!��莂��r���"��^�>�(�CQ�]r"�P��L��-ښ�&-Ȃr�W�#G��}Z\��W�
�����!����"s&��틪�Oj�^�5u�y�u��W�K�Q��C#=�_�/�j��-/	N�p�����e҆�pS ���֔�sx����hϮm'������$�.j�©�� S�$2f��oȎ�]�ޅ��I�KL?�����b��mS���O�_![���ޡ��I�A�_9�lZV�W$ ���r ��$D�%�7��Cs����|z`o2s�,q�ˎ�ٗ��U�3}��E2�����ɺG;�L�rJJ��`Q|p���0ӓ&o
�o$��:��
�|<?\��4��i���_�]:k-�SN;�vw1���w;��5#2`�8L���[��&Y�����E�����t��<���}��Eߧ���5�>��լ☧�Ѓ`_G I��niKl0?���3)������+�uڸ�l:!�iCNv���ʿ�4��ς�g2��_�#Y���a�N�:�2�:�n��Q��y��/�5�b�A���A�ݝ��0���R�*l7:���y]��}�w.nC<�X�0�Y�f�ڼ:�Cևk��e��z��C����,�`��m��t!��=�I�Gd�q��$
:p)q�����M�ZWW�(veb[M,_�$c���j��
@	S�0�i�L�j���;���@9W������V������FIk���|����;�0�Y�����]���I�� ���d�9pa]v���t#"�RR��Ai=�k��E)\؍t���/���E�)�j��Z
�]��\�������P�zo�6ͳ��L�Y*��W��0i�sG�w��PpG�+�S�;G��et����XLѯ��J�y����A���l��1� 2$O_�^��{�	��W<y�c�P���.����r=�a}L���{0��>[X�m5����������B/R�8�'�?DL~��#����3wp��*,hUj�#���n�m�vӺ�Z׋9��&�d5n �0_6��zo��q�*��2a�����I�OM4�絵L �B)Μώ����F�<,jV52TG�%����U�v�J(Vo��Ԫ�b�!fP`�`(z�"�|������1^j��W�Vh��v(UQ�{ Q���"���E�^�]�~�K��d��͠��Ԑ0�3R�x�5agcd�:��&b��n�u9c���E��nE-1��+j��K7xl瞛�n"-��ST��H4��X��<�?������^"��"�C��9��U�"�,�!����x\�4ʺ%���%�
�`������X�<m0�jwf��� ��m�P�`��{����]#��V�n��Đ.f���[g��5���S����Zj%
��l�63ݳ�m���,�����	���͚�T�����L�MȆm��(u��C���8��,�6��\��d{~g��B�x_y���-�/V��n��Q0(�<=�N&o�0��1�t�����PۨJ���E��;��+����h�� ��u�S����yR�JK]�/�jW�n�W+����8�>,��&�+ʉ����y��qq�r� ��m�@8���]ŃC�3Q"�-�� 0'cuנ��˺�����dZ�Q&Y��6��Ңd���\�;#�M]C��?��=C�ѬÁH�i	5��X}�$�X|j4���rHiF���
v)ϢQ�kt#ZS�����������d���=����v�:#��L�9���?PY������A�n�GjŮ�%���j����d1���^{�+Q:�\��r9/K�ȼ�>�t�A�TyE��e�(f���n�Y𓊎���Պ�{�G��lH�"`H�%,s��Ӈ�}dDj4������5{y�iQ�ԏBA%i�}y���~��/4h��x�8���7���"��������#;�?7C��l�"��~��4Ȁ}����Zahf�j �%K[ !�8E�̪��:C����4�(�<�J�d
-�i�Q�N��Bvl]H��n��?@�����^\�,<�~�6��4s�@�H��oX�N�K��U�^����a�3L�$�H2��-��}_4o3����,A^-�/Ew$��X�R-���@D�h�V��K{G��r��LWΒ�OeӗL��2	�8�m�FMT����3>���h���)�Vc�:b���4
<�Y~�$�t�Iwvx�`�P�#�ŢS��R��qʳ�����^�$Z_����!>e+>�f����b]�>�q�X���N.���;��������ǹ,����C[�Ү4ѿ�l��������*�5��YHѶ�Ƅ�}��N��5qb3P��H*��G�3�XFVO�fL-����i|����7T[}��ڲ�!���,T@>� t�Q=N,Y
w���^�A���ޑ������9 Nt̲)[�1�R��Zg�����	gQ[j <��=�3\e������E^�b!V�b#�M-8}�I.�����724�DvN�0ZP��x�,	2��ܥ�`��1���ْ���QՕ��6�*�_\ڱ|�%w�-�#Ba�+�_,0lfǜ��|�䨇ɥ��,��-3H�v� �|zT�0��6��e��;(6���Ĝ��PzR-._�p�~	�D;�Dc����������<���ڬ�"�az�6_Qe����E!O��;��U>V�I`�d~��V��ӿ��>��6#K&	l���m{V�PC�d4���si�Rh_p� ��k��ثJ���R�'Z�l�Dq��^����	nmO�(�d8���W����-�M@��oYl��!�Y!5��fx�y�	���F��2~z�s�H�{���e���w� $�s�gK]���!�g��	��궺j���ߊ�?�8;�jOu��
�8���	Z�\�\C�Gb����9ye�]�����㠴R�����½-�'̾�uD�V���j:4<3��k'*�o�O=���N��Oˈ-�Ұ ��K�Z]��:����W�Nt�C=mȜ�1[�C�턽�K���眬�������W�)��"�R`~1�WCxn��\���3t'p�!�]{9ޭ��ƌ�8��}�Z��3�~bH�qf$��� J�}�3v�g6G�>��U�U���P�#=�%S`��\��x�7��������5��~��׋T�K���:���Ԕc���܆�����̖�xd��Y9S�ؤy%\+�ٚX*i��m:w�GUɰ��+m
ݥie��;d�������DN�#��/f� ����� �>R��>QQ3|�+��l�����r��IRK��^*�i��DO'�����z҉}�5�j�QǠ�c[���x}1%e���Â;R��hJJ����fz��O�-ẽ�b(��(���jI��(R�~Cƛ�'T�	eʕ�����;Y��Z��W�ٓ8B%��į�`�X��r޶"g�P��m�n�^B�J�;�G�X*��ڟ�0��J_��}�F�?�)��ē��u�GJڊ>�1D���|��nڨ4V}a���j��ꊝ��7����9����Z�8ҍhF�I�|U1��*ю�mFxo'� b�|��*��<�l������F@�v5�_�}}g����a�o���U��(�f��X�s��,D����(�J4�(:2�4[��k0 �t�5)���'R􇠑�[BlZ�sZ�JW�r!��ob'v��(�%�^3��EfH	��(O��ԶB׬á��_6���$��	 ϴʰ����U�K'�����Z��0�b96�W��WiF��h7�		��G�pXhuAu��n0T�B�4�tp�^�^���(��9��������S�:�<�_�'�ǳd�:�o�.Nhk�p�s!����lJw�������ޖV��eL6��s�[��E���g���pӿ�E��
�U���d���=��[]��b��\�[�8����nf�3���^�s.��;�IYnÞ�RG�D��?����| �h#ݟ����w��
w�-����r�4v#]��/E6�{�� B��Ϙ�S�բ���!N�t$��5���x4?P�"O$�g�*�~kʔT>�.�<�K!X��1�Y3��[՛�Ī�O��7���ՍK{hbx��b�L�^��O��B)~r|286��'���L��;�4f�b�z3nx�W�Ѥ��K�=/��%�G�hA�%�&9q�H}�r*RM���*�
�;3#�MCD���aU_�k2T3^�&�N�#���1�(��=�Z�p�O��m�U�ZcD�����15�Q����8����B�Le��\?�E)�y3 &���׈ɸu!�>p�[�<J��n:�#�A�����Gi��u��4�{$��%P!(��'j��2��J�%��Xd�%�+�_�\`Ys��_xu����DO�6x��^��؂����b �$��w�>*�CcʋDeC.�̓���o%��L���v�Z���!N�� �Z�ū�Ӳ�"�w���jr$x�(0G
�]������L����;x������yC�����S_�L=>�0[��r�k$X��"�O7a3��_#kCh>7���4z��/O:�g�<A�	�ݻ��u�H`_��\�*�J� �ui�#K����	��o���G���*��\9��n)�"��Tt'�pb����عY��)o��	�rO*�pgUc���`�ʴ�;�+�u�;X�����%��풠�b
�_���&�P}��Fh�t�c��p�(*�X'��Zz!��.I,�S�H�x��6!��[��Ev�Oo)�n��������\�Z�4-j�ƻ?��W~�����!��}�\��l.��k�ˢ{'�BAՍ�������i�9-���ǌGz����s��?�%n��+\Q���fx���o����va5͔����M:������Y7r9q0(X�mŨ�L����]���-����� ���$�d�5��
��f����6��zS� ���R.�nz�v�̻:5[�A��\�4�r��y �O�����=(k�BĊ�P�_w��g�FL����_�:w����;d�G��ˡ|���~�6�����
���^��m�!��v�-�p�x��#��dd�"��m_�����)'�+�	/�����i./�d��(Kώ`�"�g�(�&_iF�卭G]�p�׫&G4�t`|Amtk�O�@Hxt�}�!�<kLC_mc>�[쒰���P�*�ȕ��M)�w��=X&/��W�����eô"?4��������;c�2zhse�i�����RZh���?⌇\�J�&� ��������B��,{�����G���ޒ�����{��yj�|(Eu�s?��p�a�z��������P[�D?�\tJ�œd@<�	EF�~#�G�),��ܞ�c<;.J�n� C^-�Wϧ��*:��1��������7_M\[�7��J�q����A��ݼ�D����MP2'��#DfcD=�r��|��@��ɔ�ӟ���������Bu4�s�$9CfQ��.8��of�O���lF��^n&�f1��X�N��J"�ߟ��;�/d�d��{�W���/0�t�#�&�\Xh�0v��8*e�:!���c�e6�v�d��Sy{~�
)�L�'�sZM�}��&ոs\4��%�4��X4���,)�.ga|�nNT�Օ[3�*:�����π�� 
����ݘNiu5lU��:v~:gC��(o��<��+��eg������Vo2��z�����d��ie����r���w��(��q!��\5����O@y7XB�E#4�K��ee'۩�Bs���"	EG��\�$�]�kx�|��g�^H^��^�R'�p�����.�{6g��-\>[��
).<SD��_YK�[�L��|���J�g`�����I���c��P�M41QE����;yF�Up�8ĝ__Ǆ]� �f3���H>��c�?�9��1V��|6��i�k�G�C[���b[�XM�%i�+B:I��Ra~�d��4iV�\xf$�Si���)B�����r!Iq�z��9���-"����#��� �i�ߪ�߆���/CJ���q9�.��f�&�8A)!�
Ў�#�̍ WK���7}����9�g�5��]���W�>����'�=#dS���`��S�O���	_$j��'������j���%Nx�)�'�7,�� ���J�Y)T�Č�ʹ�(1�����O��w��陡?���7� �J/��H�,�	i���r{�� �[����Y_
sˬq�)t��c�A6S\� �YQ�����M8�P��_�5�����.�X?�1`��b��@t�	繩( �'� �����6��0��j�+�h*V�.i�Q�V{Y1�)	��恩Lyu:fWE��x3��R<�-R*4z�d�N��(�1���HA�t@?q9��Ԁ1�F`��t~�d�}�f��=l�s��$̈́$h�GC��g��q�\�mn����`[ҫ�H֔�|hÉ�+���gO_�Ɣ�e��2^Iq�
GG}��>ʹ��V˲`��E�N�B7�1nև��8m�s9�2G�l@�^��G��
>K���r��m����0�Շp�l������t���j�=aW@�#I�f���Q`�������|%�Pg��0���G��K3O%�Y�3�:WQ9=��ʊ�|�fQ�M `,!��D���R��5sGD�^�.Md�~	�l��6lx��MK�,)�Ď�1ޠE�'%���ܩ�ݱʉ��(���7�� S���Y� m6P<�oT�z2hp�����l!�E�����\Kk}�W�Ψ��l��q !�`" X���|˳�uG:j��r��0M?�%~D�Y��������U;wT;+���Y#�'�.g�l)��X�Ȁ�χC3/
!��La������khuk�-�����YC����6�@B�v�v"..I���/�A��$�U�2Õ��z�Fi�դ'�`=��Őڔ�`zqT-a���x�q��k,,�d���ٿ���L�>/��D�;oO�'χ��A�[9��J)j�5	��m{/
;}மp.4��n�;�^�]��'	��TH�C�����M�ja��t���D0&c_��ɵ��C�(��)}�G2�4gE]�|G0ܨ��yܭ�lK5�_��X���G�N�`�X�]�Ȑn��00-ɰP��"�:���JÖp(���G�?+�2���t<��>LޘXշťW%_����bO�n����U�������Z!�x���Zf��a�6�W#�~�,%�UN�`>���,X�t����}����%<=���f�, 8��t¼�4$���hF�U���cGd��l��;�Ű5PA���Ap�a�Ԥ.~I��ZyT�ҧ�Ə��c֮.������t�a j&�N���j==
��5d�[�RL��d��A�N�ʫ�iɥ�fe��0���++��=��A�?Bm��#�xx{	�NR8A��$���a:fYȱ2r�#6��v�c���ȯ����(F`��/vh�
�?uS�t�%E݈G�Y?���J7Ql$x���c�+\�XnL
WG-5G�:W���Q�r��o��-^d���h�6��+�MAC�?O$�|���;��FLUF<Q���o]PKL-��7�����2x�Կސ���s"��x��pMy���+	I��ge�=��j��F᠕F�$z�9T�7E��B�SŖ]��^�\�L~^K��}����>-���3F_+�'D�D��T*�0`뷗YS�"Ј4���=yp�$d���hl�wJ	Rjჺ<M��g,u*�Ď}e���z[�(A��yU�]O�C	7H�g�~pVI���=��d}��4{�MB�Y���g)R�	��j�w1�� !�I�~_��\=(�Bԉ�D��Qw>��`-
6K�T�U�1���j�LգJ�u�]0~ ]�D��H�f�N@N��/�r
���n��$����י)28nH~���>�2U���ט������K���Ã�5�Zx߃� O�eD�����Z]U�^��ۅ�m����p�p&��z���j�>��k<W��!Kƫ)�oZ�TC&��+�E1��b��:�Xb��S'�k+J4��,b�0�f>��.$<H��q�&�\����xp{{�=WT�|X�l~>�������a�`$-�:���!9���>�?A��Є�S�MY��|�-���5�Zi��\�����=,ͯռG���(m�����5g�t1�-o��;1�D4Z��)VC�� t�f���d������rc�t����Z�z�[�]�.��;�����t%�4A�&A O���?���V���$k�����V��C�V�����Y�5)ė=�c/�׋-�g�i�R��r��\@wC�w���� �N����n��Ĺ�'�)�>���Af���$ ��\�%��H!�Ҩc�nEy��?X��ۈ,׶]��R���	.ÛNx�d<O��hQ�_*����C��Z�����>�ʹD��"=:�'җ�����=E�����0�ˏo|���B�0l#:x!�?�ڭ[ޣyμ,�%��C�Y���*�0���eF�MMh������*��5���0oS�[�W��������3�q����,!�k��/9�?�����#[��r-���s�_����=�jKW��c,�����	ƋQ{r�	\�Y�����^�K^�G+��L7J�͝E�F�q3�qq�f�r�e�!�d�F�ȇAqj��<��M��R��.S
G|��l���C��7��j�jX����d��w�)[�íD^ׁZO��!�-4S/v��K�Y�n���SP5���{��A`!\���傓���T��r�M�á�p�󆹢fHܠܥ�STF[�֙��I���,W�C��;8Vc����KӖ�-���	ϻ���V	��4�� %��:�!���M���-���Jv��xA�gw�]��ohns�<647��kM�P�Ǣ/���gr6��۸$�g�r����f>�Zg҅�Ɋ��Ö���z�r�$rb�@@G*��i_���5��N. �ʐ��L�6=4�QI�7��_^��,�y�7�����\�[݄���!�G����Zp^U���P^VO�Z�"t�����|�³.�֏"�?>Ph�9~d���/�B��]h�a�Sa���u��g�� ���T�	���L��?�MHLE
\����?*�jV��A��s�y���6I0�6�O�Z�7$��h�O��Ji��%�w]���d�1:0**xusZ�/uK5t��z������6����mo�3@~��ȣ�����HL�%���w�~�+����/Џ�Y:]E��������C�=�!�`�AJ��,��?}E�P��h�����K7]aۿpPT�j���W:W�a8}��I����ڸ3�\ l�<(r�LR
�=���VQ�v§���7����G¥������E]N�ֶP&�J�l�¶���
�5v������@a����p�����f[�gUC��j�T���v'I�֠6���a#�	~Deŏ���q%��.d[σ��E�}j��t�#�������T��E�#�6R��$���ߝ�bZ2U��j��%��C�j@����6��_
<ᴖ�lZ��X�� z�\���z\���md�[~yވ�w�~�������&˓�z�SG}G���N�d��p?^3���GHQ}T���mVO�<�5��RHl�����g�3��S6�N4S�S��q�EW�ZQ�>l�O,�Ǩ�<71+#n�ʊ�=n�A�捂ް�XKy��˟�Q��Nr:{��Z �7Z��{��ϯT�8�;L,��7o~�UVc|"3V�L�q�(M��شR���&%|33�Ac@\$��2�Š�M��7M)�/ �Lhm`��鎦�1��sT��Cź(g��m���q�:*T�a�,�[�d��"x�#r��B��{ԥy���������X���Gu�#.�R�+���L�z�XZ*MQ�u����G +gp��(n��I�+ahf�ؾ����.�!cqZ[�
�W���c�#�t/��]SFU�Q�i��)���u�������D�&K�����t���g����kd���.~9;�X��~�4� ���q�K�����=j^CGƳz�#r�����N�'rKM�#u� �]E;8�Ǔ[H}c��H��0-gs��Zz_�X5���*{� G4���V��N%b¬\:oG��Ǵ!
&:[ٱ��!"h�ҳ�h\$.];���4�B)�!�$��C�+���i���T��{:���/Ҙ�u�������K^+C�
LwKR���	��p;m���Y���}ȥ%���1n&vG��e���a�0�|�y����D?�*ቮ�O`5l(�UB�a��Vq�w�F"XEǦ'�O����4�i�{:������9�����E$N	�����2K�N�C��`�;)ۿ7g�W6/�:����l����3Qp�\��k�)��팩��8C'�M��S^�8�ݲϦ��T}'x�c2��������'��[=V���m ?k24���A/'E� ?6E��Pa���jM�yT��V�rj�a|ޟ��햏;�TM
��s�8t@c.���u���2J�j�%-��%NM�7ou� Jr5�����0�=�Ǥ�=�� �>u׷0!�
��Qsԭ�H��,��Ue�K�� /�\��[B����ҋ�$lكI��fS�����>��z@�K���SD�����$�>�ؒ,!3��c�A/Ԝt;�7�qK��jI�0�rB03�;�~�Tbđv�*'5��{�f|J���n����>N�$5y��VOW��gRF_��?��_�̬֞��X���ԁ��XK�:�9gu&A�os��� ;�5�����HQ��ڇ"�Z&�+-Jy��1� Ϫ��'���_���(��q������В6����:� [���9�T��t��3g�N���sd��7y�S��I/��i-�=������n���뀈2��/���'��sD��x���_L!�.�������t6��nj����,�>�I��9*M�r�BI$��H��:�f���eX���@O��P��7X,�pEmh�nj�ArH�X�V=ȉ�x�1��vh����Θ+��N�W�����BO>6YS�7��[�۩��}��@�|��ك�|3pIC7����ϿD5�,�Sc������2�P�eLژ����K�E~�����M񜒯F����q�@� ���Y^��.�����p�.�`_���f}�p����ʍ��pOJ�u+��~䒿��@p��r�Vv�ڨ� %c�Fs$����h��XI�.�hT�s�SJ�ǻ@N��5	g�UO�>%$Fi37CrMtb�u�sM�����,����)�43@�r�����S�Z����*k�_�.�9NF-��R����ņWD���;��#Й�b�l��p�[�B� �K�h/��nvt�Ɵ;(��[[�UDj�oNR�&BE���䪋^�c蒥����	E����'h�/?Ju ��:�Հ�r߲�/�( h�B,��K�\����E��_�"�����`��zgQy�>����9ONh5���ž��e(��;j�4ظ�v2V��.�v�	�pn��y���z�kc_V�+���' Ф/l|u�H]�������h��J��,FJ`N�N�	�� ̋�o������@Y�-)!��:h�6h��A�g�4�HՈ���5[`	�Z��9���-ǒ�k�3r�{�MG�8�:��<�}�0XE$!Iml��3 ��}T����8kB����(��{�f�"��dĈ��mrLU�9�\�:��������!Q�푟{�80���4|����hF7҅u\v/s�~����q �^���S3��;L���c�.����)t�#gr%�f	���b�ZX�߬��H-�%���^D��ڂ� ߓ��MWnyl���"U�CL-��S����w�n{�ϟ-��"���U�b[6s=�-'Pr��Y��D �Q�bwO����|�|�ג��<`rʿիR�-^)�>R�l��
�x �gϪe�ŧ� ������}��.�@{��������@~��g~q��v��C�F
�VA�F+=9IM�u�zB�;>��MZR�Wt^�D���WT�DA�y��0
���]p9t;�Aޖ
����z��k��}�N3�tF�Dp��VZͧ�Ջ�e0�k7�{��
�����жN��/�yI1�G�a��x�܋�+���lO�2I�U���K\���%Bz�4�hz(m�6j�Ӂ���L��M�_R@��P��@/V���3�-�5����_�tY!05�G��%	�?�#�̉E�pe�(.
%�M�d�~8�)�Sw't��砶3{���f]��ڸ��d7�&�|�"�E��W�-QfB���ε�F���dJ�|���)��>�1`����P?��q0����Ek�V&�[�r[^���S�;�Z�MAo3�H'��L����D����;�`�;ݏs:t�}]���p�����&��s˃���4�ɷ�Ѿ<:ړ�@�8���[P����=�� �i��ɝ.cK�C����Q��/�AN�T�]����B�p���p3�zxV"^y/p�5')�B�0��x[�R�d%n��2�yנ�C�쭀�B�S��}�wX?�5�Ϩ2J�Y���*��3lhSx(�|P6�w����1���;�
�?@1i���Nr�7���������+j��2Q\�����*���(ͧ�R��q�Z�֭���d�ÏM���ν,	~��u��?H))�r̖����=����%��26�u�&1ϟ*�r��fN��J�Zs�G�*~x|ho��Sh���mVE��+W��Q�u���J��7�ҋ.�<,Q��Fx�iU��vg�~�������*�n��I���vJg���ɝ��
�yǻ<ŀ/q6�>��*�r�.��X�%������gjJQ� ?ԠF���/����[��ah�To4��1a�j��
�(��$?Wu�9Z��c�����热�����!�$��q�9��C���KC��Ū�f2= 	��q�;����d76���p��z��s��%ʵT,7$������s�
�x@�)ٳ�]��� ��D�o��04�a�\k��;��g���R�d�_ �^r�'�^5�<l9�{���q����-U�ϖ�D$��(��8T�%����s�%Z4_���uqLz�������F��t��`�1#t6Zm�����.��a�.�/dc�|�i)�@E�g�@�ʺ�Ȁڟ�ӊl��辨��t�Q��*=p���.����s:̔@3�\ �Xp&'D`	�)���N�eޓ��ӿ�m��/:z�Wϳ\�.4+/q'Q��^�S�S���j�!
��WY��f�~��z��d4�W�F�z�H�4��l��J�zq�� �D�R��M\*
��9*b�:��et��lP���E7GY�{T(w��7�6M�IW�5ǥ��l98X:D��PW"����ངR{�V����n�n��S�����w�1���W�����7��O��Z�d��\�8KV����f��U-�]%š�'|\x�c�-�쎯�7R�?P{�Q�l��~I�($	td�+�?��}�^��c������İ�f�U�j�,>�t4����)���=hO�����y����ƜF~R�{��0	�}���7E���)��J
	���i�F *���,j�����HTN}ɘ�36i�{���=�ǘI7}���(�S�r8.d�qK��\z��j��ڙ.�$��)G N��gq�����7���8�(�a(ˮ�JzC��c�\�B�4W�b:����O*Ύ�
�������!�٥oP�boP��_���ȄC�Z&���M��D�{����#���
a�7e�G�����]��ߧ���If�����0�E���?s�75S$ԑ��"Zh�X0���)<��G���<������|�g���
����#���,Ƴn�y^�"���||�n���p�hZ��m����\TI���	�P�ɱ��g1��������\�m�PY�?�����S�ۙj��jj�Q5��S0i��\�%>>�Xes��Sڥ�p���ͭ�������ǩCeR��\�);���=���p3ǔ��wF��:��)�2V`�Y��.�<`8V���W�L4<)z�g����4���gRCa����Yu7���!�đ	�FnkhM���t��wU�T�)�{��BE�����o������
H$2��M��i��m0��^{Zk�-b�5o<�!3cO�ŉ��&��H�Ɋ7�����%:�ͮ^
�(��ky:X��(�ҳ;���j�iK��j�\���X���:g���fԭ�"�����_R����^ҩ�(N� Λ67����p����0��H^\r������$d�?�	�u�oQ�̜� ��E��'�i��j}`Y��@�A���as��+�.ϒ�Ζr}���K��`G��ϭd���cJ��{�.��o*�5�b!|38�������e���s�\�\7����!�{�ʢ�p��7����梺�����f==_Wu�!��-qͮx�z�7nd�6�Lq��1��#^Sޭ�,A��jV��J�/�޼���&��s��x�7�>rY럎kw��)V��ř14O�$o UBt�J��u�>��֙O �3��So�NL�`e\m�7!�֕�	,(�>N �����gX�^�*�����Ĕ�j�Px�2+C#7.�9��)�a�>�'�xV\5ݍ�'_�%��al����-|h]��5��Ag���/=��-�Q*���理cB@:B��0�`�����;|�z���n 4�q6<BxS
�'���v@<��_�!�Kn�������PӶ4�!�fW��,J�&Z�^�&��n������,\����$+<:e�Ζy�n��P��.ଟ7	����8�g)?������3NCՕ�[<���V:�`��GI�n��[���ry{ݐ �yX[Z��t��7yDҼE]ETU9|ժSu��]	�Y~i�a5��~�^�4�4
�D?�m4�☈y9s��c��l�� a�7�����_�%�ԙ�rM�ɠ����$�Y�sh��_������$�����[JY����{(gY|�R7� <ݒ�&���M���J��d�SLzc?��HB(��!��v�bG�U���|
�z~ ��9�fe8Y�Ѿ��m?����x�́�{m@;u8 /)G���C�`Hh90R�F,�E�O7X�2�ݯTX��n�.��,��(RF��ǵ��������X�I�Đ������.�&e)-��R��Ƨ�#�I�k�e�~=��z���Et)��IϾSW2T<�]5Z�?���G�0�m�����565�>0v�@�9Rk��C5_@�7��MEpB��O1x��h͹�"�Wc�����q{��u���P ��۩m���:�{f�QwXD�ǦXv6��$���zΫ�4(D6hv�9٨D8���9�=yb���	�Uk�a�D;,��$�ǝ��z;5'�ޘ�Q]Af���f[WS��� ���.w4�ˤ�3FTǀ֊���U˜�ħP�J�Ґ�u��ٟ!�F$��*&���:���X�L��{,�����͒*3E�}Bģ3����������!��y`ED��d�pf�3��
`Ƞo@����mp_�籂�}���o<]�uU�G�b�ΐ�A��1�V$���Z!���X�pg_��s�ym�WJos�Iט��x��	�IVL�0gz��FM��b��a��B)x��q��̢����=�?S2�F�i lؼ�S�[��|�P�ֱz���zQ��㔰*��?i�E#�ŠT;��k!a�^L�,�\p���8��p�Y>l{��ɐ0`|�x���Rr�+:{ױ\5�0�u,ԥq�X�M��1�#�Oy��O��SS�b�`%�)-I�����K3��p��S�.[-�u_��g@���/G�e�e�SOԧ�Ď��8�26��S����z��J3����	S��~ۉ�������3��A�6�Lӱ\�H5���,����w���2���3>O]��Zo6�=}�߶�k,�Q�!�v��=�����\x^�I�pRi8����}9T6��?�:�4R�Ҽŕ���
��SVGM��A�Oq'�!�L���>9J��!V�ΪĢ~~��v@�>���T�C��)�w�M�� ��#
b�VUı�w1��3q�{V�mf�2�v����0=<�ڢ9"4,�'࿊\~����c�M��1"_��߄�24�ge��^��J��R��lk����k�%��g��c�gKT����X�ogv'4u/Ȝ��h��H6�����`i� �ϑ�;�\��8���!"U��1��|1$ϩ�gU�9��q�w���R̽0��j��Pc�O7E�J�u�Y��8�N�z�l���*����! �Mlj/Y+u8�:_O��.Ω�g^v'�~�{W>Jq�(��b�cc�hi�ǧ�?��wZ�:��2u����qf��gUź
eg5J�<;V"v� h�J�&"j�fP������!��q���^j��ԭ#���~t�Z�������Q�,�F����+����Ⱥx�4;u�<}X{��EK5��]��b�
�wV�x���m�pX�V+�C�M���'z���0?���O��Mw��#1��Ш׫`��a@��rC:	�}�*V�K _��@���� Y����,���*�mUȰ�� ��$��	�<+� Y�O�5+
k����>?}1F�F|ɉ�dB3��\3r��W���J�wB�v0��2'�{���jW�Fj�(�!�%`/i.�'&X�{�j7`��B�GJ��x֬Gd췢=: <3"d1j=�^YOӨ�>���\S�LT�Eo��:�ʖ���r=����P�q���阬�K�G�YH��ؗ���VE��eL��t;i0�0R�Z���du���}]Uo��Qz��f�+�loĲ�\��8��׏�D*�>�����)�Ѳ�!�z܅Hv����W�QF�x��<���h��	��Q�D��t6}nу�p�� �4=�2���@����%�[4>-9���V������=��-�� &0
N���S��I;�D�;��lS9��U2g'�Y���⚃М�'ۅ�w�qO��D�a�k����Z�=�O���k�s��#�{�U�K/���9����Ft���߇�����n��L���}V�Q���F��΢]���'50��*/����TXu�<*c�F�޽������k-[Mڝ!���]���f2���ڦ!��*M�Xfr����ld��A�'��Hc3)B�y��DÇT����0�B�� =�Jcj����@oN�e����0C^V	r�D��$3	�>0Z���Dto��k�)μ$���8�Q)����G�@4.?LsI�u���|��O)z̰Q���8Y��zK�����̘�ܦ�=�,�F##�n���W�zp����e/M�f
��-����s���`ܖ[���sБ�Q��0�{,nEń�)��o�r�`��f�49��͵�CgZHH �q�?R��*�$_���옴�폽��v~�Ւ#:�=�%�|l�C��ׯ���z"h�u��g�R2�J��;#>�
�6�&_�F�>����ZBC6Ro���G|YҦ�Rd�a�$z-T�}`���vz40G�^�z�K��j���E�9�C�� Mj�. (Y�o�4��f�/��n�w=�h��Vl9:���T���u��
�&Q�����1HeVڻ�do�t+l�3�CC�A�.b�3v&J���L�l�B��QU��n���
0`v�}��"5��ji|�"�I�����9�/5ьS�!Tbӑ(A��)Ӥ����������/�o�Ϭ�%ft�D�ER:Ou&� ���6%�.���vx/|{Dw����9	�p��s��Trd^���a�a�T~�&{�ܽ�l)g��/L�'I�AjE8�������!f��gu���?f����[�}T�����2vh:p��VO�]8��Q ��k�l\�^HP�t�)=H�� �,��bR~rq�\\K���5_�ۿ�8��RᙾY�� �a>��e'�@��v�o����3/���������������/�"�]4~�˴S���|d�NB�rC
��
3��	��,�
��c�Rw�M���@;��o�*�i��٧bE�o�W'�=T��
g�O��5Y	"4���&(��x2��nR��Ѯ:!�Q���dU�մ&�I:u;��zQ�f�$���<e�f���i��B��@�f����x<(�/}M��"�o���:x�������̯�V_��b��;��Ug�q���^�]��A5(~����pD`j����`��u����m�7�+�_(E8�"�����R۩"�����<��˂lP>�)obk�����|iIR(5�/�'/ o����95���wd'A�Y��Ɇ�g*��3��q�bqB�f%�Ӧ�%tx"c�?���nl���-έ�Y�������g(n�߼ۯ�J�#&l�Ƴ�?��@S�h��ؔ�i^�3����3��4<6�({4f�O��p��W�0iB���z���E���1���w����%� .���?���Ykdt���4�<p�q�;M��}���2K_\t�ʯ?Z\�r���Zk�Nhzw�*K"�J�t�>Bq���{$��D�����>�3
�v���M!.`��TO�j9'�L��ІTM�Md�l���I<�Np�>��D�V�2�'��n�V�)�8��$�Ŭ%�N4Y4�����'-��m����b��^���ӿ��`��|;��΀н�Nd�����6�� (o�� OW�}|]1�y���&��N�cu�q�,�4��Tpn�K�w�s�>�7��U�T�  Q��Q��2( �[�y�-M��XE(�\��ƫ��Ћz~G�]�T|�w6��>�D�Bh�>7Xw�l��E�hh3���N1���>(�ĜϥK���I$�K������6Q8T���)���rײ��eM;}����H*P_Y6y����5���O�w�� �-?���m��d��|1Ŀ=-⒈�ƃ���T�Xy��'FR��Jl>ږQHlW���Ɣ}�o?��g]E�V?}��d# �*e�A7:�_�z�����r�D���?NGC���ٮiٝ���cK�Ep9x�ܦ��:|�3���҈4M��r���Q��|�"��Z��b6%b�-����{��S��cr�8��J�4�$��j���R��&�w
�X횸�f���~�YK������c�aMq�
�&j���l����9腏�Sg�	H[5�j�&V���^���8�߯���Qѹx�}d��W�D����(�Kǘ���N^Z>����~=�91w{�DnX�S����X��8��'�va ��8Q7���ŋ�+������5��<rw�<yq��F��7e�Du���EU�~�UF�;��ª^��� ��юI���I�9��v$<&ln���N���%bzT�]Hx���qI��s�3e�[�����RJ�X��ڌ���S#�24�X�ĊG�W��Q���qF��A�Q��\�iur��<��g���v��e�4G�$�oE�R�8�P,���2����-8B(��l�P 9�����0�a����*� ���:��.f��}Q�V�Q��v����0�����zD�:�ǯO�
-���{U_?�$�B���/�<�c� alb�AL�ę�,���B>Ϟ5��u��jA��X�G+�������>��-�63���d����(a4�n����:�7x�G�A�	]���H���jp�/o��&���8#���7��Uw���b;؈T�#��c%3�8�r�9w�����{��Ϙ�KYB�_+��%E��m��+\�zI�V;�	�Ѱ��	#�u�L0���U8-���ێw��Mf4]+0!�������5D=��]o\,
��2��c'��(˒�g�i.晍��7������s���vE/2ӎulu���Ю��a�V��ո[8dׅhN���n7FtpwH�8�0��B�@D�@��]5������>�AGW��ə�3�[7�J�\�y��N�_��P�nPIg��@O�L:0P��?U=SH�C�&�]��GĖS2��֋��l���a��u��F��f�
FQ-.�7ڮd��}"�c;�3��A���/��k�:��䟥�84F4V�n�1��\AH��p^t�<�$����&��Wv�p�dՎv�K!c��tʅ/�!����C���I�������G��q��'O�8�2>��Od�3���W@*;ƅ���:��Q!����<ㅭ�59�Ie�NԜ���hpF�FV�����%� -��RS h�ϫ�U ��K�})�
�VͿi���>ʪ���Wѧ˺�h��?�@1�Hr�٣5������=3�M�E�@��ܓ����[��
�/pL�?�/�	���s?P����D���V�dc��L�NY�i�&�mbtL�D$dAri請��j4n䧃5&��P�WWq`ߓ�傃���@��ٌ�UlGE��z1H�5�As�4�{��t�W=ۜ� L��&��wq�5���bv�h���O%�$PL&W�W�r���~��u��Ō{��jL'���*��Q̃;������K
�D�S�H{���"�+V9��؟R`�
+�b �uՑ���~�7e�~���%�2� đ?hʶ
�65��2Oŷg�<�@;SMY��2~��\s.'�y�X�^�_&HkT�����y�tII��/{�)�U�?���{�N����i�v���K���O�/�6�+���|��������5]�y�<�MF%�!Q_d?g�l%�*P2��I4w�ͦ�|0��a��"�S(�QD����>m�k�!6��u���<�(��G6Q��� |�u8.N�Xbl��K�%NdH�1�����r\����=,��cG�S�}�=D�&H���~��vD~t��6E���p�|!wV~���!f<��Dn��iz�Aƌ��m��|�fR��?�Pdorh*\�����;+)�$�|2G��@�� ����22G�1�X�y�T�m bc�u��.g�[_�1����tU�Kv��u?�ZB�!�Z�TOe�����
�y?�uUo\J�-�\�����t����`������ie"�����ia��[P���u=�F��H�(%�����1-���+,�/�r2��ͼ��֋Yu��y�m[#��
�����R��Ȍ�1��4U%�� �V����e�MK��ʩ�ɽ��Qݍ��
�<Jf�xQ�� R=���	��ԇt�e�7��mTυ���4nD�s���{���ƙ��6+�e�j��!i����w�|6��p��ȿ,]�M[�U��0��K�!�����(�� k���BL��!���y���1I����*-�S���"uG,����pnYI��Fj�T.���O��r��"C]84�Ӡ�P	{^٫C���Aq�*�<����՛�c��!� �M>��o}��P4�R���H���	���K�x�c�B,_�1��Y���j8����(��o)~�P�en��E�����+Yov������/B�n[�Ql�_��Gh����v)�)���z�N=!�?�h|f�WPh��T��	q/�gߔ!��D�a^�<�Duz����C�iZ�oΑ�\z���Ě@zs+�py�@)O���Kc�㈌�������d�}���6�V���i+w21+*��s|�':%Eh5Ï�X�{�$6��2��5��#�VP�%<�z��]���t(-�� ��/Cib�O�ҧ���9�G�y�Ŧ �����G��0�ΫM�ɤ�Ú�`�ǽ��Z³2R����x��� -�xC^s9D�5�P���I��;p 2�e�7�+9�hzG�gz�%��bh�n*Җ[m�C����z{���m��e�Dg�QQއE�/���f΍������o�o�_k�b�e��K�0������-�S
��[?O=?j2[�S760�����Ɯ$|ѥ�wW�S�`ꜟ�INgc�	R�aE#i��%�Z�j��8�������$6\�����H���9i�~�և�si��Υ?�Z�`���c��K�nױi�����+����������-��;�l˭ҩ��0�o�G��-O��Hj]\��3�@���9���Y�K����2ٛ��=]�+�R��ŷ�4��r�6t -��b�-�a�58H���l��p=j"�/3�� ϡ��s�@���0�)'V�źvS�Ϋ�<��&�O�|KY��c����B ��nD�В���ێq��Yc�d��*C�V7@MI<]¬��\�f�y"�b�q�n���$����w~��8%ah(#���Joqm8{>9T*���|R�`NV��v�w�%nAq�x|í�ߦ�Q`�B�����Е����� �{P{�ˆ�u�]k��x��"x��r�Wc�oD09?�Y��`���X`� �ٯ'�U!.7�ρ�+��M�TFu+�������� ���+8hŧǜc,CM��]v�����.sX����S�K
Bsg\|g���q��l��Iơ�.π>�S�"��~�+�aV�H��2���J���q
	����;��˨m���ԟ�Hm���hT�u��b�+���0��'�m�κ d}3��Z����M_K�e�Ŀ�,���QDYX;��lk���̙*\�M�Q�����V�ö`]p+�Q�[�U�QP	�^.��;1�R�Z�ʄqd��O_�x�a����47%ź��x��A�u���`�̼���8��	��{|��0��w��q!����n���p�A�1p��D�-ji���w�Q}�~��3��8���WA����}�<�D�ϱӷE�0�ƣ�1�����X�ϼ�f��ej!E��JLx�=D��Br{��a_��cK�o��b�	���Ú#��Ö�����dgQ~]�p��Q�?D#)�h$]�<;��
�ry'SΟ�����s��2�k�k<L�:1�;z��w��~s���/���F�R�m�����b���H��'��Ŏ�;k����Mҹ�
�oU˂{����ư�ƈ�G�iX��	�9IH��1�A͌��w���u:��
O�����0D��w��R�ؔQX_��W�2dI�>��	�e]�#�4��b�[�l󫴋A�q �[=�΅YPC�^n�:6�y^�4�+\I}*����fpA���~ph��
���b�n�a���f�n��`�^��|ˤ�(������tӪ��E'����lO��S ��YR�mM�'��%v���ٱ��)����A��)$�q��/�ܐrc�����,�sD��O�	�F)/����0�t�{b���̦J�'����Z�W�2Y�"�P&`�+u�~nպ�sӜ�_�)�]C�k��l�WD�6Ml��V�~����4I\�������q�������B�uK��2qQxE@�޷�x��pD�2�������Y�_銲��^Ȉ�f�o��n����������?̚�I�!B1n[�5{z)ӗ*9��/)��gy�n���
MC��:��b�Qj�(�`�x�V�u�Uh�>��N��� 3�~��aB�㠉�y`߶����@<H+?����!�p�ݸ�6�<9綅��0��@?@3ѓ,�Ѵ��%�A+��yc���S�UǓ��m��$Hx@�$���A+�2Z��Qp���-�A�7��
��/�)�Y&�B�$�S�C����S��Zo�Dp>�W.M�O���J��`E��(��E����d1�n.�|��q6l��x�G��?'� �,Z�}~�p9��]%4�{�|x�Ϸ!o#��)�MVg�?��ǋ�L]��f&3��,Y4g�VR�>���(���(,�-�#ɛW��Ú0�f^+NIkdUF�q?Ů�1NS�����"�!�^ m�krB&s^�N$
��H�Tm�Տ�v��FV7\i�1!�w@����@\]o��/9��Fe��Z* _�rJ��,��	 �n�z�K>K��9�"r�՘�H+eZ]�,�oSA�)�w�N�>�p�����e��'B�6$�|6��MD��(Ԑ��.J� ��
�H�}1�I�k����	�}�.��-u�C��t���@4�N4���j��	�=á "��LX�;U�)�itt�y_-�E=
3g����U�w������	�Ht�V��d���1vI�}�ج�(t7|�X�^�@�mm�����(ХYR���V�Rj�7J
��?1�9b��؈�U��)�r�]N/͑�R���{�{�d��ή��6��U<�]��D���p�G�?1�����y뷖-a %�w{�.�x�0z��E�\h�A �,$8k�v@�2h�6I��AeB���a��_�A�歏#��/�$&0�(�J5�a�}�����������vM���2<!R����\�k2vB���:ҍ�̅~�hk��	��Y�7K�B0�	ܕ����o�u�����Ӿ�#��NG�IԊ��t����mQ5%R46�B�O�^���/���Gd'oׄ��͡t)�R2w�/�C?�}��d?i3���;V�7I!�1ʄ��5;�ӊ�9';q���D��t|)��!� �~�� j�����n�7�ղQiֵ�Q
R�<-��s��䰦|��\%,vXP,���J�z~Hڎ�.7�Yt�r������oƂ#HVa=���^xB���'��xՓ�X�i,H�M��n�X��Z�S8O��@m�3��Zhॼ�@1����]6�qr`Af�n�`a�P&�@�
�P����"�����Y�����~\��<oLl}�i(d�1��"D���T�_�Q߼��ރ�D�2Ip�g������jb <��
T�{� ̧ѕ�
����RW\P=��~�J�l���wCp�R��{i����+���d\��z��Q��7��Կ�"ڟw/J�>��-`٤�q��:o��h��X��w���ɼ�#�������y��+̝���(�������=Z�|n6��P�_̕����H����Z鴼IY{{��=(g�C���l���1�����y��*���K�����D2�>N�qG�6��0�n�v���Zy�+
�`�l�G{��UN�j������%]�>��������o�%�L��tp���!��{�cw��!Uz]��+?�#�u���jq@�U�b1��S|�m3]�rpK��+�^��.�T�T	,B�Q[V\6�W�B��2�Grsw;G�H�ﭠWv2����zެ:�����]N�&���!��H�xˬ�����l;b��l��k�HI���Q���.x雜d��k�t���1��[&�m�\���E�g�&�ɷa�Y;a;;�~�^�״��P�}.4�#�ש%_�V�1)G�F5�e�~��<+̤~o���.�>Ϋ�� �W��3�_�k�Q��{?��l*��)Us�ЃM��x#W�7v̼�i��j����r$�S/a3.M�5��:�3��K/S�cƦ1�'���8�&�����:!y���gҟuͻ���&S�� ��úK��
d�!:bWwx�l�^E�p�@؀���Ay�+9=������H��P�VC�*�O��j���@�"/�`�?=�)YU16��+���Ek ���;Ӂ��o��2[���ձ⭡�$���Y��*�ÈN����z��/�iace&W�@��0����;�����˅���8�#W,GC#�*i9:O�����y%�������H2�ϣ<�'v<�����%�Fk����m �����-xq�Ӈ2�QX	�y.&�K4�R&�ξ6����3�r^@�+@���g����s%��ش.�R�6"xz��JNTyC�,ɒ�d c�Ff��\����/0���۩XU�T�!�|��V~�c�Tt��V��
�}��Ոе��)��q��(?Urr>��ob��Z Kgё���ô%=�0�X+�|<�ۣ{.K[�b=`����	��|d�M���	��'۬�E`��;��
2������u�J�<1��Yy�I��0��T��Tv��f����2��.f����d���L��g��?�8ȜW�/ ����
Qfqx��W�ڮe��շ
���[u��Ѵc�?�}�2��\����J̃m ]���6iR�N�e�6�]�}47�$��M1
��k"88PK�n� /�\�c�?�&h�Q��~�4�n�v�ƿ*PL���h�	Q�z��|y��Kr�6Q�W�3�C;�d�=>�1+��N�ܒ}�-!
a���g���j�aL�� ���L��#���P���`Sl4�H�M�� ������VcX�Ey���;�$o�s]G�m�=�_�	Y�;��>#\�y���3�TE}]!)ߋ�2��W�3hLU��7�����s��
͉�4��&�<�4ڡC�s�&<ub��L1�m�6r�wꊢ���˄6\T�ԫb@��J��뤜>�a=E/<���x�����%����-���p>���WVad����޶݂C����,��!!F���������I�Y�Js����R}�l�����q�~5|Ҏ7=��y1�>Cx���v*�J�e�ÉU���}/�8	���r�M8ۉ������:b�ј"���ڐ��;�Q~������?��-�5=&=ʟq���?jX�q��Q��7��z	��T��P�'�4�K��Lu����gR0��e�QP�f��KW���I�u��t���J���#�N�������\�����Y���0�MԾ���TN:���_�\�ǳ���t/�t��/Ν��E��\��HZ<M��w/&˾-�BV�iܢ��@�x�86��^��@@gC��<�ꗹtb��Y�f�0�n��ꑚ6	���, ��<�YXM6�TiR�l3��G�I�ٶ��� ��ۚmf�h�������ߣ�#��(���?;�s2��~#�����7�#����OcCG�B�����ۻ�Wi�:R�ފh��;ݦ�N٧��i|��-دQ97��^2I�t�ڃb�j��;��*�M�C
��	��2H�������h���IS�VS��ʕ��c�OQ^�w|󘗺��й�L�T/L�N�e�v
D���ǣ@A�F�2��nraxp5o|,�Aj����id�$QQ���8�͛n���xu��Z�佑含��d�3���̲č]5�`ul��슛�v.�󞍿�c��E[�'j��Q�Wt�����P%:�<�w? ,��|��87��R�s�4��Mo_��F�����^���'w�(_�L�v�QwW0ȥ��bq(�O%#�v�*4ij���RAl�¾�X���������ח������*��b,E�]��Qe�Z���e��c��������Da���=��	�};�����|K�u�;g�9�xa�%K'�?�+둸g�Q�g��G����G��Pm��'b��*�%E�gL J�h����Ā�����`u�'+c�n^Ӱ��ЬiPU��_��bF����O�ԞC���#@��Ъڸ�r���/���ǭGX�'i�А�Ie��Н;�+��*����0+7l�ى��w>���u������;��<7���n��9�5����:o�����=��Z�����)W��	�t��-�;�T�BN��)j�<�{�!F�F�@�AyE�QV?#i*�y��^t���o9���)��6{��>��]O1)���Q>�!���]	�Yey�,�vA&`Q�	Oх�����`�
3���P'&�S�X�hN~��W����2�s��ӖXG�$ㄻ##��]!����b$�u9_��q�̤���W�"8�#D����ǌ.�
�N�^�4���{�d&Ң6ހ`J�wMi�m�йMan�j�_ߋ���Z�DT����!��U �h���ףR&���b�Цy�)�D�VN�鑚�h�_�9X>50K��EYNT���^XCdAt�6�R�4WF�<�%Y�Ltj�:4��Cs�����%�~�!8$ol{�j����^����b�xDES^��!~��	�2�_��,������i�������75xqe�}�P0�,�/�1���Ñ%�W}�z��uf��@�-�;ūd1�h��r"��w3��\�<���*�1�1�u-~�����ʝnz��D����f4F}g��ayxW��O�d�.���&��.ʤz����$�����kc���گj��R4���Z)��J	H��W�>q?��E��ݙ�a��;?�P�*g 6x7H�-���������}w��7����� �
2t�[d�/�Eʔ�\�a�|?�G�� ��{���!<����Km$|gV&;�k�߃�
q�}9Ԗy��2�M�t���<�fy���Ӥk����8���u��O2��a�������I��r$`�qJ��qg����pM2����G\f_��)VQ���0���o�O<�'ţp��ٖ�ǐ�1Z<$��z ���w��t���gȨZ�[�4����<h�K�N�q1�x��6�ݬ�5�%ڀE�#�3�6�ŭ�JĆ�h��w�$�-֊Q��Θ����7߂��G�|��4�a$|�.&Ǟ?�@�$������:}MAOt�B�|w��o�*��-�J2L�1��!$سyq�@�%T@����	�2x��8��P�#+D���N\��"�n�0�C��Ï��$So�^���`x*��%�E���f��.��A���\���_-m�i0�6&#}�`��jd���ц��:Ǜ}CL�1�������u�M[{�)�s�1��O�wCJ�8[V�ן�ۨ��x��Ѧ�`�^�:�$���4��X���΍��M�4"+*��cV�r��?���h��U��9�G����K1w$,/�H>݃���x�Љ��`��(�]����M�G8�v�4FZİ[&�t$��v����f>dD�8�r��2��~	�F8BO'o狗HT[�_\M0�cr��l�����=?��������xJ��nE{Z�P9z�UP�g~:0\� �X�r;@�~Y��� ��tg0��1?Fց=��.��U�+ק=Y�������[\	&�Ye���}�Y?$�VҖv�K�{�).e�'��E ���Bՠ9�E������ّ*y>��ol4'C�&$>���:�Uˑ�Z� �O����&�uT+���Ÿɘ�n��g⶷�����ƅ)`>o�k�?}����� s�(��
w@�U���}�R��4��٩�lR���ݪ1�e*�(��p'��R��m�U�䱎?�R�rnL�4&&=�Y��Oh#@�T���`0�����܏�H�H6����8Fk��Xo��PPb/��5�P�[3��7�f5��5�F��k��8jx�����Ԭ��F���D��r5y�y�ʈ�Jqf�q��c ��o3�0�F�>��=.bd�9h�+8��&�c�a����GF��:�j��WO�$'�^���v� I��l~���I��4�����>���>�V_�&m� ��)�A�2��`R��*O�qӪ�HJo�=����2�F���+}m�B�,��jǽ?�]�[+���Mvʪ��!�V����8�rP��f���T���l@�l�;���B�d��� �s'�c�� �*Xѥ������bY�g��I���i�O�T����u��18��t�>����t#���k��n����+_֐`^Bo�������m,��I�>�F؉3C��5+��9	k�",5���4�o>�`TOs8{����?7�G��0g�x�0�j�&�6�$���N��Ho�ÍY�رHC�*g˥�Et ���0)��'�j4!yV�M�P����gL� ���+�Yڙ�����~A��[��f ��cv\>+"{r��g?
PZ[G��M��9��kQ���{1������f��m��~^9���KA�s2� "t����Qhi��A �ŷT'�;eI����X��z����|ٸ;|!��)/�"{�i���< '�?bă��ˬ�*��R"�%�g�;�)Gi짐��&� �*��~�7�-LɄ����^'��4s�,XZ�w� ���1�m��].���&eB�u<��d�M���F{%���,j>�X��M�Aԗ��(�����G���g	`�Xz`o̟(�� !��L��*X$^D'ʑ��Yh8�Ɖ��q}_0+3˜��2�ǚ#��m[������9�q��_l�3��0l�V}cd� �� �{�/}�5)�o�[�2�oR������ӿO��$V�Ic�b�����)�7��{i�8K��!e�%�&�(˩�;j,x��'�XL���Y�H�'K9V�@�*%�D/�#���tp�(�����a�HXٖ�(;��ȗRg�d��s>c�8�Epʦ��*�.iU�8����� �2��͖���y��Q5��t��ſĖ8�������֠'����Ǖ� I�{$l�-<���m�p `R��@J��H�2w��[�r� �y�b� �eҰ�`�-�]�6�&�P��@(�ݖ�$����pϵ�p��O0V�c� �)�tT�[HMܣ��Q�%�P��:B��g���E~���+�e���o�+����ӧ{p�B(�vz��u�i|��٣#WhH&@'�ŽW&��Ѡ�X��"��׺H�
�
�0r�:r	��H���j] 2Cg��DH2���u0(�8H�o]�-��XX� �Y�؜e����P�yi���s��%���wW��Uƛ7�l�ـ�hc�ZYUd��MaS�w�FI��6kR�z�~�zfG֋�ߥ|;F4�	�n�%d�K㺌s2��!99ӹ *�!e�&�b?�|"���[��-^wߵ�;D"]s�u�Tbbl�:��i���
s�`)�,c���v]�ӆk���	l��;h����՗~��4��q:��*F�9?)IV��h��ȼ�3��G��q���=��o��	TcuOK�T3w��$r�
�e@n�E ?�g�x�X:���KN�4-1�����E#K=���"96�J"�� �b[)�@�T���B�J�P���\���>��1�p1������������k�B��]Z�nIw��yT\�ͥ��Ӡ7��F��=>������O��IH����AT�P���h)�R��*���u�K���5����H�Q���s	 ,n`i��81:�
��J�dm_�B�Rpii��,�Jr�,�<�O��~?M-k���$e�A�EV�
--��R���1>F�pïr�A�!g"��A�\�?70��7�@@��B�b�ӄ���:��@]Bm{�I{��t��$��q��-A4��r|�6��q�Q���dPo�FA�7t�ZXdqD����u�P��s��W^�����]�]�c��x
L`_*u��[�^c���d~���l�*V��?�0�[oK���CV��a��s7U��DKj�\����q_6�vDj�����FX$iF; x�;�����5n�q_ZP4�m@�&40� �s�7	�-�s�owHy�G���|�٢���2zeB����	�6��w�{�L��O#��hPe��ˇFmۄ�m�o�v�-���x����+��h�h|��T��tf�)s�q��LdJ�m0��-R�&ٕ?��,�":hJ`8����<ޖ@`��׾��.���"���]�:�f���b߁,��vMsǏR��9�hc��ͱ{���
g�y9Y�fdh�|#7�N?�� y#�/���.:k�RҏG�� ��UPf:N�Ic�m��z�����͠[���(�=��c_�W�Ԋ��{�y8ɱ���[FE���9�W��w��A��/������j-=��?��VN��)��(�j�DP!�u8���yyc�ӟɩ���R�3\�7���c%ZA�0��V>r�fU��� ԅ)όb�����G�ago�V�۹����k� r��Z/�F��igOv�{&ox�
Q���S1�k�2+�vj.'`?����&�s6ꄽ�吤Su�_PC���R���`�X�e��aQ!�m�) �q5��ɜ�*6	gT�s�sx��r��ʍ�w��2jL�I~ %5���l�����h�Ru��o�Z"���t:U�v(�Ȃ���Tn�ߛ�e�ֈY�v��/.ĿD���k�P�u����܉]]^ҳ��8����ܵx�?�����������j��H��L�s(�M�j��[�|���v$Cfm��T��Ь~���2���߹�HD�`�/�:���P��wt�L�K��F*H����j95������I�~/&��DFY
�$���Ս���R��$$ڀ�8�֣�
������� ���& �T���qnD&���ra���@x�`��*H}|�^��j�J�7j���, �11�g}��R<��C�a����K/����e���S(����B����0a6J`����C�*�~91v���4��v��i`ˉ�m���W��'`�JEo��)�GF��=ϛT�AM�`j�{�&,�+R7�1���_���ϗ1%�P�Rx��|�45�Ǻ.F���¹�$���W�Sj+V�n ���O1��q�GB~Zo�ɗ�;��q�	:h��SKN���V�7�Z���LU-�x��|f`Z�No;'Q�	CB��*�-!��[���T�3����$���+�%��b�ۻy�ɷ�yG50h�Z]���!�����J�lZ"��L��(Z0�7�ٿW7&�| *_��>�&F�{�'(�KA1�(�8���)�B�1�@����S��=�~�ᣦ������?p����0>N.��E���$����r�k��ۮC�iE*B�6D��woQ� ��K s����m�� \�"���W�X(Ǯ=��,_��J��1)�a�NXM�����l��4��tdF�1�B;_1i�++3��jΫ*���j��۴�� �๬²4����ZϢ
#e�H���਀�/r�y}4�-hx`�?���wc��K�������ř��E%��\�I>ѽ��"�����L2�[8�D7�E,���PO��0(��]!ٰ����ٙ�)�X ��SR[�uV�Zo���Y4��؄�9P�r��p�V������r�冼�T"�|YB��B?���}����q<�۟�U�*7롂�OL��aX����cm.<��6P��"�ԗ�jq���wcJA�ۼz�eTB�l#��#T���>Ǡ��	������]gIs�_�X�$it�������y�\u��W������`_�-�srL36�>�,~�Wj7�at��>��� I_���B���%�K������y|j���oWI�"2 }�o�����V�,�w[��C���@	φ��	���
(�u�:���bw5�
�����J2sJ))������,F�1\���T��!G�8�m7����ηX6�Ȼ�KP����{�-;��p��R޳!C�tI�3����
d�-���A^��z>ɦJ�������V@��> �
��b�4ON�(�$�'�u��T��0��/B�3!bZ��&�A����Gp���$�-p����z����~QYV�w�9�`T��>�^��Rk��®?J��Wg���:�2�i����"y�'���w�/*se3e��2���=)xЗ7���R��@��~�ި��=��\����#���T�� Ł��p�ų�hݡ��?�nJ3����9��_�Gޟ������+���pC`���̲8�ӽ�;�֖���=k�>]iGQ"�z�z�S#��v�a6�O�gHeV]��3��KMN�ez�"Y�-� �qvo� =��J��X	>A��`��:L�AOޔ������M��8v��}� r�ֿ�E�����C\�I�{�׾����a����PM����j��N�mx�*r005ur�f�u�ﺪە�����"|?4	������b"רs9�,55i��!4�`a��/}��C"��U�ė�u��稛��0��d��JA����l��h�ML] �X��פH@���Cz���#�X�sb���Y�\��r_�����eY��Rs���������kTE�_e��7�9�Ù,�>�@Y��+�\ǳ^�y ޶|�4�6��\X�h`ލ�0R�vr~��S���ך���$@	�FBM.��\�ʁf�8����5Ch:���,��"}V��w���r-��1d�\���S~�1��i�b$���B2)��c��'"��d���6� ƈ��aj��]�rA�1z��7O��N'�g�2&�AS> !a%�[7�8f7�����5��Okf�_���P/5��;��3h�����p��	%�����FbB[϶��ZçԠJ������7R}����C��CD=��!9�����I�J��:(@p!�6�c�\�7g(O;5��l1�UQ��V��?-���޲?��ǇZs(��e���V��� i[i�ϖÞ9u8)*�F/ъ�?u 3�4J8��x�ە@��;�3S�vP�лޙ��*�0��1>�����!��|5�L� R����0Έ���Pi���P��V���E�jYS�sz�FH��럍�V�c���Zd\�>ϐ�Q`�)#>�ҙH�>�z��wC:8I�s#VL��T>�?�e�����<���&���^5ä9C����?��\������@�C�:�о�SW�b�Z.(Q�i����7>jS��r�� ��Qs��[I���l�B1C�l�\�󭅷�J"��?���>�.��,i���3�zw�]%���v�����|b�[ea
��6��8z�}-d�$�m��}�e~��TR�$92J���]pJc[`d�s�x0	3�e�����^$JWe�g��JQ�-x�8m�3Zmi��{�.�b8�:�K��Ҟ�^�a�4K�؇y<*�#���RG�룠�W�?�zW%�����F�4]�.�'�a-jCBУO��+�RR3�c��c���pG|�de�{��UwK�&��>]J�+�����$3�O�4����7��8��D������+d��B�vT��u��ܮTu��㑣��0��+��3���v�3cZ84v�G��w��v�Q��W�+��-��0�}���W��ɰ�㓌�߿�c���ݘ�jmH��>
����֐����ݻZ����W�>U�[^Ԣ���L���Th�c�[��[4[�7KP�m:E�v�K���i�!��]�5��qH}��>OQ��>�$��� ���+�1�d&a��:V`�K��������%���/�ȡ���扔̷d$��z8� �F*Tc�	dƹH(�W��>�2������j.oe_��`#���mE$hK�.�C"��t+BR�K:

��s���g��!j��U�ǽ3��P#�ʳ���|U�|c����um���^2 
ŕ!��YL�k�\j����g��3ͻ��	�n��F��C*��]�W�$�J��q�$�])Yl���HZ����~L?3m�"�������ќ�ډLm��5�&&�R�r(�_t�ʇ%��=�p�98�_F}��W�oP4[��V����u��M�(t7�r=B�<,��'���M7��j��}����j���������>�cs�p汹5�Y���>h���и�62o,�΁��֥�)�W�~X�?I|׳tA��?q0�V������o�����>b�l�6��f2�Y�,B��Դ/XA�*'n��_n��Z����=�v�PO-pV���V��-?���G��/i	�EV�m5�YV��닓8�Jc��ca&��N��5�q6�F�Q�YDyf9�J���A����H�@V�w{O�ҢlRŽ�^��B�`�}:C�|1Z��,V8��e�n&Z]2Sq�G%>A���?�$rjۯo��j�TM��L��2�m4���彘����Ӹ̉l�5��߭E�.:�1*�H�]�2!cP�����~we����[�Ӂ������/mG:IG���R�R�������*������Je��O�#Hn�;��6�o����O�#
&y_:��u B��'��k�I1+�E�6� yK��aZ4��f���tmh[2pI��/�d@��F�B�'Yϛ��]��E��D���XZ���/�dͽ ^��oY�X��'�8�̍�L��ZSS��Jɫñ�r���ϙ$�O��Ψk�v�&�_�\��񭦦�1�O2i	��@�X9j�Q�k\ _xH;�7���6s�`�[����C��'�L��|7��*ͅ�������8�\\sP�B*ҕ׈L���h�l�9�����M���q��w�ӹ����sl3ܒ�V�7�}O�ij\�D��y@����O�"��1���ѕ���}�N��AӒ�OYu���n ǐ��e霘��&iV7��Dejn��դ����,h��m�Ϧfa	Jw@D�EW ��'s{H"�#yy5����f��k��D�L�6�<<C�a͊��W=�&d�am<���{�����
��/����V|��c���o$�ň)�,Qx���y+�P��fZ��{i*P��\9VUo��֔�'��\g=�ܚ��$
4��Fl�z�������!�ey�M핛�7�h��"2"p�������m�F��"v;�>�7S�.�;���rzHڗv���9;�Uv�1y�T#̦֚{����oe~�(|-����Ƞ~F�?�õL@#���Sm�8��]ؖ5�:]��,�DA.e&ri�8B_���f�Bθ�	�B�^���Q�D���]��v�V�k��D���ŋ�,@.��Ң3���W�7X^�l��^w�A����y�ߕ�U�&��LX:#�ZS��P���[����@�v'�
,荟��P�S�&�}���j��_��,�sN�́e��ӣ`�T���ahyP4X`�}xDS��������U?o_���_�q%�d/M��4��.�D�6ʺ�!Ko�|�%�̾л�;O^F�i�+׮��	�����j{�shYA���Sp�\��i��+o���u��x	>��0_	q�TE"gǄބ5/�oK�!Ut.(tjG8U�T�D�狹�##y������z����$�mG�U[�}�����D�T�nZ*M6��쀞�gs���|�_�d��ӡ\e�6��!<*��b��Lq	����gw���)�#8��t]��1�lX�G[𕎯+׶������e@�"����
e�%3���,n�Gs���Bu�9� oC�"�;��{���x"��L�vhQ_� �F*]	�)B4�&���(�P��@+�3� ��v��l��~X.�u|Q1 �L��L|w�!߰���1X`�(���S|Noε��ZN9��$^�q�%\;�J�O���X�1�~�3`��r:g���G��!�Y��+�H�'�E{�FK����嬂��^��h�1��jF��"��
�k6V���Nخ��:;f��d����pӲH�Ys���	�pվv>%�ڎ��~Zb�F[��od��p��{�q���=���Ǳ����?�]����!��Q�k�C�Z�;Kd�T�c�N�[/܁d-�G	�
�nb�w���������l:�����!��2o��Q�_$�P���9�9M�N�Ͻ"�:Y�൑�"�	�5���l������pꮮ���q��������������.�/�;�� X14�3���?�tm�f/X��5�ף��T�N����KIe�Pvh����Y��4�<ws=6�^�g:f�ݲ�d��r�c[ ���V�}Hl��
��Nݙ������,gq��M����aF�^��<u��Q�N i��$�K�m�w�Շ�ٙG�]�5�GeՁRV���vjx��c�Ϝ�����74��.��N��ȋ`����֊�ek$u;�j��o�MG��F�E�}�h�.Q�
��	��ޥw��b�#{���M( �7�,������}��b�/w�����op�7DQ)��f�&��v��M��YEh4R��r�Y��GO��;�
ϑ�l�ӬN.�7I���%��F�"��Z�w��Ⱦf��)e���e��{�$Y��jD��o>F2�u�]^~x�=O4ǳ
v���K
�[�S'I%E $��y���w��o�Q���;ЁsE#�JN;)���x�U0BA��k?7��S�ʩ��ݫe`g{v���5��4W�?��FTC}d�?ۄI)f[ `�ȼ{��뻾u�2jX�1���_Q~$��5Pl"�CR.g)w
ln�B����?���Y\����j5���=�u��}���a��I��#�];K�<Y������.N���)����">o�GF��,�i%@^��G��^�V�2��,j��Q�T���5R
�i�f͇F˻m��[�gg籿�K��eX)+�k՝��~��O�������t�L '�G~b�0+�9Xj���3"Nj��:�b����i�8���j�Xq/�����*L:�nD�)k��s����
.����L_w��{N�7l1�݀��/d�Q@!2�9g�&���Fz��Ӫ.�W�%ӹ��.Y�Mt����ō'}�k��Z&U�h�� ��O���ٍVݡ���N�|J"�,´�q�-��ʻVKhC
��x7��F��q��P4X�ٱ�3�	v&��<�%�#�(��H
'a �>�
c ����=ˑ,H���f�DQ�$2�����hw�g>CA������tK�?#j�>}��*�qs�0B��?�|�i�K�ޝo�,�y���e[���}���p]�g}�z6���ǁ��Y3����1��ī�Zm��p!%� Q+J���"(�l';�t'<��^aO$ߎ�F�fp�ty���E�^t.��0aWd�^fc4��{KT����y�S/�j�W�"/G�v�`��^��8��c-2v�S�Ų��.�BL��$�|JX�6뒟%nP��M��t�(�-�u���>0������ ����7�|zn
*Z�q��2&�j���Fp���ޤy9ό�V�8'vr��l�y�;"����rp/�8ת>�Q_��n����◷ )�}�����E��6fO�Gq6�[�l�˰O��ڠ��'�A���pi������6�d9'T�p`T��W�+�z���K�`�o�<�<��_N5g�*���У�TG;q��U��}B	f�h�>�U��k��N����]g%*^U��v{��ind�&Q�/�����<���¨x8�p�}�2��;^������U�v����C{	=����UHk���|�>��ߏCXy5O�ܩ,���,�㔭gbhI}�8�@��u��`�vA�F�-�tG�K!,�(���]�p���̷*�=�d���rR�2���t\�)����a�̸g~8&'��%���p!�:we�������	�䚡���q�b�Vr�S&M}�~����a�X�?���O�������*�-V*6_n�	���x)�Y��I&嵬��~�>�E�^�^κ����K�f���2�Fk@��i!h��h����A&S�P�-�Kt�	}��+��!��k�j�����:�JBq'���^=Tq��U���"^=0"Q<[m�j�҇R�/�S8���d�X���j�Y��bb��EzV��l�<�f �\�P�w��7������V(<}G�\�6u�O� �ň�~��B٢�$���p��2νCw9�/6߇�d�.q�y�ǂ�±��Z�o����Vk.�Ў��o�����Eu�����%�ݙi!r�Tmu�G�����-��tB�f0���%%�T}�'�Լ����|[mC(�r=G��4|H��I�χ�pd+w@���*H�l��^=��w��^�胢�d��7�J�&�;᫽���o�/�M�����1̯��[X���
V�r�-`I+�U��Њ���2��/�T�d��3C}��>��cr��XKȬ9��.����Iyz%��a/i�b{��9�@�Zޛ�P�/&�-��N��Vy�4���r��g�C��3u�I����ZI�Gr�/Q���[yq��5�k�6��~����א�H�o'�wv�%�9�e�����(��V�X2��>�~&3"��@�9���z'��q��h��d�)f|��oߌ����f�{�c��Ѫj�jVp����^Y��G����Cq�䑛\��L�	�!�D�Fێ��=����ڑ�����W�[�
IfĤ��jp^�.�����(4�p'0�~"�4� FiHQ����_���C��Af��+�x�x��um���kw�����Ve�����^��o�g��f׻z��̅�nt!��bv�)��� ��x�t����D�E�H�L�JJ�G���ѐO��Yr)��c8A���&��b��agw�*�`x]!�d{��1��Wn�6#%�&�chwυR�uF͟���R�hR<���
�O�Y�.��Ǟ�`N��cRxk���n��-�]K�O�;��f�������1ΨS����֘�e��4�k��O"�^7T]���Ґ�P�'�~�S��r���2�t�6����A?�L0L�@�_eGs����:͡%.$@�ɚ���F�[��r� h��rf�ߵ�����y-��}6��9 f��<B�	ҿB´S�����]qȽ���!M��d �	:l=��M~
g>6שli��j�-��r Őe�r?��7G���o�s1%���-}g	Gm����
�k����F���`j�M�v���D�������D�/�5�"6���8��/��xJ"�j[N��҉�:L�~-!��ZZ~�Ë�|@uP?�ܜ�^�ًf��Jko��R�8��(��y\�;�o�I�}A�W�px�@ºP�݄lj������S�����Q� �F��}6���T�8QM��~M����Ebn�0�DW=�������n	�7e��L�w�o72-B�k&�Xˊ��v�x�\�ԩ(C�I\w�
���$<_WG��D�{-�f/JfI� o�f��4�	j�%3�O{�$/���.ݬq#yg�{v��/�d�w�uܹ-K\;4O����{�qu�vq=�G]bF��l�%Z�#��<���	�����mg/�z����$��f��u|"N��i�̀)�O��n]վ��P@��t��)�@� �F����.��o������������e����@�c�ղe+�������`R�ʓڨ��ܶT��Or �01��A�(��s��2sS�J��OF:�i�ӾLj'#8F�3�4���z|�ÀQ7Vz���]���a��	D��G9������YE�4$���Wt�`�Yac����ko�	����u�0V�����~�3�V|茞g\	�V@T�7��t�h�����co��1��<�g��J��\��ةO���@ߤ��:كh@.�*~x* �r���n��؟��cIb���37]i �4��;���44�9��'��şG��;�=j�.?��*���P�1 P�ED���S2�&?��h`������F�d�����,U�r��B?-���
���2��Q@�ԿJ����:��_șV�i}�s����9鯇�d�� y���K����9��/)�Nj5v;9���>DΕг��c޿���*�9�J�XB|�͐n����j����:�Ȁ�b���R��̭�w����SoՅ���sh�ꔕ,h�ԋ�m9���ӸJ��W��衧u9�����bq���)=��A'�-�F�5����w�p���W�/C�_� �r㰵�&��������pD���^���U��rt��N�c�]	�8����z[S��)�����Ym�七�裳^��ak>�uUb��7�L�C�ϋ�S&z��!+����;�B���Po�Wghp�M�uiՏ*^�S+�S�?�DX��CvG��_׸FX4~*E���U<����+�9#�Cb��L��`۶gUX�wK[�y/5�Ǆ
z�ʷ$l�%�О��e��������J������?ɉ���!Gb�f��T����#P�i��g��3¾��Y�N��m�C-ħ6+�>>K�x ^�@1��ʶh=�I��l*���Kj[u��o <D]�d�kz(��I	3�$��/VDԋ,�1��U��W6�����{D<o���Kq��Н>i�$^x�}����������ј����Ů	n�=�d��X�}���#ɏ캧Y4D�v)����j<�n�^�eڵ��rw�<�0�^� �X�Q��c*�*�'N����n<͙�rF3r�I�c��5[�"3\�]`=����?��b+˴w��r��k�=x�B��MG�ۗp�U���3v�bU�#�W��L^o�c���+J����Y7��esCK��R��� oJ�(��4\ol�:*�&G�@>��0<MZ)�����k�v��|mr_;IM��qk�������8�y*TDJ��0��d�fU�����q�PՓ�41s�#����e��>'���w��s��`���:5(z�3�j[N[��`2A�^w�zTE"AS{���w��ӥTJ�c�<!0���� l��v�1��$�!�]��ːf̺��2pk�E%$L��S[66[�AU���dnkd��8-��|��R�*-�1c�%���U����!G浦�~�۵�uN�e�o���s��d
�F�֯����؍8X���v4�B�ަ�O��(�sd��d%$?�bݝQUm�3A	��6@Z�M�b�^D����FXE��tu���jf�;�e2~~�ң�'p�	ūoX�6�p{'Ͼn�D+k;VD��w�n���b����	-Z�zoCz�q�.�0���Y�1@�3�\����v�U�r��
�Y����[EJ%�3���3:������G�E��ޛ��?�ЙCL����V?BN�K�;�2~�K|4� �g1#��"�9ʹ����Ɩ���Lm�C1��h+V�x��=���J���N{(�@wL�B-�݇x[L���#��T[�9Z��j���V��j��*�2����d�`U�I��qo�=����
 ���Gz\��f_���"�
���V}�rە��<Waq�M���a�Q�p�4t�V��?�u�d��d�6�LdL���6A�e��#���P������({�rCL~�:����>�Ў���LWΘ(C*xO^�wdͧ9��c�2�����0�'�q�w��1����i�?CNuA���Y)<D��u�keŉ�����B1�,* �u��@��{���_v����ψCoE"�WQ�?�X��c=��'���2ê26?�cr70�Mh�tD�L�ʿ7���������F�	����\ޟtMT_�;۩,��͢���k�m��$T�۟�L/n�L���\�&�&�0�(^�P{Rzn�����ϗ�IAe��:ۭ  �3KK�	��>�%N�Mf���^A��Lu���5�O�)���%�cޚ��M��i�m��hte��ܽ�%:�cX5�3�&5�]4���l�̒�~�;p,+%p�BY�]�a=����M����Ñ�R�
�mNO���븊S����)<;,RX 3h�B�1#�y�f�6UmX�g�� ��h���ª����Փ �o^��+�6*����aw��r�U#�;�+��yL����p+ ��FCK9RH	�$��_I�%��5a����7���)�_����{ƚ���^2Z�x�d}xiϭ���#��5�V��L�l '�u��a��c�9���bR���������[��c�UQ!E]�Աgf���4e�k1斋o�Q���g�1�S� �s6n��^�d�6�~�-÷�[m_a�M���\��G�P���:���P�Y�a*7�Tx#!�Ҏ�:�jDO6�7�_m�r��;��κ?�#Q�8Sq��"��.�-yL�s���ћ!;!��,��l!u��> ^ru�S����%��Εi�E�1#CiY�����6���Į;�)���,��j��F��e��s�0�B2�t����b�J:�J���p��T~� N����9������(`x�����X���[p�� wԌ[�� HU��ک��l�|5g��,WpC���jS�a�S��- ��͙aӭ�0�n�"{.xJ��Q)��
z����|L���@=�h+ɈrB>YCp��1�j\��x�u����L\93��F�1J����*�p��i���T@�=��S�ߘ��l��^k1=��������eP����1�!@��oc�@�i��a���Z["�p�:R߃����SQ9��!�H����j�-��Z����V��X�ML�)p���nQqm���h��B%��f��),4SͶ� ��5�܉�xi��V���*�zk���������  �t榧�(dɋ�<Չ)���<6'�ѝ��1����Kl6W�$g��s@��*��ϸ��&�F��a���4�xz����u��XҜ&I$}�U�����F�R�F�d%�	rW$T �um�YJ&�X��tX�J����5��d��m�1w����̆9M�}"�Z3J�k,$�6U��e[z��[��CQ���O֖�$[ի^�-�'��p��������4�U�A�8����$_̅���L��sTt�ݟ����������7���MeޥM�a�Y�}��d��b��M�anh���K�V��\6�z�"��[]����y'^���L!� �/�AA�%*������)<�F����ԕ0-ԡ�%ӶH	l�+J��
�	�C�*f�-9�&���.���S�ARl0ɍ ����3ⶒD�kܕ|��4;Bp���'KY�E�rYJUt��/�~�φ��˝=��x�o��!s�Y�Hz:�Z�D&}+=GaZ����*E���8�b�����y�dd�TKFe�幌��@�]2x5�џj=��Nv�ZǊ�u�V���Nm��-�I��ܘ/3�\�4N��ۍ���rXdoDº+>�^dy���z{���`�#�����q�Nm?��Y�?�y���g$�Q����r�)k	r�#�ֵP'�B�u�'Y`��ON�2w�rBn��'�^�QW����}O���P�ȣZ�x��#�`�,����0F�*���
��̦�����+����j#Fȵ�dL�H��op���r^;��ڇ,$�}QP���#c@<_��o��]��P���4j������_���M2)5�[�3������d6`Y�Z��Ʈµ����O�T#ږ.����~R}I;���"�z�I��&7�����7�������ۻ�e
�>i�����{��8�C�2� �$y��:���/�7��#Ж=��]�ŪC#7z�n��&b&�u&H���W��r����V@�L3���q]i�R����Ef��jo+�!�}n�~Lw�oi�l$�{9�G�^�~[C�'O���X
�r�'
�tJ�I%ά��N�q����8���w��Y����M��ga��Ѣ��P����²���,"y��H&���Ś\��,�#��/�t�1�&��_	�;|6G
�����6%eYL���¾۪�N,+��0Q�F���9	 ~��݄��o��\�WS����r�>�QM�U�@�DW��K�;9~�`��NXl�ɺ�����6�NZy1��B*R���X��y�l4��HB��zC�e>#Z�h�j��h���Є��o��Ȅ'�T�1�xi����g���,I&�l�I����v��#�b� �M�s�z@i����;
߾�I�%1�d�_��ŭ$~Μ����s�X���t�����b��ӂ���N�S�L�V��z{?8���z�*��\��+�$W���skuk��$u���L�#��Ӿb�'f���d!������w.�RRy�D���o�x����ű�����m=��h���yk���	΀� ��_�6�|j.} m�ή��Q{�ڜT�#A�0`0QgpC> �08w����Xszȏ�vI�H�(���2nEz��u�	��cUHGN��c��� 7��QP�߰*x�f�����Y�_&��9��G�_�ʏ�	dcu�% �OB����o��~xQj%�����>>����9=ܶh���!$�`�z��6��>�v9=/ޡ����+8���v>i���!��؀��D|b��Yo;xM��\�GYM�+,uP؉� ��z2�{>K�|n���.��d��&��4țVP�s᷼�V,�J��l�41k�)Cn�M��������2K�i�^
B&|�E��-?p�ڼ)m�sij�%X���`n��� Lo��m�1ŭ0f��9˴��-��[2>�7�,[�}�����=Q&2�Em(h��嗕����-@�����Drr�)�DR}���<ݟ� e#B�U�)w�_]���vR���{[eW.�H �����N��x�
��C9w%�.�첈�/�;��8ND���̜͑0��p�#>�{�9!⫽��[�t�=�QI�z�$#�B-)�k��z��fa��LS���y1�j�b���0���8�^N�>A� ̻�	uԔ��L U�S[{k�Hƨ� {]��A"[B?�Sӫ��O�b��2�����ja�>s�e�E�͒���B|SI^��j�JFq�ay���=x�NL"C��
�ce�b��P��͖�@ù���l�$.R!�iiKN5�P���c����}-���-����m�9�7����}����˂�Ofʪ�Ei<RT�XЏI^3Q�*�lD���V�I�	�o��� eJ�Eh�0�t��x��=�& h��cxj�q\�[��w��5O�,�����ov1U�A)RW[4����3o�{�d�[�za��o���8/E˧:|�.�/<��E��=p+M���6��O�V���g�Ʋ�v�k�UZ9=�[���}u!��C*����p����v5۞�s��]�doޝ�2G��[`�&�D[x��S3�ڷy�x��˧&�k1�ab�6�Id��kP`B�|O�^g ��t0����W��btHjo^4ו�W�0��*��M~v�i��_�� 	ڽ����$8��Ot/��S��,Z�Ul��>O��z���``�x��R{S�9�MY�x̘�D0�c:?0&��X�'ؤ)G����TJ����Ɠ�ƙ"��$��V�\�e���̓ *9Ϲ��(�\����{�v �t%�h�h ����d`�����pG��N���ю��w4䳶��8��i�wT�������Q·�ɴqx��.<�\�^�,|�y����%d%��l��i��<��-H�:�l�c�J�}!���g,$똓��;��\�5�I"Q����*|eU���U`rlg�*�W���j�[S�$F���ߑ�h(XE�Re�0����]�� ªC��pB�
'JO�hfo����7e4Z۝C{~(n,$>'���^2BI���$���^���G����Λ=�ǚ��u�^�cK����R���/s^���uS�fL��A���^��( ~`}^�F���H�2�%_Xo�f;��vUrc�x@�B��̝#����~�$v/bXr�w l������I��Q��MZ�1/�q:�I8���|�?4��XK�kЕ�ϫY�mEЅD~���?Dl��8�|�	�:A`K�����U
.'5[�e����
�g��Ϗ}���ml��u�W�!
��f�b.�i=��k�b>^�6���(Q�gT�l6�̞��ω&{p ՛&͐�k�{�#���M���e1j���.9�����D }-���>Ƨ���V��~�L��XX��+%��v9b��å���E� �t )�2!��s�r?A�?�sU|���1����d�	ؾ��G˦�Z��8)�!oM.K.Bȩ��(g������>^���꽄2|U,�tXF����F=@��d�`�����\A�ϻ�o�r7�H� _� ��#&F��O��fH��ҭs娳�
�&�+ە�����x�>ĵ�^���l��)lņ;W�#��[�.0� ������P�Lu:2/{(c�"�fƽ)��_FRݼ���5�/wlƠ��i���e���Yݻ�B�<�F�IE��}\��)�a�������GFw͟���.����9T�l�Gcdӌ>��xx~�^�~���у�k�/)#�D#Z��b`ݭ���xȀ	�Pa�h���jE`�ӵ˹ƭ_�'�]��(���bp�}�l��ޙD��]'�'����1s�Ԉ��$!Ď�J=�%��\�֫`ͤ�v��7��A�9҃K&B��9'9���-��'��`�W�I/�̆SS�)ǅ|�4��bm������+:��G�LF���S0���H�����(B��+��'�S��S�kB$�Kx�Ȩde@Н�"
��#���Ď}u�CU0 M��b�Cm�H��lJh�ҝ�!�����j�ƾ�Z�$z [_�d����(q}� y��l����e�Z|g�@J�&:e�,/]��X`M���E7��d{d=�N�H1���[�a�y����ݨ$�e�X�FkHo5����\�!�*N*��J�$�$��f�*�|gż,�p��B�5��҆cBi�QmH�`��6�+>a�pl=c�Z�[�������>�Lx�c�K��W�w؍R���]��x];4O���1�`˃?D ��]���Ъ�j�!��G�~�7�q\޴���|T��Ѿg�I�3\����8k1�~^R^ͺ�9��b��uƛ_�qE��};<L��f�\�m���}���O�z�+ܓH�8F�f����@���n5۝5
0���B�5έ^Xku��q&�E�p�74�Í䵰Ob�՜��i<��G0����e��ˁ�v� 6xJ��H� ]��6�B��ұ?����sӑB���^�&(iUK,v��:���k0��V�1&ǌd�l;�oKl��Ѐ�d}?�v�*w�i�eq�D#�|�	��.�k�o#j�ϲ�)��ax@G>�J�\���ɕ���� �R��D3���ȧ%y�ۼ���̤���ˤ9�;S��I@U=�.|tk0*�J+n7)�.{�=�N���r��u
��L�<����$н�3	����n^*K�-�2I {l�5qI��J%��-����jP²2_��Xv�?�UĪL�?�M"�?�F����>�H:6����{���`<W;=�Ui�;���?��ޢ����Z���t�Aꋡ��^�>p��^��	�nR�Ҝ��K��G Wf[%:؅�gDc����!	(,����n�X�T�,��#D�u��wsH�9%W�Q�&a3�����!~0\A�h����rA�jY_Z��`0�^�}YK�+�)2h	Cq����!����o���e�#����@_~VnP�O��O֬�r�b��a�͞/K�9N��x���~S����L�Bg��o�iX�|�m�uY�@~��;�3�e;*�
�K8��:�U�.?����'MJ���
͒��Ѱ��56���z�����8����[sDHU�mBG�.���޿Q�:���W��=�)��w����#51{l�K��]�ɦ�3N�ubδ7Qf}���W.����w8Ih��`?~�p�'}Lu2#.�x�SgB!�;�W���=c�Ӫ�}��+"zp��\����n�l�릦�'
�!uS�����
z���mk�Y�k/P�U"�_���%�xa�f�,Ǣ�)��lW����4?kk
,GH�̱���;��X]��M�m���4x��4����]�r.)�J(ja���A��l���Pd��#�J�	��kkI�W/� |��2X�	�x��\`��*�U��u��Fh��(��Ŏ���QrY�Z��/�Ѓ�T��lլ��y�D���P��ώSdZ�]X�>:��X����CU�b��N��w�+��"yڙ�]�K�Wy��;�˲��rY��t&,H�mcI��4�{Ɯ�@��� N��o�e9�]�pϰ��Vuf74��Z��~|���+[	�Fy���HTW"%���r-n�}XJ��oݟRbX�+Q� Ll 'k��G���f�#7���=�;P<P��.Ͷzb���e�&݌+5@_��N��)ej��u@~Ch��b���+�8	q�������U�ހW��P�=�uGSF��kC	�f(�	���@n������!�_)�C��;��i�%��;�#a~��A+��D��Q���]����V�R��W��d�#�uxg��x���;�@�	��d8����cG���]U�A}����IȒ�б�bM�����O�7@�BU�5������j����Y�V�lAH�%ߖ)���@��R�u6��ܶ>�C!>���-�������V�q��6vt�+F��ٙ�C���t��.�R;�%�'p,M|�2���d���N� (ב�H�D"�t].�y��f��-Q��g�SN�p�d���	�����?�[���&T��t�"��e;���0������d�T��V/'7R�� �1���b�`IB�w���7TȽ8��]�;��.ק�Ȟ �h��)H������`�Qh(�DO�|O�x���mە��
����Їl��*i����N��巯Q�>���s=9��W.=�U^�pf�Z䖟�oҔ 	�"]�$$yt��r��u��M�cn�[�9��D����h�%#0}�ٔʟ�@j��s1e t<#��;�Y*���~�u��*�e��]~����a�"݇e�Er��J�o��~��Mä��!�͸jz�$*V�B�����&j��6 ��g�S*7��7O+��^B=Q�6��*�}CZ�I�� Gs
J�s���"�;�3M9'|4�n�<��kc��0�s�;�x��n�%E��R���+D.�JH%P����^�,Pܓ�����K�8op[I�p��]a��4;0Rg�K�� ��.��?�p0dJy&�U��&��cE����h��x!9+�V�`�m�~Z&�x��[�T<�pT�N����U/)x�{��A3M���_��U�C�k�HӠ�<1O���5�a�v��
�
�,E�?���dz38v$Ng�r}Z��8T��w��ޘ����E;/N�����.�
���Fw�x�/[N�����O�tRX,?�+�C]/L(�.8J��||����{w��𿌄�0S�����I�ln�4��δ��	�2�aZ5�J��&խ��8�3�47��Pi���-�&^�;R�8��=���k#�X���[��m!��!��dS��� �3�n$x���^QR��h�����s)kh>��6�W�QOkyo��v��K�u�7T��>�|r���U�R�L/Xݞm>���S��^���t��f�Z$�n͐)��p/ebs%�qklJ�SU��� �+ox�{m��� ^�enn���'A��rM�"l�ۋ9f��J�F:�	]�u�S�Շ��hh���X�|����
� ��LJ|�ir$0�g���Tg�@� l���F��˲��j�0[^�[����YӋ禜��J�做�5�ns��[|p�r��B�HP��eì/2�5�`����}�I���q��]��-9}fuoGf;�'�
��0�?Y��`t�ک�R-*�V~0b��>bD�|d�^�s�W糺,ʔ��pK��p~�%I�k7K�����~9ja��r��_��%p����m+F|�uɲÒX����	Cb�g�?b탛�Đ�ܟ��Sl-f)+�?%��d֩j6�
��i웚��� ivs����b���c��~(�ܚ���x4f�d��0̉CDы���F���^�O�PX$0�[�~1 gE0�`nk�[i\��L���g܂��t�V�ghCn��n�!hYt����3d�~��0%��{C�H/�	C�,��Q�E��̄c����Y�z�M����7���=F���!���R/�#PA�����=t�S��U<?
w�L�q��~�g�$��Ǡ�G
����7��� @��T俄T�"����4�����d��\��/�*�0���,�nd֝�x	�ʏI�P�>�7�z`�ۡ1i��h��\r�Ji�l��� ��t�o*�Ֆ9�Ϫ�j�H�͂g^_;.�������\>�n���o1��E��"|bT��K�)��!j�i���!�4ܰ��q���ٲ�E�_m�w-#��F��m�:���L*ڼ��[d�!2��M�n�N�V��r��>��&,"��6�o �����H\��*\9��~;��j�?���m���0���w����[@x��:]�]���h����������0�i��X���R;�:���i�X��cL�[5�a&�SD����Z�� �*���)r�R\�k����#۶�>rj�gO�bJm�r�7Na��-���ڜ���l�3�(�t�c�A���d4��nA��0�c����îTʛa����Y��HK���Ɇ��������8��s[��e�l3,��b&Q8�j�	Z����nR�lʈۢ���Py��hZ?8C�l�f,�� ����$�w�8¥�"T?���@:ό��x��}O��4Au�lug�H8a��
����YP�d�0�I)cѯ��)
cC��{#�uǑ,�>�5Koçyyq�"�a���F�۾u��=������H�P��\�Z#鎟�d���^ɽ�R�9�f9%x�DMv�a���(�Ϙ�/��0l��W7�ͮKt	E4�Fk3�x��c~05���ѿ4;Z�sFm�;X[�����bU5�`�m.2p�0L����0|�c-鄨�����(	�͝2$�0E^��b�3���&H{�{�)r��!��v�k(��2yR�?��z*�V����ns��D�aKU�7���[˪j~�����m���P��j���!Z?<UO�tn���.����zO���8*�<��-�����(����84�n�Md[C��;������,��b�X���zKQ���d(B�Fٿ ��h��}C�t�l���|L&v �\z�|�*�"5�wyb�#ҏ#b��
��[���4�/�W ];i����0�@*]�krF����)�
.��{�l&4��®0&,�Ұ�9+���i�{P��v:{93���w'�ޙ����E�;��oW�<�y��KN�z2�ʩ�R��f����x����ܮ��Z�楅֗�%��2Qm9�P۾:9�(��2�+2K�9Wx��\|DnMZ���f�au���W��u�#\��@��A,Fŕ;��9R���=N�2V��0&��%��&D�k���k�6�"����56�v�Y�O��)�ti�^��%2OlTK�����0y ~��$)�rH�ʑ�x?�4��sm�t�{���k婲��oFc��H�i�w����d9~������5�\�����:��$�|��x���t.��s�˙\�[���0E��wL�r�AZû���l[�q�%�#U�x�%�ׯ�^u<|���)���.��v+����B�<�
��Ҭ�_�_YN�V])��7�~� �	Oz��r�[!��|v;��ey��%�����n�{>߁_PJ�ם<�ȳ�
��d�66R�|9 N�Bğ����#V���b�Y��Q��F�[�3!C�\��r���ɴ[��A���NO��-gT�Īa�ϙsǛ���G�:s��F5oF.y�����E�C+�O����c�xa��YB����ӝ����`��[�Xi�S` :4����5=�S_�4�F%%�V3��5�/C0"���AnOsi�7��y��Ve�{5����o�����F4{�;��L���ZZ����@N�d�R�I!�5��Э��z���-�ζ�淾��:�!�neZ<��UYEy`������
�k��Z�����IF3�fyC8��u%Y8=�|�f&�HyC��{�fv��'���ƒh������R7<�=���������p=v�%���O�#��U�~�i➡�}����Jq��t���{~p����'ߺе	�#�-������~
CV��{8�*��*mDx���1��TZpd��j��{�����i���]������S�#�LyZ���KC\��C��)Z2�U��ǈ�N��Z8�c��e���n	Č��٨����6N4���(���G� �e�sNcm�(6�\�;L�s��%�v���[��g��e�M�c����h���a��o��[��O&&G�Idn�\a�b�D7��Y��8�I���0�~�bfZVnM���q�ֽ?g&�g��"%L%��)lr�����Aɥ)�X]�۟�������Y�km�SՎo�,�]�*+��*0`��j	�}4&,c�^��Y��!���$-z
��h�򄰉j>�Ԥ�K6���3Z*Sy0��!SveN�����_ )������sD�@��$X�ҿ_�е��]���P���7_�J�?� ��ôMY�dr�;,�x�/��7T9�<�q	���r5�u�a�VAK�E��p�=�$Ն=m��[��e���~־E��H�������K� ��KgA���8Q_=I�-����bty�ҫK)�������$J7���f`�Ő��Ox#����9�{��G���oV:�q�z1���x:ũ
Yku/syt	V$����N���|p�S�9b�1��}�;|��"�W؞����E�i�PXǉY�~�_�	B>�"� ���BJ�8Sͫ�P����]��Xee��^S�t ��,��C��0�GAb����d,�Jd���Y͢��Z,��6ʔ�e�Ă�/-O�Y<~T�����}�3��i�+���2$�M^����&�^U�i�J����Y
11�w�|Q�ǽ��d���k<[*������D�o2�:����9,¾�	\j��l�k�:�&79DnʓT*~��:q��A��c3������#Υ�JW���������P<Z5�;�_�����F���&�O����]%�MS|̢�b���`p����]a]j�D���}Ŵ�̹�D�!G�a��d��r��gra���;J���e��|�� BS��R�O&xB޴,���_O>�#�:l����OoL��,V!�����U�ȫ2���	���,�h~���m�g2���Y(��	[\	������z	x��U�6&]��>%?���nf�-CB��uni�*8�,PM*��I�K=^+e��X�cH��w��H
��U��_�.�K}����i/v�#�]!�S٦����I^��\���8��
%)�B�g�$�5Bj�N��-����,+~1���u����0
CK�_�N���N冧 H5���Ρ�v�&?Ds�#���m=������$Aj�r��֗$�Ѽ.Oߟĸy�2��1GK8:�W�l���l#�����w�� �����/�����u�a�`�V�	]zGD�|��`��;�/b����h�d�*�̟�8I$���ZD�W�d��^�"0?�&L�(�e	D�9,�h�<%EĔ��6@�ÚY����je�G5	f���0*j-���z�6���;/��I"C�ٝ��>�0�:���dHW�Q\��ds����Nݺ%^���p������@��C�i�$?���%�bY?����i�
tV��="�`u�(�Itm1Y�¢x�)_������||A��@(����Sb��D-[5~����"Sԑ���|�!�<���D����)�9Q���H��)��"�v\q���r�(��a	o���t�:V?s�v�@��?U��J��A8s���������&�y~�Ųt?=r��۠�9H���#uIϩ�4Y�k���H�b�K@�GRl�a�q�rk$�m�/C�O1k�?���Ν��4\}��yg���>5�xUF��G��Og\0:��Yq*��4���@N�����~�_=�j�^ @��S3ɫ�8ǎ���j BB�גanK���/��n���X�H�i͟����>\�f����K����(�R���Z|�b�� ��3��ߦ�{%��[�r����%I|[���{��&MH�%3@ao9�3������KQq"d@BԴ|G�Z)�8=�5��9�i4g�p�i���S��1���r�NB��+:�/�V7��i9�`:�\�^Y�&c�Y�,��H�;�{���Sy�{�P��ӣ2��}�"z���7^��-L�5-H�E�VI3/�4+q�1X�P"�T�f����ɒ� �Z����
����~�%�S]U*
_�:1��<�2F!���^�<�F~�e�f�.�1Uث=�4��l��±��� N��d}�k@uN��d~�ͮ�z���er�u�z33�)A)>�
��% z��L��u���6vX��#�D�u�c�����|N���Acf�8�Wl�ƕm���B������;�G�����L���$M��j�i��7�T�R8GG�܂
�/�F��_�>�'메���h�Ᲊ��9R�i��7h�䉇�Û��[�"g�k�>�z���>W��H]�]�Ƒ>%s뛯pgz �q~
��I%>�K �e�p����Q�9h4��Z$�%�UM��	b���Q�j����HCS�K�\�}B��i&b�a�VX�h#�$��e�V���b;PR�0�A�}�\�-5��/�(6�e;vO-�9jyN���X���X��=�m�VRd8�������r�o���ƭ��ߜu��'m�%����щ���FɦC`-?TQ��r����	B�
UۑGWf8DN��(>�������9���P��8~h�g�Hǈ�u9��9Ȳ�����w�Pw-��,5~RI��:���6�K(�"�d�Umʝ���<+�jTQ��Ϳ�"8߱������@v]�Q����Kt�����I��g��ۻr�D<�g.�<(�?q�n��'5��LT�.f�yfG+D%9\���Kڂơs�߿q�it��%V�E��ѯ����Xf]C� Ŷd*�-o9��1��	��[��P�>X3�L�j^�ʩ�[Y�t0C�ٸ����@�������e��J�c���	�-��@�a�l)%�"�$����6gs.�쭅������s���Τ��w�B� ŕ��E�]��*1 �:���\u$��d�������?�;W�Q_��������Uyuܤ��ނ�P���W�r��l�ɛ��<Z�Od�rQ��ӛa�����y��ئ�ɳ��gN"�����܁�ͿYVV8���ː2}�T�����J����hNxtiψ�"�/�_+�7�#^��� �7r�<�O�:����`������e��z�:�}1J����	:��<�߮�N'S�L��w�(LX�Qe�FU��*\�ُ��y%Y��1��)��$
-�C_�uwG����1)nj�%ӮR��O�dg؏�0|E�������$����J;$m��"���{3�h	9�
�I=�X��T-%3i���L�4��T/Ys$%�'N�lY��n��>���pw��D�b����+U���I� �Oo����ʃk�ۊ+5T����:�G�m*�0,Y
����S�l8<vxC�>�p�N$&nq�5��B|^��U�u�5zLG�ۆ W �X�^I#�{ �gv,�����5]-J2I�T��*�$�kJi�s����-��X40Ir�~�����5�G����g��:��dCT*�c]��Т�\�AF%$������3j_G�آ%�9��m�pp]�҉��~��"n�0��2�<���L�T�a�5�Mį���[z����2c�o�B��M�c���-�Ki���,�݃���j��+	�x ��x�Sx�8��۾�3o���� ��`Hi/���u�yv5̒��{0����M������`q�\?H��f�0��R�/��	����{CG�<�`Qg`o�!�'�T �BV�c�^�nO5�a����Y�ی�U���?�l#�`��'I(�E���lK�N�u��Z���e�*��6��]�Ќ Ꚓ�s�j:�n{�>���+׮LC�?jy����nH��.�گ-���ٍ���3KH�F�G�"	�.� ]A�+����i�X�`��!D�;4|u��	�)��[��<ee��7�-���*����	H���M��xJ�m9#^��/[~�� ��Ne���f�Hb�CE��n�4��H#�N�I$�����q�zJ�)O�KCoN�V�F�GQ�~�?���p�/`��$i��f^,´Z�<�n����̓}�Y��"��=} +���C�f�Ո?,�~6�O���(;G!&����)Gheoģ� 2�YoA�b�
?���3�5�� �£�K��D<�w�gD 37������(�µ!H=��9V���n�9�]���=���T,�
��8���gd->�)ӥ7��F.��$��@�c�Ӧ �d�[)���k��6 �ʂ�c |
y��w-h���ik<*
Ky �z/���𱩛w�yȺ��vB�:#�$̤�;�T��=Y6vE"5\[t�mn�#��|NJ�V��s�R<m�8�ązQ�sb)�t�L1k���	A#)S@u�廽=�3��ͮ���
7�6�4�Ì~5ݯَkتrx�Lo�=�Cg|y�+������7]:��N�Ȱ*��L5��7Ӷ�/%rB4����ӂ#Z�Ù#�h+��7�i��i�@��l�T"�#��C��	4�]��:�Y��#o�'�uLfn��n�x5J�݇]����\�Y��9Mzy+�"�;oy���$�-��EbPDu���(�S9ׇ�"�b��~���*�G�;��V���bQr�:�}Ƴ爋)��?��־��g
AG%Qz+���oU��IV�D��J&���A������Z��+n��*��!K���"p��"�ց�vU��aS�e7��쮄?`gW�#�N�����z��:���㝔�˛�`)�_�s���lmZƷ�-�6�C�5���x&;�a*yض2{�'6R��f�IL�D�i�̙�I�+]�nr@+�#���_*���lR��cW&�C�w&��7�v��,ߗ]H"#�.�$=����Wھ�ͯ�0�� Q`��Z���P��4�n��x9�:���tD؂^}<��(L�)yq��&���#9�	xy��qL��@W �y�<-7u���CI�8����V���MT�jt�p��hK�hA���:E�0�:�E��sm(Z��V^BP����3<Z�?k�D�4#�V���ކ`@�W���c}}@�G��$LW��I��vM�b�_�Q����\�m2EJ4���L��O{���{��h�`����i�k`QUDj���0�V��[Z!�V�oG³A2a� ������y-����V�NbeH�^��	�|SU�ʫ��O\;.�n�,�2Fj�I��.u�M�,爀T�[������hZ
J��7-�
+�y�9Oٿ��i�M�;k�		`o��C��������� Ӗ�;Wh��#U��S(�/8ܨC�R�xUւ�����Y(��sk̖�=|�������p6�+$I�z��̓>�um�.�F��)�U�.����
�Y��V���K�[t2��y�$���;��5?�'¸ Yw���֝d�ԧ�b�
�f*%
�&�V%��`1H�vIv�Q��?�~g�P�R�w6qIWK����;B��L���XB�D�>��<��#�w���4�ֻ���ebȎ��qang��l&d�731PIld.ݾ�Hp�tD0'� ���R����`Z�Q&���"���u�����2p�H�2�׷5Pg,�_�{P�e$Z�͆�$r ���$q˫�(�i�4cߋ���n�r�L��h�|�5K�� 4�4�X����7S�L�e&'g�b?)�u�	����{�.�Mڳ�����|��h )j�U�҃��}���7�
�L�|p�O��$H/c̾��~䱦���-���`�m|Sо���o���� �'ҝqm�M�����I̡)�����n�w�y����M�t���}p�w\]c|���~�\u�&\k�HQ>��ا�K�}3�S���Jh|� ��7��]E��Su��)׾�f�H'L��:��-x±�����,Ĵ�OG˾�;tj��om����ȧ0��]���T���޴���>�L�J���9��gM}�L�&�6���jqYk<��9�>	ΌV�ŵ����{Ζ��K����v�hN^�#���X�pCY����q���qn��V��3��°��#��v�R���z3�Qu��j?ϭ��q����~�ί���0����!,eIK7"nZ���+���2b�+֘2\"����G�kH ^�!��"���P�ʖ�6��vGc8�r����.�􉚳�g)x#�\���nD�OSY�\�{�9_��e�U$:�[�q�Q��?WV�1�K6���C!:�ћA�o���K�[�����Z�B�U�eق���/��#6����pt���A"�sQ�%v�b�e���?�g�?�hm���>X��������2�zn#�����/����(���B�z1z_���Ft a��������)�D�s���:�����������AJ$9Đ �	XJ��M��cl������af���1z>(?�4SW�!�l k���R�oeM/>l�U�)�֠ Q2���%>���LP��óxCg�pB�t�l��� A���1��`���+�eI#G�{O�m M����J I�	6�<F��;�'](/c`m�]�OWX�C/�ʀ������A3'(If�Dt$G��:�޳��ޘ#Ϭx��3��ܿDh1.؟�xm�)�+4l �����ϛ݋�2��h�$���[��"�C��u|n	/����B��`�"'�DR����|��=�gй���.t4�J�"	�����;,�(�:��xv�V�t"� �� ��#ј{���[��j����jN=�м׳G���]�Ti�'�'��|h��%�z��/g[������&)��E#� �'�=; =�U�qoz�C�!��ءA-z|���b���ٗ"�4y,|�X��f�\��I�a��P��I8a#�H2c6n�e��VY���NdЊx��G��^� ��ɀ�P�ϟ�s��i���M6��&H�ĝ0u�$�;{"��z|:�Sc��@�^�-��a��r��7�'�1U�rͮܶ�o�%_>�Z
��N��*I���6w w�N������� �X�ܥ�暴J�'t=9o��>Q	Bd�E�Mh	���*tyù�A|���]�|���v�1�u���.f�����aǺs��z���x�zu#������%r1�~�Ɉ���L��!��ɞ�'�m�H�g�J]���/���H��Hיּ��8{��v�Msg�Fy(J���/25:�iKҚ����C�Ο6)�|����@�������6ZǙ#�i�\�X����ֹ��-��l�vU�{�M����5W�(��2P|H�&
��Hl�w�`�Y��V O�ߎT��� ��C��� ��Fv�=�N�VU��i�~��F��F�C��������+S��q������}��*I%:�kJ(�|�RU���H��mv�>^���o�4T1��/��_��KM�p�]�ײSR�Wd�e2
�v�˴!���k���%��J�ȳNS$�G�z��2�4�m?�{���Xj�O�]Ig��h.TK��I$g*�۟Ue<4"u��~������F�����jh�7 �����	��6U�4۷�6-3�(��H�أ�S㘼'��Tn41�(����:?ђ�R� �F|���6~	�n;o�	�	1����[<�A�6��|�vT_X�]AM�.�$-�H