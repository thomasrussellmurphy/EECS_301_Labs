��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��V�^�Z��g��*3��7F�>���`D٢�*��k{�fbq���M٧2����R)��fCM���jGZY)�B]�M<�b%Y�>5s�����$j��t�Y67��HC����O��BG��p'(Izȝ��c�?'�ć،�@v%银�!``70��9V��G.�x��d�KcY9�LJ�&y�[ʌF��|I�����I��S���|ф�E���#�(?I��o����6���\x����N�])\2Ke �`A���)B��Q+�C���t��:ޟqo���֛��Y
!4*(���Ќ���ʦKYׂ�'�֍!énYG44¼�3�ش�6`���pՔ���<a�>�a���t^�8�w# ���:�y=f)��8rE�apݿ�Y��y�哛C��Ih�*�z}�Nm��#�b[�:ޜ��/�k߃)�w��C
�n*U�Qg���K.]ɸ4�kU�?��i�.�q��/�Q[�����"w���-Ԙ���1�s���ـF����"R�_؄h+�#��؉
��)n�r�6}�cҧC\�Qy�ls�#g�E�X^q�zT��R4�|�/d3TYկ�Of��-����k��َ�����&tx��������n�TWmV��_��
Ml�ӢIc�c�~[��c����fioZ0C7&AI�LUi�)�S���]�vY�Z����i�����M��`��	���v�GA�<�|	�~�1[���\�!^T���h�J�q~����]�2�B�m��^��
=Q�h:a��Uf2+�T0_Q�[6�ܡq�-�E��Q��e��8 p;p�L��� mv�S�^�`���#��Ow�"��z��c����;���ǂM�����EA�6|D������H��� �]�V�=�
��u��d�DV#(X4f��2+Q(o��MC>�s爿�,D�h%��Xcjl�>y�V���u��1՘��	����(����_�XEC�f��)[v�?o ��[����_��� ��[�]�b�����J�>mh����X�q	,fQ��̞'e�T�Ntdˢ�\~�����y�����k[$��餺I�:�[�j@�a꺳�]��9���;Q��%���a3�_�]�z�~��5�������x��bRf�m>|���;���Q�ȏλѢ�D]E~�u�(�.�=	}�=:�Kr����#���y'd�
X/�O����m^�θ,�.t�*��Y��
\�$;:�ɻO)�f����Yn��=Z�X�oX��le~���,�1�i��xK����p�H�s�$�o�n��+�&�+�*���( �����N� tY�'�S@��g�������q9!k_�x��X��iָ���v��OZ��vav�|� ��S�5���3��V��q���V��D�\��0�~�n�u�؂Sۊ&R��n_����09.��d�Y��>�ZC�x��ߏt6��E���n��ɽ=��Q_	�UGM.\!;�t!�U)PZ����,=w�%�ɏO6+}�pIl�"4s�_Sqb���RoZ��=�����9빎/��:������V
��ū�T���Cg���S��ڣs�i�9���c�$U�:t$8�Jx��%/a��}W>��Ė5��;5���^1�v/��f�h��12��|�Ͻ8���s(ǺFzѤ_dF�(���	%�"��fâ.�RB��D�x�C��j��I�O�Vf���]B#�{u��(A1�ɚ��v��'L�,� ��ioE��d�>_)�&<���dK��Up`M��|$�F24�]o 	`\�|Rӿ˶{������j
�)�	�$b��
�>�+�p9�1P��U�
�2?7[z�P� *�Q�sspV�b����YaI�̋z�Ƶ���(�UP�-9藦��n>�!�m�W���f���c������<�ꐃw��T,�͝c�'�>ӓ��ٷ;�zȦ�^�b���Y���w�Y��.QM�e����t�[ƅ�T��+Eh�ܵE&�5� ��jW�f-�O�Z�L�����eZ��� fE4��qO"�b��a��c�Q��Sp/ ����H������_qehׇ�򗜢<�ڻ�\+����7˴�]f�Q̈́ڿ�B�o`�Z�!P�g��A��t����e5��k\� �3Fi�O�>������m���u8����$h���a�����hǯ�X�l���H�7�Y�J*ԮS�C�}�qU\~�d�3�nӪb���fǹa�a,�2-�kIIި�E�9� Ħ(R�D�T�A��Ů;g܇K��og�u���A@��*��(�G9;�Qy�I�6 �_�4_��4������2��| /`,v������4D5|:
+>�Ɯ��!:��/�=q��m�X����q���#^��-Y+�a��-�̿;���
^���@��/��u�|�pgl��Y%��	���1 ~g���.�X�s���6�l��:�E�2?ɪW-C�K��l����-Oq6��*�i�R��0�
�6��U��c*������Jf�Q��������K
=b�_�إ�u$&v�A�Fah��Ws�+�[I`�G��<��̼ڽ�3���-R�i�b�T��1y3Z�.�G�X����d�@���yas��%@�0c���.��kU� �Z���smR++��H�@����ed���5ApBN��mΨђ|��xϨ��JG��:^&� qi��|sW��OއC|Q��|)R�3+�C*Z)H"P��%�`�*��OkY;`.���B��EvP";O�e�˓�ib=���AE��=���u���N1����#�M,�O��^*��������O�Dҩv]x�>#PL�"T�`���\���2c������x^P0F#�>.p��1 ��C�+��\�e�8h:�3�:e�B�,�c-�6'�Yj� �a��Zm�F����-�=�%t��Wߋo������1�0o�"$o^ ��f��EK����pŅ�XP�|ݍeu�.�	��Bǘ���?1MQ5p���|�N��:d��>�F%�a ��L��7}�'�������K�1���q���Yr^���-L�R^��`��N�f�Y*�2㒴p\f�0I�Վ3��Yn���4��Buȅ��jz����q��ve�ױ"6��_���I@ouN�]>��ɷ��W�]íN����g�j�G��O	��6Y *a�+/@P��	�/����=�R~'����g\Q�db���!�����T�4��~������1�2�7�����C�Bl��%�ׅ92j���?Ӷ�YQ��'���i������N��!��`��^��$���I���L��|v�^�#=��$�F#D�����=c��&�A���E��R�̈�����@��.A&�P���d�uL�]���íkP5Q�ԇt�a	>w|C��XWF�����^j���ǩg���RwV,�,\�Ɋ�@��V?f��Q��>6��[-#� KID<I�6�Z)��zj����F(�V�Ɩ���R�����ʈ�.�Sp:V7�6[�78�s{�,3�R����n�M�Y��wv<�_�Yb�hF3��>����\s�$�Ȩ�X��eE��+E����E�1��!�|�Uq+_�C>!9��I�$���@� ��u���"���.��%i'���8	ٮ�٦�0/)�ThI�b
�.�"?6}���I����X�h��n3��B%� =��G���L����)����v���]�6�Q����v߯��r��G��*��HF&]AHn݇wzZWݨ������!��<+���]*��,�߀�<8�v� \��s�d���~���F��on��4x�ođ�.� ����8�M�b�y19 j9�kk�����\	��}��}���/���TZ��=��W����tK��Z�]L�B�,%LӚ'�q�!bttfE��nl�\����U�B>ɟx�=��Y5`gs�̍{t�j�&;�o2.sؽ|ښ�
ٔ�����,Ef�Z�5L�*��	%aa���Fa3ˍD&���.��5u���0���k%�Y�Ȱ�}��/=��k\�oy��kP+�5�<LI����JTD�B� �8'Q�k�f�0�ax,X���Xϖ��>g��q�H T>~o�?`'YE��qu��\˟�p���vp���=@T�������F�ӭ[M�\�����?UW@I��ȉi����C��>�|�v���8֓�$ư�'G���B����M�:~�/���������<�����S���G-�Y�mT��{vd`��{WR��EA�G�>nZQ�;ړ5!y�6�妀V�"b�Zb�g��p5n{	�be�;2�M.�����7�����T��W�.)�WMR6>�����d4�`}k�;�u;^����~x�uY@v�/���@
<7�YԻ���9��; .���f7	F�ī����}�5�!Ɂ��ڱ�hl�}z���[qy��@k��UCN�y�m�T�y�ߒs��~��ڴ0TB7�7_���mi
�n" U���ms�~éi3,9Z8*�Y�.�V��Dx���&8���`Dښ�h&�A�`�����"1�	\`*3I� �5X��p���<j�#�W�W!=��KT>��T�":��,�l� Z��?ͥӭ2����N	[�(���j暑^������<�<����O�]#穅'� z4�D9��p��u�Yr�9la	k���BU3f��ߙ�/���X���A�؀،�c}�H����ކ�m�Ϯ.Ò ݍ��=�*��m�����=<��0j�0����Z�[Z�$������'Y���u�)rU�܉�m�Jx�Oa����R����P`$�����̕>�A�7�#ŢZ��,]��m� ��In,K���B��܃$��	��G��D�F)��,԰�;Qr�6��n�T�;��}O]1���j��[^�\=q�I���s��o8 +�����jE�
�Zy�MJ�q���eL,��r��;!�zPvͰZ�;�m�r��5�J��"���4!{��*���w�z<���t�/X�������=C�D���_65$#l�W��F��[d�4�Ifb6B �1ftB;��D�˻l�5��<�-7T��Xv�vO��Dvs�%2�[A��<�_f�1������5���t��p@�-�]�s��q����=4����d����>�/��W<	�$C�6��[N�O4 C����X�h;�"`���	u����U.W�GȠ��y�9�dzl�#Ρ�;a?�IډBqBz�"�$�l}p�(���-!���/���cc�sĶ�7��V釸J&�N8X���0�kf����ɺ��^>�r.�/����%)�i�ҵ(�Rʨ���*s��w�0�,���C����!
�3��C�C���A1�U�-^GA
�z0Z��~X�Gc=g�"䰻�\O�p� �lS;�Mg��Z�����_F�d�D���D��E�y;7�̒�4��
-���o�?��,��G3�쿹*'_�â��.��d�r�c�\J�Q�NR�[*lʻJ�2���*�� �G�^o����&�*|�[�3n/�S�i�:��&-��j�h I��2s�4��|+	�!����]O�$�����l�O����&��aTf*�^�4&��}��!Ó/��\�����iM�G��)B�ZĞ����lxV(ܸ�g��[ 4K��Y�t�#ʇW��zO��a眄]0��d�Jp&g�RI�������q�\|7CC��0]~Ղ����r�]#���"in�6fi�9ef��@�ˤ6����_��bJ���/sQv�`^�tȆp�	�8�SQ4��N�l���.� ��FO�RY	���¨�v��yKf:�Np�������z�Ŧ���"��w�"H�������3=���kM�F��Gw�cᘋ2��P�iՈ���spS��y�V0x��B�3�Ӥf����q�W>�vtys�ƌ�ۚ
Gg��aNpI�� �\ρvL�	�Bi5t8�w[ ������Ѫ��x�	�j/��p�w�$��G�b��M=����Um~�{���s��dnD>�wIvL� 9����)2�2��Rı��X���4����������)n�<L��|�I�	����{/<�.ް�G����J��
>�=d�P^�Q<�Ϳ���^�i;Y�U
kNϛ*xm2��TZ�bKJj�g`m����5�-^@�R�YHr�r�^a��|[�J���ݻc�Q������q��I�N���<��������Nފ/�k��H�u�ƕ���L���YتrG8}T`����z�"UHM<.R�Y��_�>�;�"}-H��9e�<� �^�?*vh_j6��NQ���9���9�I�0���uCn�S��o�{��k�3��� r�>X�`��+S�9Dl�Gnb���闬\u}�>г?�54
hvjR��9*͞lf����e_X�2���!�L�h���0���yN�����-�c�� \�9��ܚ[�G�MP�N�*!��<���NIg�O���8�K��e���@k7P�޽���A�û�G�5V�#'O���@~TXj�w��]���~�9��9} �������[+V���r����:�qW���W�?� ��ݮ�4|��ҫ�e��tT���R�f!�@�_�y��s��ʴ�B�%=�&�TY�:±�eN4x���/�U��z�H��Xw��ð�9��]�l��sơ�Y�=L@V����>�m��y��5fE�S�y��Ҷ{`��NzPTZ>s&��Ғ�s�d����U��h�TKP�_��|��9Yk��xX�/��A��L�e������e�):��d�G���f��Р�-�ة��0��[A�s:l�5@����B��̚�x��p���ݡ�é�G�*�c�ޥ*�a��{5�'���A�kd`ޝ�Z�C/�&˕Y�t�նx�!��4�۠J�s	6@��f
@��m��ZA��I���9y�
�x���6�K�g�ܻ�Q���BF8ܻ�=,�,��^���P�r�`��s��_7��C��#�5\���[�������w.�P�r�a<�~�H������ۢY�)|��챖�rh!{7���MKyg��W��Q�ԫ��	rn��`)+$�4�3of4�T����47oT3ȑɁ ���m?޹X���nq�S�@]	�&����w�l�twL��=�\�w�c�N�o���h�h �ϳ��/�X��빽K�>��^Z������)���V��N�ԕ���Ie\�$^����a�>Ը�g�ۉ)��k�J����:Y�D �y����JU��n�����g���͞t��0[��/PMq'/ǧ.$x���SA�A���$F����K����qB�>j;���q^��,���wz�F��x�˰�N{[�K��f�h_-h�N��E�gĬ$�f��0��za���!����g�X@6[�u�_�4��o�X/�di{cMt�w��yL��i[]�iF�G����yy^|�50rS9��9��EX<�2Fh�W��A�ԖN?8a��ٜu/�1�Cs�����A�#+�r�N��?��\J(9R���U�E̖Y~b��C%o��L��hʧٟ���g�8����Ċb�O-x�+g����8�f���@��r��0������oi�