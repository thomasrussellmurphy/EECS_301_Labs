��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\���V�fnvx��ÍG_;�ȅe�~�>���9�>��Y;�0G���O��������Z��J3Q(J�˪�-v{�]���������f�\s��\�>K�Y������2Z��di�������b�5U:|M<�T7K+�J4ry�'>uT�x;�E�K�)�l����;��?��XRј�3J��6f�"<��!L}�'c��	���P.��4��zu�tT R|8�^��;pK��'{J]���,�2���9����10"�%nvG��ؔ��s��I���n��8^\+8�%���ΛrZFm�Z^b����Oy7��YFtP{�ھ㬣�{_U��{��m��F�3g�H���$R�1��Ÿ0�s+�����2����5��7��&�kB�S�3�^�B���#`c=팾��1�"6*����l����d�QMe�v����(>V��qT��Y��4�V �v����|�'�*�Q*��L����P�"Ɗ/��]�Q40AF[:*;�#��>�x0���Rj+=�I����QZ잡Fޢ�Mf��g,3!��T�[�.LN�T�d1%�JP@�~�����#cj�ް�]a�w7�^��~��K�e<��
q�>���s�&ǋϠ�'�8�0b<b�D���ѽd��;�ww����،�8U��e�a�AR=�r�	�7M�,�Yvy��b�;�&��M�a3�Sa*������z���^��_���a��(59D�;?E.A&�t��:/������)M�="��9�|�����(��ܪ8[�<��p��%� ܓ򸒈)�ǃoU%䝟�#���"O����Ξ+�����ܐL�z}q�Uy0�yPU7d�#���\a�kh*}y�LFL�|O�I��ɫ �,)�#yuiP7`�m5��r~���c��/�q���=��uC�R�~�-y�i���$R57׫N���$G�Vi�\�{<`��Z�	�4�/�p�wzfd0����q�v�بd���W׻b�9$=�&�!�n`���XA�O���� ��PRR�m�6�@)Ug	��r �6� �.8�|�;-�{_ʥ͆�.�/%��U`�k���>�)T�c�%Vz���7�tG6�C>R�ކ�ha���Ŝ�>A��wH�S��͍v����������a\/�������^I��SD{2���?�F
Wa��*��/5��U�B �X�S���
uE���TT�4��X�����I9�  ��|�y��Zg!i�+F�s�� �_e2u�k��=�n�E}�$�MX��[?J1��N9Ѝg*�#9��`k�߸�"��=�­��i���p���eM�q�W��6kH~=�'$�
��2�	��D�8��U��'\6rm-�����B]���T���K5���CñuƷ����+۩�>��ZP.�6Ͱ�Ā�5�yU�|i��o ��p�U�[�@�
%�(���U�$C��B�a@2�+x`�i�i�y7�@eֻZ�m�b�m���Ik�IA}�	�p�NG�[˅�)kO�>��h���}�i� ��^����"�YⰃUX��&�Uϛn��ۗ�Yv��X��0��ff�7.'eЍ�|��eF���E�i�[��|زމ�w3��ǽ�q�>��!�:�A�R�X�ꉁdЈ������D\�8IlM͂�y�hIQ?����Pa�܄6������=MU�Ii�,��-Q���>�ii�Xf�>�5ݳE�\�cQ�R��(M�Uƥ]�-��`��C_"�t�b��4�A7U�ኖT��p�xӇ��������+T틏��-oo�XD�!^p�7�X�(/ˍȟ����va���6�J_I
7LI�����C�~+g������.��Z���"��Hê��3� �źW�L���f�O�ފ�Bm�:ToA�tuT:�i�$#�ہK#,Z:�䖩
5��0=�D�����h��R��F����X����m�����K\e�t�:�N��Zɝ�#�79��+�6�٬+�-i���P��$�|s
A��4`�ܞL"z�^���7��V:i����s%˼QB��*A&;K�#;٤LA�>�m��O�� ����< �T�AD�Bn~�]�N/?�c���G���7pf�W\șk@�_���.�7����-��eW]�f����G�F2��͈�C�g�z�c\���8�#�Xp�&z��{;�B8_��>��;�Xx�'�ʟ�r��`��������qH}z5/��Dխ�Ize��e��5�����ZR�( |�q�[u�sZz�u9�b��v;��V�sY`)�R֘L��/�E�v����V��c�+# �bke���W�p5��©�3�1��P2COd�M���]�`bҷ-J���*���R��հ�#�.���OH��#����O�&�`�F��d	��AP� �"Q���&B�^�@�f�̂��l2f����7�ޫ��eHu�U/���H��e�4���a褫(	��Il�۽��؁yW�j1<<����8�O�]�[�^aŝ�$��@��X�sX� 1!�@�Ʌ[ �́���`��@5�I7��������Ç&�^�J#t�`�gP
�K|&�,[F`ȣx���Q�"�P�%s�J[���<1g����-/$@�}�v(��e����3 �zI��pג�F�"�8���G㙔�A%S�:Orlvn�e2q�G���щC8o�Eky?
R g��hyg�U{ m�]��.|��ݽ��M�uw̐eb�8�M���\�����1���Wy�$�A�Lnx��{(�-����$�N�jM�[B{�:��f�Zp۽����z ����%svkѓ����/M��{?���g(��M���L��̃[i[�;Y�z�Z�v0Te+����ف��"7\������g��n�.yst�:�+�R� ��&�����p_ɰ�@^>�"������k��A��VV�����	���P#Q x�����Ȁ��$�d��<��'�	��6�&%^�.�a\?G��t+|C���u��FXG�L�O��ݳ���ΡD�9�E��H����O�]�*����.�&'��ݲ�i���m1��V�4�A7�g�ɂ�� �(�;�x��0�έk��1�xzc�
��1R~��S��S?2Y��Gʲ������nUagգy'��A�E�ﵜ���F���}�S~\E���'����c����� �g��M\����B{b6K�&��S�A�M����]!Nf�7[�CA�cJ��rNCv(�ܑj02D׆`��єH��s���!���`� � ����{oI��S�a?��ZL%��O�7�LO5��oY��:�-�;��"ip�i2��\�n��
O�F�C��i��@&���z�u�:#A?}�<��������R��JXo
���|5-��u�C��֩��3�Ͳ�f��-D�����/����[�W�~�Tb����z^���m��Tj{������c����� �6��\�E�ӝ�!�8F�z���;Z���k��t��Z��Z����<�=���&���������=�����9�z����L�O�]����wz&�� ���L���� <krxKa;g�Z!T���t�3O����ƙxV�(����	��r�dI��v�?J��	��
���6�I��=ڎ"M�jŅj���Q׭�(�(؂Mr^��.	�� /�_���2kB��l�`7V�,6ԑ3M^��T��������3�*D��{���8*��=��2D3�(��M�
�������z����ʖ�����eh���w�X��V3��#�����bHd3GPG_�����{Ή{kx�"�l�YQ�#vs����!
�adI�<��c+�#��b*�^���K��z "�YTS���eX�H`e��:^ ��s݉D�ӂ���~�^8\v��u�#��(���w���/����7��/B֡3�%�wIF��5�(.
�%�I3��p��~��|�HKA�XT*�RU`}�x�|vB�a��œ���`?��G:8AZH4^C�-Oz(�b�:H��"]"#t?���C�7V!nV�:@p�	A�f.B�S2�E��EW��j��S�!�g��s�F`I�wxU���n�f�\�"ZuA�\�"��4A\u<+��cθ��ū���V]�"��r���31���#w�������0��xr���h�ᙱݗ��(�e0�f����PW*�E���f8�#��<��+
#�<�;�����	����p��_ٝ�-�iy��e�SH"g8�B���&<�n�n�f�I�3]��ޖ���2s[��t��j�;nl�cI���
�!s��:tC�VY����E��/a��\E�&�/��7gw?�e�r�9�-���d��4����b,�QҜ�܀r��j��m����3��@9�)Ko�\u,����N���opV2�P��c5u���sw�0C�Ċ
��UA��>���d�\9DDZ��t���Qb<BEl�X:@��E��a���n�[*��D�����Lb�탬�$�h��N�H�7��]���H�����T���}*�����~�t�Tۑ(.�"���Mr0��G���d!�|�h�s�K�L^ɩ�Y`[�/P�|﫯gz��x�S3���{wm�S���T�x=5tB�7�y���
��V�s����pV��YX�
�l������H��@B���lGU��DN���GG�x����J:�-t$о�u~�1N��Zl��W7T<�y0v,�e��h!{P?�ĩ�c�iIG'Z(2�'�O �o����v��rs*qK�>�0׼�kJ��b�X�H)����&�<=�LΚ��O	�B;�"������1��2N�� /��@���`-�#nlwgS~�r�#�+���I����ط�^d�6�t���zPR6*P
2p3Ϫ�KU�H�Epc(O��ɜ9�g�����cx�<���8 ��Mi������םH�00>:y�h�~+�\�jR�	Ѽ�.'y�c�h�3�̭�nK���7���<�)s���-��T1j����v���)�E�V˸��b� t]�uS{����+Pp��%n�g{+U3�*��ה���ax�����p	wS�v*�)�_�yT�����>��{�"����C�Q����7�N���"�'*�N;��x�g��2Th�̜�}�F���C`�iZ��m��/4� ��p�i�������Zp���B�����y�u�֯���b�p8��*��r�t������s1�?%-Z��$q۞ߟ42'J���R��\*��GիґӒ�9x�K��zt��P�Ú�:���L@J0��627��n����\3:f���S<�%�G�{�(�w��ݎ��L�xZ�۬b�}ݴD��|��Avt�:��|�|[mCN�"�~�<���+@Ϲ�$����X��n>�*�K���~�h	��\�^�_�afu\cB��Jz5�3�?�(�?�[TiN6�#4�Wd���ىS��45��q��":�ӭ�b�P�����-�����i�,�N�p�zh���NŃlZ���;l�L#�������_��p[��r�!��w7�o�HqT�����S��,F��!%u	'��F>�J�Ȱz�Xx�;��.��lT s�t�M`*�Z���q��?q�|�g�v��p����*+릹��.!�Y9&��ޖs�k�D�#�2γ;;���������|�_�bV5M��6�>�k2�v/xh�cB������i/X��N��S�BƖu�?�\1�K!-�v�uI���3FQ,&���{�tG,�;�d��Է'\Y~F?L�N��Y)s�4��E��2�5m芆2g�]n��H�_�?o =�ͣ,Ӂxկ�g\�T�}� �8�� 0^ت����	�D��rP�LM�E볓�@<yKI-l���r�S�耶b���Fh��xY-�h ����; h ]9�=<U�>�$��GF�Y����U�c#�d�_�8�{2��ܬl���%(�;��<�T�����컧V�[	թo��Y�ic�u�#�?�W|�y[����c3�9�o���f�w�<O�)uP� n�vF���@y�U�>+�j����;�ѺD,�K!"b�}T^v�ڐS�p�3�����z�Zw�C�+2\�I��:vз�?w��(�B�o�_�·#�t�f��	`Kĺ���1��%	?����&���1Y)ф��.�CȐ=ǟ��]���$_�T�+o� c��m{�:ER|�RU��O�!պ�*��ެ���U��������;����M�2�p8t���w3����y_l�tv8��)�`��i��{1��u���#k��CY����a�EK�?z�;k��6��J�P���{���$�3&����`���0��'E��Z�9�����1+���K��#��#@3$�i�0� ��`�<���D�"�-�.5:@����# ��^%"o!|P��(c�R���u��'�ډk>��د��N��R�l��!��k��� ���w4VG?�A�pBT�3%J�tz5
54�G�����s�0C���X.�5V/S����ъrmȶC� �?y
�e�X�rm.k�N����f�I�.%L��<�Sԑ5*O?{k��>�TI�Wi�Ǯ��);=A������7'�yt{ʲRM6����C�8'����*��Cȭ���T=�sAH�U�@�Д�2��u�|GX^j�(�|��x�=��+VS�'��S���Ő�*.5��ff�ϯvm�aO[˗%�h�Y�O9�7R��ֲ�9�j�Ԫd'�!�!���@�9�Z� �y�썻�&�H�R"���s�Q�(�P/7�{(.���K�4Ik���-�L����ej��[���}��5����͚z�CI%�v�I�p��V��\/J3�@=�LCm'|V(���CL��t+��)@ː�o�'�P��[�(|wdb��f?/Cl5��|�Ƭ��~]�7Kw%ެ���(��ck�&�R�@-%uA	#�'gL�b��v����\.0ñM��A�znQQ$��|�omq�q[R�w�q�a�B���\�q*�؀���Kh�#��s"��N���鋅"���Z�8���=/y��	��h"�� ��,�{�����&m��m����-��CsA[ H���v�&�p� ���[S;�c?����r�K�+8�Lp1%Q�y+�%�V���E��{��Xߛ'��{��5��)]��sB4
3�q��9������9$�e(�J�Ė�_
�1�W�\��a�}�l۽��տJT�4ם��͈s[W��}���s!ce�A��:S.qPZ�y��T�\,�$n`!��C�m�bf&N/���｢���Ԭpta"�A�����L��� ���b8��lX榋��ЁD�L��m"I5�CE>mm�����^��a̴ς�;*�!s�Ĳ��ߨ�)��ʡ;����퍚XI�S�ȼ�z�ñ��.�ZB݇^�����ѓ@~ځ��U&�=R@����	~[�նY���.uB ����2�bci�Ӯ?�nA@^EpG-��I)Qx�Ŵ6!7+$�1�q	g$�`���p ��l!(�@����34bؒ�a_�]a�آ��IF��sJ�Ox��Ԛ$s}UY�*K<�2lPo��R	'c[���x;9�Yƨ��8Q�������� �����9b����B���[�:G;qv'&F݁���� ����`�5��E��Oz�̊)��+���^�z���]��9�f(=�s���m��6
���5��0q�(���B>���U�9��ಖ���+��֠��l�)-|Ó���L�խ|J!8-ʛO�ݦ��fIT�>6��7���
����GCj�B�kዖ��V�_"*5/i�b��!�bVׂH�OKL�^=,�.x��!�W�;�d�@�����`>���^v����#uۇj��s&`s��'�=p��Z��=��~y)���Vu�u���S����J�A��Y�W��Y�� 4�����8 5���U�#��{x��uv�v�U������Oe���$4��|�E�ՐI+l}�Ȩ{�?��]gv̐����E��y�[v�`[��p�dh�e /��V�z�n�l�p�W�@�	������mU�C��yOY�a�k��F6ճ�p��H��� ��##}�O�Gp��w�V`�|�1�$~��~Ks�����$d�畷�t���fjp��)�������~]�[�iݲ'h�H���j�=���YJL���ӈ(�y�:f�p	YP�+N�8���6�i���ܘ"-�����獙��o� W0�¦S��[�J�������d+
V�m�ڵ 	!~
#��l�=i\t�}9QP�6)| �I���r�i��1XW/Z��y����Mc�\�2�d�������5SՀ�;O>����}�8��^���xm���IЎ����c��TnT'f�3~p���v5�2	9ڜ��\&9���W����zi��P�>�w�L�������J�A��3C�o:���!H�l�LO����yTR5!P�Sεn1a=���y�S2K���@A,�KF}E��_����̎`��J�5Gç?����vVY����-���4�E�8�*������ѩ��ߵ��f)��mFU�Į���3B>q���~�9�Y�S%_��G��.�(��ޗ�u���0�C���(�x�H���bw���~���L�+
�:�Ěϊ��Cgk��A�m:;��H��X��f[l�ę�-WK4?f��Q��eF����yƧCG����k!�X���������2�\8�`p��\#9>�#F��!��
 f�}��F:�6%FHP�R����lyb[���ɿ?k�rw��T�o�C��4pu��ЃI��������X�]�,���dGj�:�v&J������X�4�C�_�I�̍�M��6���~Oc
��ŻH��F�q1lgi�g�mñ���
�B[�޼ݸ%'뫉H��d���A�	2G�������X�)�r�[(�Yx�|I6�'��h'.p�p-J�պ���{"A�$��ҷR�G8�{1�7.Y�`I��d�ָ���+�n���%�%O�;5��ٲ��[��Z[~�U	�\��,��X���
s�e�:��s�h"<#؊?8������S��_ݶ�E�;G��o[��֨����'�ҞN��#{]��5�jO)V�����H��+�̽�md�¯�gVd��U�"R��`��F����wA�+�<O��.W����qg	�T�DzۋEH�ʳ�bD�	�y�H�5�Mf|d|}D�nJ��?��űT���ƀ��(�q˒��>�������#�ւ�ů����s�aVVd�e�p,gMї���Ȳ�%ٝ�K����7��q���z�wNQ2�y�����[n�}��f���>����>v�/�J���p�B/8���a�(�~��Y�yL�@;h?7�`��a��ʼux�"�`��A�!9�X~����տ�׾Y��*��%�HB�	7�t��T�Rd�P�E���m���t��޵�Xz��zi��ue8z���/�i<#<��o`� l�p)Uʠ+\6$=�5|ݷ�d�Cr�\X}��[�mM"R0w���L-T5�d8����@����T4�C��co*�����dS���3>�d��%�U_���������B	�E�t�VTF�J���	��-������7�/R�0��_*��q�Ѱ���KÂ?&��ȒQy����/�
��^�a���j��a �x��0����s�61�Jj�������:6����!����V~�x^���ey)�O�Pc#��j�͢�T� �ժ�\��Y���M��P���tD�ަk4-�m����ޭ�h�"Ǫ����h�慢�4��>s������<�)t�+J�] �?4?Q�#Ӟ�a��WlgpB��J�+��������Щ��r}��~�u����ϗ�D"��ٲ�(���8^y�C�03�E�v0�^Oc~F�6"�C��lq6D�C�����w�4H���w<ݥi�܃^�M�v�<P�⫩�Ÿp�yd������sL�U?m�l��k� ��#x?�P�j��
���SBTT7r�;��y,��]�.�5a�A/�����3��]���|v���V6q�0G�!	^(c�㊶egʛ�o"��s�r3�]q/�'�mҡ���U������+��)�`��5]�v��`>D���O�
�*h�'4�ZF��2{1k�"L.�A����JH��]6W3�ӌ~Oq�:���M��p����Ta-& ��ȹ(���th�U��_܆�-�4��g*G7;�-�v�c�R��H�@;��J��Õ<��=��ΤU�N�N�V����d���W�a&������5�z:���}B���*�:�xȦ,�7L���$-ϧ&�Aͼ"����{��&Oߟ�)D�h�q_~��|�e����I�͘��pŊ�]��-��fYW���@���1n���I��#�Aɸ�!zB&C�Ә;!^rRr$���c�nP�"���ckhy��i��7����#��w�P3X���k�8130�'S����*�g����ɭ6�^��jCe
h��mB|�4l��~��:G']ֽ���g���G!�{0���O/�����A�?�k#V8��B"N/o��c-&�Cv�/�#XxEg�`�&���f�Zq{l��R��h�2ܫ�t��^�0�V̺���QQ�O���E��MIeΤ��i��?͢�L!B��5�0#ړ�O�9��o�/O�P�&�I�]�& "���me3��0�<�P��Q�)��;�{Oa�ּ�KWLz�����Z�|��xQ����*DM#�V�8bd��{i~��.���2z�i@��Eqh{��T$Z|�"5{��꼘�g2n�@��-1��j���zf��P��}y���{��r��Wѕ�.l�OD�,mN�<�E�Q7�~jp$H�=�O�gǲd])!8�б���)Q�����VT�ȣ�'>!'��1l�}�Y3\c���x��FM�I�f`'C�`�8m�Q�� L�hx����y8o�ir���G-���o�#�҂�6hxf5I�5*���}
BAf���r�� �L*�����8����}��:�Y4,·�)Z���9}�KC3@rdj���s��)�j�=�?�dJ�P�Y���}���^�ک���fg<iH�?��FbB>��j�z�s/,���5�{�p�ҥn��^�d��|/��Κ�_ǜ��ܭu�ظ��~Y;�ZsM��O�#��MC��>��G!DA����ɡR�1U�A�[
甍9۲w�S�݌IG��X�3)ެ�]Z��T����u(�6BGrh(J�dv����=zI+)������s����z~�5j/��/�s���Ap��>��֤��VBr��x/�Z#��oT��u#� >�����&<h(T���G�\�;�p&��/	uoO:�v3�]�U�BPQ�t5n�����
��V�H���l �Y�Cꜘi^��a��:�ߵ�sz.���yC�(#��0�G;�z��ۓ��ђ�$�G��s�+�$����w��M�_w�0���V�j�&�ϝc�P�����q�M�)��}��\��Q�N��`OEM$O�7Uw������μm+-�5��G�b�a����,J����T_�.E������0d���@�E"���ױЀ��E�o�09����Й�5x�p����U!h|!�H���v�,�3��CC�^3k�( ���2�ա|��: ˶R�|�
i���[������T���)���xR9l��B��BG�U�O���3�1!G��~�@��STz��OO�3��N�`_�P�΁-W��d�f&�2@�V2��Cd�d���Eys7eC�iФ �Ѯm��#�7q�TD�-�vv<0�GzR�� ���_�hqZ(F�����ݓ���$X3Q��?�����I��Z��.�c��k�A� ���bLEL_���p�ƈ�xj�ζ�}hSD=i$vP7 ��������ex�2�/�]� �b��AAaҞ�"��n�>�I���l�?U�8e�17��ίl��2ªn?!�h"t�Ϻ>���W�x�,`��ű3��*�~�:�Yt�{�SS�3��Uߺv���x��3K���6�u��z��<4 ad���荽f��;_�!��|�Ds��m5��p┃��&� q �n|m����� ��PmX�d�PiMш�p��i%���U�i�R90\��Q@3p}���l�=�B��h)X�qd�
K��P���鋏R3/�w��v��L!�� @*�:<��⼮�>MPY��/�F��{�P ��Xu�θ������U.���/\C�M��{�x�u	c6��4�
S����&�<���blS�˽��s
/��2�P�G�S%C���`�����r7]�$(�N�H�N��4mѶ�c���`�VT�,6��^�@ A��:�{������rr���ǨM�Z���D�w�/'�I�/		�.&�؟�9�;�+����f�}� t��3K8����Dduz?���
����|~�H�#�����$?�^���\+�W~�� 1���F��<F��ǙpV�.��0QE��Ӭrw}[���Hz+��
�;�c�V�[���Ƥ8-o^��PP[?WtO�Lk��|��$�H��֌�-	ݎ{)�!����3�����I��b�?��ףq]��`f�(�f����*���i�հp�q,Qwz&���:�:-��ө3���^�+���̑��Nvu�.�_j��}