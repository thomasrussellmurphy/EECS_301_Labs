��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>,M�Kߤ�I�;�b���}W �XVH{P�p���Mǚet�ڎ8��iZ�g[1�� �	�ݩ?{���%����������
��y��b��@�3'�^w�YW�f��ElLJ9���{�Nэ�B�����&hb��]0[NY�%�.���r +9�ؤ�+,���
�_"*�)>yg���(�>f�Q�`��P�$@�����h&=�R��X�&�}�:�7y:x�F���n��n+I����ps�QL9������#��N.qw�&�� cѧ���VF���s4t�HOĬ���.�a��c�ó�OWz��;����xD�Gcv��U�D��<[���,�	�=0־1�Q�t���}���EN2j���a,i����=�4��(�p+��̕��Ń��%g ����h�b-wnh��B��B>�% G�z�u'�8�w��v�N��/�Ʃ��3��u���"
��*�m��F�t����g�`w��:i=[톚������2,W�Caa�̌�Lh��'�TΔ���'n���mr��9%���	���e;1۷�l3��7xs����Y\ ��$@h/�E��?[��0���ˋ�R/��������<�C;����V$�e�~��E05�0�8i�;���ɝ�����Ʒ}�9�n.��2�"�C<8���^D�����<�'�M�L����CݽZ����X�:��7EC�Br+1���_�n��t�P]����~7 o^������-��*�9H�6�,ٖ�mj��b�9L6�j@''p��Ƕ�U�ͬ<��1񅐥�Ѕ��)��m.Њ�$��y	�p�M�8kd���Hs�@'Vw[љ�/Py�J�#T�K �)�ɺ���GHf�:���x2��cwC�
���Q�Ƣ�)q�9M��Mʒ������z��r�[�ޜ\�-�o��;v�h`�&]kI��?
���P��) ��Ӵa�6�v/�-;��B����w��u��++d���n�q�������dq西�����w����e͸y~�f�����H���HkȈ�~�;���i��i(�� �9b�~˵k0��訴Ա��͟3�8�,kR�ݒ���㋰�3^��Ԏ��m3{�;;��]� ���?�'���8=y4k��H#ȅ#K��	�,V�d��Fy�n�z��x���'x�hS-���W�y�ڴ���a����A�kh�8O(�k3
��f+/��j�L�%�'��u�gL�W���p��ØJ��y�h�
�U�A���֋�8 /9X��	#z|{䱉rx���@�X����G�,��$C�5��RR0߳a�vi�=�Sb
SeL���s�0��[���,�t�2�s�(��FL��A<��r0N����s(�U:gmt)�B�9�A��/��P~u���?��^&j�Y�@J�
{�^��Z���p�m�Ju����~�u9�a�0Vy�:����@R����K����j�]*��l��gq�	\��L��F�v���i������o�#�ੌ�X�|}��(;�m�'F��p���^
�s�K��1�̮��#z��#�yh X�<ѣ�ch_"�󬘧���Mh��[���d�K59�U��w��m��������0T	J��智����Ȍ����;m��?�B�{0�n���y�+,�y��o/��{�~�#�p��TW��˨n��4H�p�m�wf����b����K�3���	��IU>��܄Ǵ��w��-NcI|)��K�s��!��-(�{_�C���r>F���mX�IZ�0�ޗ3x��T���*�m0���^���H���O��P�_�N�y�rR��
޶F��L��Ǳ��ە�@K�TY�:m�]�>1RM�d����.ƌ9,=}�Z�x_�#D��ރ���������ǲ�:�By�ݖ~�ɪZ�N����]� �Ffҷ�K�h6�I�vàe�%ʭ1f4�x�2�o�-�`v*�U����a��ezn#�+�+�Ґ=8L��r���q#g�����g1���Ø�7���:C?S����&X�=>I�����12�킌��4�F��I?���N� Ҳ����+\��@�j����?�%�F7|\�����F�����6��"���P�k���|ƻ�"�y?����g��鴳�)� �^6BC��i�W��=�vl��b4�k�_�)^�HJ�lc�x���E��sI!�'�w�4�r>���m߯sN�Ii;jY�e}�������rľP��(M6L	�<)�u|�>�F�n�
��HH�-��o<�z�*�ih�l{푬 O�U �m�� � 5��Oje@����+�H��\�<��	B��"A�qsE�k�aR��x~i:��Y�g�j�����H�=-#�~(a0��y"�����9��v��keM�����P�K~���y��u�gh�Q��L;��An�,\#�K��R+#$ᳺ-��(�B������/{$8���gFh�{Jhz
�V�� ��jF�˟���ʹƒ%/���b/��"����q)|����+���Po��Wt:u3��H�0���O��zpT�8�&����w
�qM_$Q� ��ߍ�x��r���kQ��N�g�� ᔨ��*]Vta��	cC9�/���d6E@�^�\d\I�� ��k�I��P)�t�7�Sg��Yf�KeO�k1�*�½[�aQ�F�j/�d&�5]\vKpFf�a@��	�@"C������R�S���n���� Y�~�B�*��M�;c�q;|�"��
����,c�#&|.Փ�1�՟�$�<3�B���ž�s2b�{���&	����H�*��Z���	��N���')��-��b�����5<-���>��r�˳(̏�a>+,zP���e��R��'�T/����X~c^#p���&�^�.MV�FXD�Q@�E_� Zi�n�J>�-)`cf����x��w�@ryێx
�S���)�:�,f���u�c���3{�nQM���J�I������G��o����P�W�_����h����ݽ_���y��H>�UǕf�$��᨟S��WX\��JF����$�0G�B-�~��SKc��F��+��V��y�m�52z�Qe�=��l�_<�2��HG%פ�i�w��S�1���w�q�����G��o+��垱2�p����q�)�5h�G�������)	����1�ŅV����G�e��_l{[��|d9�6)4cN������_rˡ��2�eb9�o6�_Q�\K��c�yR�-y��-4����㏓�L~����r��;�z����g}��[���bI�v��!B1%��r�19���줜�#C�H)N����p.�n�@��pr�)�p��m��T��	�d�aG�Gc��J��|����O�y������&}ʋ���s`y�LM���v_F���tg[��#]�+�hԴ�o��w�d)�CG��rЀl�7'����/���ʮ3h�D��q���fE8M}�P�^_kgm�c�W|o�~�n�=jp��6k��O�5zҩ{@��xG..5*C3�6S�5<4���C��]>Ʌ[}�B:��4h�+��Sr!9�G���j�n�z@B۞qBTUp���ĩ�,)~Y������c؃o��! T_�;ؠWZ�(9h�N�՚Va�G��x���%P�a'������11��d�h|a��e÷���K4���2F�e_�`�Dאn�̈U��}�P�_Dj�����4k�l�
H:�b�_#ހ��02Z�����P�>�[�)e];�����{yJ��jG^�$��Hg|��N��g��p@dĴj�Y��+c�;�8	v�y�+*�}0i�kB��xE���B����:be����d�j���/������X��ܢ��X��,P���r����х�z���0r/W��V�N�p��V��+bt��Ǌ�=����U����a�\����L�k*�%_����Ф�4c��{���yk�c��1fF_�NJK̆T�����
��J>�3O]vk�*�4����J������̏�P�3��1=��c�<��)�`tʒ�!";NbVMP�Y�`;�̺R��|%�گ��KUh,�N�Tąz���åv�f��u�ذ���Y����K|7&����������� n��O���	
�a}��t-;R"~���x��i�/����ME�>�%J��@���fy=�cj���ۏ�i�PR~�D2U���E���!��3w#�pa:�p��`3��j�FZ��X�Um�<5��F��ʞA.,u{ö-]�N1<��2�V�}��|�W_1T&�H88����4[tN,��=H�|G�6�!���S�!N�}V�K�� �)`�/L����E/i��˾W%;��ڠ���m�i�#L'h������9�>�W4�1���c]���2z`��>4@�� ��p���f��31�������
0U�i x��SX��jO
�݃�?�z[#�*G v�G��`�W}yMpj��|���ù�q	��eec|C�UYi�F&��`�	�w4*��qZ��s'�B�>;B�ad0���+�YOjMu�:��}�^_s�(ё�^�;�k~�ca���Rj�U-CA��uAo:%G��Z�nл:�9���/����Z~|&,������0��L�O�ܫ�W�k� ߪq�G�AQ P�Dc�W89P��f���;�%�/o�Ȼ|L��;%ɀ�DG-IS�C!��+�cZ=�5ԅ�-�b��2��GVg9o<Uj�9i�'*%���QNt�]M|9W��xJ�y������|,���Œk��Eq7�G�I��H�(ש~�ؽnW�� �a�4��O5�8�Մ�'����,�R���[?�@�1`�9�~N`�/�1�Hu�4O�E&xᗮ`���dz�����s0��#P,W�@]���γ)8��K/y�z0��qZ>�Ϋ�:��t���g��x��Q�7�+��mO�E并/'�zt��F��.U`�S.ՙN�3?R��]�YW��v>L=�LJ� ��é�>�W��gW��oP��������/]{?9���v?4{8
�-_&�m�(����F�?�o8ߝQ�:U.>Sg���D�A�bw\���YX�"E��.:����\�U�w�`�S�B[,�'�U�79v�XpӼ4I)Q������&�4۽��܆}�SUɕV7���F�$1>^�k���
��i
Bc��)��C��*�	�ΆN���ы6)k��Y��#�3sA�eA�:����T:!y���*E��VL���^���
uAt�AX��}��I/f�4\�<���2nX� �qv�7�h"�A7���.�����ko�fw�<�$��y�}+5m����	w�Jq�9�����d+�r���ͭFP�y.;���[p	,5��Zb߶����`�c0��Vt��X^�,���2���'��y���h��:X@C��)`�i�5��<�[�0�`1��d`m�;����xS4M]+�A�E��>����^�<-��I	%���2�È?���f�r]x�2Wn�^�<AZCC-�LQBW�|2�Kf���oAh�I�;L���Pn5���!�h0A>?���� KW���%7]�>�[������@�B0_�ʷɦ��⮯,�E��T���S>i�����_DV�����hP���$���$}���h7~�ZLQ�
'��n�і�T�:�+dI����Ԍo��ϥG�2� ��R�f��}��ț�{j
�4*^�N� ����(×���v/B�e"�'�YܕC:)ԣ��{����=���"�~�9Y�57@#�c��:^j(Z;ύt��q��Ffl���Ì��#���(q�X9�'"���MJač����#$����^n�VČ�*F�*F��i��3/����鶪ߢ���+w�3�����u�N�}g��'��1b9	ؾ�-r�;�\��]��_ԤΡ��I���΋�q,�]���RC����rߩT�X���N5��h�Y�	�jM�#�����_�0��߻ra)cV���恖��ķ�t����)s]sYm~�*(�Cۢ�t�`[��zir̙phq��v�@����1���	�_ʖ���az�i��SP����>S���Ş��1K����w��y+��l|x�{e��m���J��2}����c���"v%��K,�+��ޟm�tJ9�ӥ悚�8�*����픁�=��pZ�Ɲ��E��x�X������{�}ztk���q�Gi攙�Tk��q��A����G�V����U[9�6�|�jw�>�D$e����Bz�w�E�2�
��J�冪V�v׿�@�%gz�o_�n�?Ev���/F�%^�,�#%L�YCn�������[�2K�䶲�<�}���ي1��z�/$0������Ƥ�3߼?���3Ge�[�����v'ӌ��tR~Zw8�,T['�~zj-�w����=KV�Azן��.�p�	D�WF�������V�oݪ�`1��R9�FK���9���	\@܅��]�sYh�0}���\��0X�r��!�_q<�`�m`���/��g��zk�����!�;N�
a� Ɛ�}����){���<8
�(�ũ���s�5Þ�J�o��Фoˢ��lcp�eL��o�6���݀�]/93=���B�6�	�*R�BQ���%I�q��G-x��(�>U���� �2��F��~7���D �&h��7�9��<?��_˯G�^u<�M�ߐ�#F�Bt�i~��,� ��ʹ�].5튺�e�o�4(Ϩㄶ`��Zӱ�\O��1�!�7�-�vL��D}���ˈO�܊��A���*56���,�-6��������;<�cO�C�j���hB��
z�����U:�?����5ǯ� ��i��ÿ�ß��SP������>e�_�T%�_��_E�Q�1Z����z�cx 
_gH�j���T-B_c���=�FtpA��t0I����E>'x��|�*�����ݥ����"-��e�����]g��j6�}_��H,�d���,[��!�@(^�eM�7q��XA���I��\pڐ�6����d*�1�wbYm����j��n�"�Ȟ�;���A��!�f2��6��}��.,��D>�����E�"��P���\�f�#�Rܿ���u+�0V@����ճA Z�b4���h�>�ir���j��>.��pު�����<P�ě�%Ξlͺ�cc��{�c|H��9�!�a7<�y���@!]�嵹bY�X�<f����7����j9�q�#0� �A�m��Ed����aW]̾<�����?� ��̂J�#R2LҘ��٭��u�M���іƦ�5��"���6.��(꠾5,�f#��@)l��N��Z���\��Z@W�X=Te�/@{+�#�.�/�㒣O�S��12 ��v�����ƾ�Y�AF�ӑ��ͽ?������4*?�������L��Z�]A�&�E�������}�*ۘ�����X�Q��ܒ13�lڐR���N�<��@҉f�m��w��?t�<�9(��e�%�$r���?� �:��XB�%ּf���W(ꡎbv-Z���_twե�a-�d�;�|�K�C��t���+t�I�r�e��3�����|�<3��u�B�j��RhYB�\��Yy� �YA�9L!5al.������L^1��|���5u�=�{��o����Q�	�'_k.��es�J���͉�aq�Uf�c�j���c�k ��)	��.���BڝG��4ə�t��nq]�1� ���9�S� sB� æC+�vU����`��/��k̴(���B�y�L(���a��nγ�g�$%1��RM��0mc���omX���8�"v��]V�B#�{�\:�|OMN��n;-�i����/9��ԟ���3�^��H/���{��Y�`���?�	|U\S��n��z5����6��N���l��ð����=x�<+Uבv63�fA4�1�:JS �Q9=]㫬�$��d9�WS̏qd�����0����Qyĸ�/ʨ\��S:��y7�u_`|Ͼ�4�-_O�_f�p� o�du�:r��͌Sj����լZ(ŏ���Aw  ���7v��3��	e'-�o*���"p:�wt2����Zɩ���ǧA��D��|�K<�b��t\��������D��{ᓼ&-�1�s1��9��
4 d��3c���R��ҢTTM0TAM�ɢ�"�X��C?+�Ja�A�gⲹ��-T��נ�N~�1IAw�{	�[���{V»�1AhhNQ6���I�Ջ��D��DB`�+?��Ek���ݿd�pI��aSj@O6�}�n�K��گ��zFY��?lU����c���k��X�~g�Eq1Z�%��ٴvu�S�fǟR��D^�}�xiMulF�� ��͈��?��Z�㹹ȁy0 <~,v�QN~,��v���}�z���fh�4��|�l�p��QRM�B�w��]F{�r&Ɨd���6;/�f�P�Y\VбN1z�P��|*�ak�i�h����Ϗ������r1�G�� }=S�xF2i�Y�ϥd�cPt�8;�Z7�� @u�a�^�ݢɮ��EG�B���L�W��2����5�\d���8Bi\T�σM��g��A���G����i%n����[��1�2�qiCc�ݒ���J�#&�Ӵ�3�{��e�A�xe��[�|-UKG��rh�,YF@���X�)�Vm����&�T��S����ȼq�!�u:!�6�x�M�'T���W����&8����˘@.ѫ_�3��"��s��㖫ś5�#�0�g�������ߢHk:\�>�H� 8��y)����`�G*f�֑�(�h�m�`�k�f�tUx���4�m� �g��E)B� �w��	�m��D��+l��s��⨊JWtT7rSu{�,�$~,��XXoF:��pZ��К�_�;�=��~%�,Y:&ɝX��V]u��o���5��=�чJlFG5N�4���f~�H6���j÷;�!���S����-��;�i�����(�Jp)RAxl^�о6E�{/a8ab�ܒ��..Wk���*<?�py��O�e��^{�����[�dPah��J��n����a˫`G�t�w�ғOX�A
R�8���`���X��O9���Zw���n!eZ�A
o�א֯n���W0L����`��ג�s��mZ��!���� ��
NqX�ȳ�+�Ő��� 3��)|^� ~F:�f�K}Z�R�a���(�_��Ysk3ǜ�:�*m�(T7��#��B�G��g	1ߋ
&���n��$�2t �ѱCAn����$�[�n��[�*8���G�U�n&䐋��XU���<� ���>!�5���A�>6��>�O�ޤ֘爗xZr(/���^�$�/�G���wy;��r���s_pA}ǈ�,@��MC�����/H��~H�m[�k���s8�@-�������՘]�W�o��D6H��>��{�8��J.kMo��=��m��1����+x���8��DAш?����u�=�Lz��(9�~ؐ12���Iҽ%�����Kq����?��蓱|�����"r&�zg��J�]��~C��SI�������[�x��i��r�+�pP����'��a����HD������rj7T�M]�"@F����j(��v�d9�/��'��|���)�0qѢʵ�����,q�i�ޯ��!�n�S�� �E�h�^:mXOD��s��u��>�	5��g��
Ҳ%W�\sYa��>S���׶�YON�
"�VjSݵ_��Jg�������ǫ0v(��!���_��	 �v��kB��J���+Z�n�����y��yC��*�����[M�W@а�LKj�6C7����Do��6?�:�dw~��(=�3h
N��u�#�,�Җ�q"%�"Z�ˇ�-�c�8V�LP���#���?n/�c����2�Ta|W����#qR{�Z����A�9����x<r%���JC}U��'�V$-����C_���,A�9Z�0iJW�)�5����H�F�0Z�Y/�����[��+�Y��]�2���23��N���w%+N]�'K��F�}�n�����\�#t�A?!}�����0�wJ�<
��DZd���aj.F��{u�~}G��u��w��Պ�l��5�S�$�[>C�Z��n�9���OE�ю��F�e�d�KȁΜ���/ L�	��e�����g��)���n�w��fL�����M��AA�^`́�E8k�� A��>\�U����r=���+3^�r����-e���e"�x���"�e`s�]o�,���	��Iﶴ`2���IE��������׮i�U���FY�p��fq>��LY�]V.��^99F�Hv�Ϗ昅�%D
9a��ۿ�Hυŵq/�Ɍ��V�Ne�q�9�w���`�`b�J������_�"�S�*[�>�Q���O��Da4�M#R������5�bU�@�����	ǤD}�s�;�c⥤<Ƕc�v�2��o��`�!!�� �1*z�)Ą�����7�^���(pX��W:obh&�K	�+��"����k.��&KP���z��胎�� 0_�?zҤ�w�������y��J<�Hg,��U؏�|F��<�E�r���[�	 ��P.N�?��!��.sC�6�WQH����D�7�p�:��P�d,������?T�P���>�	%R�N�K�U�������&`�T��8�%�Qp@��Zd�>�������|]zҢ�D���U�z�ݖ�x&J}�5��b�X/}p{�Q}�-T�VÛ��Ա�h|������#��QЃ�P�B����޽����g>�u�ض��x	��{}fYqc���;Ÿ|t�
�_Vf객X��L.`/�n���~�A�ж�v#Ws!t?W���6��D]^ǡ8p�ra�4�똫�G�Й�8�m�g�:��O��#���~��K�:q��>��A�c�+0�@*�9�U�O��N:�	�ۈ����EF�8�|�W\;��7�|�sJ�j�/�`��Ng8��c���;�յ�vK�>Y�i>��/��\s�