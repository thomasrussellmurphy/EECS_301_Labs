��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|p�n�U˟��1��|p9I2:7&01r�
���ݭ�?�-�|�<)�!<7Itā]�̪���?�~l�Ku~�]�}�:��
lf<����yT�j�$��Z��Y)���$��W�n����QP��%՘�,���n2��eݘ�
ʙ.�:7����7���:�B���c\lδ؇�Ѧ�(L��x�&�=s��<�nVHU�&�,~ݜQ����,8>t��F�j�F+i�i8�q(�^=C�G=��s���+������犿Sh+��ܲ�Ν)h��~7#���+d_̨ 92�ǋi��Wݒ�ȞA푠���sF-�Pp�ܔ�*㲕[(->Z��*�MΈ���5�\�	���c�1;Э��dK��v��
ςK���:��8�6�=P*��O+X�-��0�gnm
7u�1�h��߂i�s/ǧ�NL|�d����-)���I�a������ǎ5��R?�fX�%\Кp�����o����\NsF9f-��h�;����)�\�KZ�ڃ*���EVi����~����K§ꆹ��� v5�wg���"8R�b��r��Я��f	�!����!W����PP�=|)�l����O|2��;�gI2�i�R������z�8����V�(�iI�"��K�Y��"ٽ�$;/�SQ����XLpp�xv�	��×r��`�߻s�簬���m�H�償ض�7"� h��Xݴ��:���:��X�2��O_�n�4\��-�!{���9�ͦ�7m�BŊ�̮��:0tp7����](��c��)��-n�ԶE�ąe&�K�P�1�9��`�9~��5��:LQ��>���r�4�J}~(�aޟ]ili]��}">�d|�=͠���I����c �G7�:	kUf����+�����ԕ��E́֎'�8��O�9jj�$+-'��>��:����jS*��Xf6	��ZZ=s�k���ͳ�N;�%/��`��_Ӳ�/*K�O����Iۨ�f�XH�"��#t�Ǒ��ksa΁I���)�@�V� "����~8�pJ&p���P��`9�{G���M�!�&Q4�A�y��֊S-���X��Y�q��Q��f�Ѭi������%�ʯ�ǀk���@5�9�g��d��^U��s�P�i����ρ5��졻5�q1?�JKd��ǜsԝ8�%�ym���%�&��09�j�ãv6=�����}���շ��ͻ�I�ap��g?��l�x���l�<v&;9�WM��N�Y�X��~��֟'�#J��y ���ܟ�h�L|e�m��x;]��H�Ԟm|u/�j�7PR��T�<D�q�Kw�W�0�B`@J�"�l�F�8����~ȋ\r���pJ��Z�*���)��<4_�a=�������ُdB�ҩZ�)�������g���B��#�޳I�1���U
.#�)_I�[��" �L�Y�A,;v�Qx�#3���D�ŝz�� ��A�0����"=�7%Y�LPp�Ge�b���]�P��=������CK�����Z]-��_�yt��x��z�؆u@�!hE�����[D�U�Ε��ȱ��Ӎ�z����KtfpNf[��~�z�En:�8�Z@��ׯ4l���WPR�g���$?o>I�v�8���d�<[[��s�6�@�J�����Z�}�K�#Y�����4#��"�d_�e) @Ј��8��F�L{ ����/]�VG��'t�x��5z�卙�8ē��u��|�k��>��|} ����!��NfȋF�(|����,�/�Z�GV=sx{�7.O��@��v�)���хB(L~�l��@���7xK��Ԟ<�a���x�Mr�o��	�#L�� ���(��_!7���)ԋ��9��Lps-8�{�g��wg"�������U�`�����%����(	T��.WȂ`��55ͪ
�ϳ��k�l�sQ'�lk ��!��j�Z,�q$??�m���ž�c��|��Nл6���T������HTb|��a��R�0�=�^�ҟwmnBi�-��[{�ӄ��4�	T֚�����Q<n|��7��Sf�8��t��>ݼ�e�$��n�#_�����@�,&&m�ؼ�����%CT�,�����=��dF��G`��&�tM���K�K��!��7�!o �2	U�n�l��f��h���a�*��hP *t�&d��Fz��C�a���`·�P/ �~}�@z�eÄQ0��^i��Іy�6�E2��Ђ��v�D=�qXL���1���奅�����P������G�JO��2��,��:w˻=|���nj��G�g4�eo�a|��KAuO���,��$�>?�{���ln�X3._�M�	��:;��Iʊl��gq���9��@fƃQ�0�xs��\��E)6�.�	 ���:�?���*��2+�6�Ț��Cm�D
��g�i����f��3�H�?�V����^��n��U�d"9�-Hb����߷A3ӓ�H@d�X��4H@[� �9�ѣPHy�d�.���V�Of��5�}����?�#0U[����	�f�6�ڸ����p��a�}����>���
��P�����M
�szӿ΍��ڝ�Ǥ�oz�?�x�*.�<!�&��М*��tU�d��0(�jF���A�|tB��w�?����� ����Q���:�[iaOpT+�&Jɚ�NK�J������3F/Dw#=��["]n�Wy��PoM�����H.Y-%�!�$5
I�wS㼻tb? ��1gw���hr\�xu�����2�rDD���;��2}�]������7n(�`��0)�l��&\Ξ������W�/P--K���0bc�b���J�!Y rR-+�`�Pv�����`���2�>҉w�S��7g����3���yi�v2�`[���*�#�)r�e�9z�)TS�m<"Ǽ�Р�%�Qm_�UŤ3���Ѩ���f��Sf��+>��ЫS��v��\��,L��T�x���+��<bA��dµݬ|����F(>�����AJ��Z���0n���)%,b`�h����0+�I{XW�Y����P�B~ISb	�E�z$����fD�*n\�����hsqv�HL?3�{ՄR��YaQ^���T����q�6�����[����@��k���{�p?-xǻ�(;q*E�y̌�k9BJB8�Ѿ�I��Ȝ��m[��d&�Љa�^�r&:��;���	��f����FDT����d&������[�5�y��$�~�!�����Ɩ��F'��	1�}���`&BO;Pܣj�S�OM[�Tʢ��)q�଑Ο\��XLÙޔG1�Q��0?�wd���Hx�'z�_
�3 ���)�8r�}�������ɋ��& ~4K��2����j�����e¹wi1��E57OL37B�9Ȁ�7NJ�Y1@�#���+Py����a*����j���r���Q(����x���b<��dP�����x�Q���M茁mO��N�<e��4o,�3�����#�]��fcnm��t�8��1�r�2�	Oo�'���S�Df�]r���6=k����a.�����h�%)���
t(��!}���U��N���i|�D�Z��g\�6ʧ����]Tg�!�����`���́���?��dK��@:�@�z����s{�7X_��Η�*��L����b9��u6\�*�!A��Y��3���B�ҝ��
Ĳ����l=P5V�"ˣ܏L�����8Ȗ��E?�AL;j�Ih_�va@��uD���J I�}.*|����q!�e�f.j��X�wۇ1O桵R;�r�@lg��΍Af�tg�j�\ ^��^U�a^���d���P��P�uDH���q��03Fc1o�ϴ�R��������+�/�W$=W��fWZ��L���*��e�Բ)��[b�m�@y�s�VU4 v֞�^пI���j���1dѯG���b�����4� k1��1��"+�
{�������ܽPh�����r���|t�$���>t��ݖ��%�YIt��v��F>YGvj���bkyGJ���1~�+�y1T����G��p �GF��7~�6'rX�ɾ����5]��s5����r�r�vH�W����5٘����U/p<���b��
Cc1�eW�i�Zb�VE]+=�5�FwJ���0�,�9wD��U/���O�<@�n�3�9���$Ӟ�؞��&@��[?#b1�	�:���)+֗ާ-s���kM?8��/-��tn*S��؅���}&�y��Ȟ���O�?��̖�|�=Xw��%��=�'4z�c��5>=���!�_O��������h�4��]T޲8� ǣ t~Kc��=`]�E�lOН�i���$���d:K��t73ѕ��^�� e/Gٕ�}�E�\:ӳ�v3D�=��5P��?�����pW�)�P�������;,:H�]DFA>:�{�$��y�eSY!.;�x��ʸ�G��aY
���ZN��)���1 �-�u�K�`
}����9���"�m�V+�5zΧ1i"�p~�z4z�xv�k	�LAx��0�2�9|��rB!|*���ʟ�5��n�,��	M��a���E�:�,0��^�ci#�>�����C-T� ��q��eM�:ó�]�k�M-
����M�<*W��+i*]"��;�*��B�/�}�Ԧ}"��͈ C��zF�-fs��t��>�^���)��㓷w�}\�'P�X��|�q�\O�\����؈�����/�⨇F�`�!�9��S3�����eױ! ���]�V���M�P2Y 8�I�)S�g���z6��!�I�h'�Sa#�)U
���v�k�*QЕ-L]9�P��� � ����j�h9�b�Gj����D(��%�r��U�/X����K�BFd�-�K�Ŗvt� �R��h-�vP�38�虽п�-BX1.�!KY�����3�������@<��|���SÒ(ZV�߇���&��]�L�~Xk=%y؎^����l&4^�z���1V���}����v�YGW��r��#^ǮL���mPítI*�ɦ��@��Rq�˱b�lr�nX-%W��P9�؈��??��Y7%�cW����fn�D7�	���p��Œd����t}yTd߽�������L�.X�."��w楮4�?�4h�[��X�\���N��}p:�����}�(�XŻ#A�����KR�<��;��'n�0B��|`���>?v�Ub �z���(����@R��8�;<Uf��i��1�<��p��!Z��T�j#�jS�Fp ݺ�M�fV3�Ol#=��i���i����Q]�*��m����|iF�4������O����_�$��΄��B>1��,{9�vZ{\ؕ%�E&���p�I�T���/�C,��6�i�;W�W24ؓ��\�c��c�vɭl,q��c�v4\u��T0�1M��K U'(G"_�TG�J�L]"��xxx6�
�TA�ޖ5|�z���:+�jQ�
̅mSt��?a?�,�� J:ݩ�{:K�U��X�0~��S2
~��gݞZO��0b�">\��d.�덀�'gc���7k�����}�pRJ�l�'<V�ɩ�Q�M\�F+���σ���L�4[�I\SF��uv1�5W�lħ]��k��	F���Δ���_p�B@ q�d��*ha�1>�<-�6C�7��W���P[��9��W:���	Aq�IVh�y��}˸�=�p���Re�$�PAm��\�u&۽�
�S�BS�b6pR�̂�����JybĮ��|}�\�!�
�3/a
L�)@󁛊�!S��ƫ�.��M}�0W;�Í뼇i	Xy\z��7�O���{	���d�yO�i��US*�N<���/�VJ	Mfz�ЦR��O7_<��b/˲@��f�״+�^�j�%>���I�`�:��I�#�>�LRF2�,��O]����)�Ul6���\"U��!�����
�h���p��2��	�bx�S}kE��1r��7<���^�j0�)�?��+�*)R��Oy�� �Z�_�Æ�&���?�]� 1�</�;�>-[*�wrT������F�����;��t_+9
���k��׎\�h�[�apw�N����NŎ�:�%ⶆ7���bw6yb�:L�WE��u�[4P[k[�W�DkVr�H[!A��&��T�K�P!ٗEY$�%|!�?�(f�������>=e(�(!�H�υ�eg�Z}�jd����ω�N��#����?��c@)��2�@g��-��'��+��d���K4�[cXh�c֜x��q���!��x ���S�⃟2�Ɯ��a�WR(�Z�Ѷ���곟��K `Þ�_����]/��h7�w�@�Q�p	�C��A��j��_J��vd�ה�cf=y}qܚ8����B�4�'��I�fӜ�7���g:���N��u2/k9
�D���dg�"Sk�%3�����:�Uda���Z�dRF�ƘJ�`���20�E������!��0P� �� ���L�2�D57E��ـ����J�5�@�B�8z2��p�3w$l^7���Sf�WÓ�#�����E]_ᜇ�ҕ��i��x��H���&��+e�d+�A���4z���z��x���Ҽ��j�j8XB��j�~��3ܰ�m�A��~t
���6�ŉ�Ѐ��-�@V��$�iD�&��V�qx5<�bQ	}�!&��n#���I3�A3��t�6]��I��&�c���lz��~1kH6T��yg�Pg8$���&���� -�f�׋{g�b��y�)�t	��s�r�*�����+�ͨB��HmU��(7'��+�x�0��E��y�O<���%�XDY#���nƐu���~�����"���	�.���9{�9�>&>��,[�;��.�\�d0�]������pf� )���[H��%�''<�!��AGl�NT|9&_�N�ܸJ������9�j3gFj�n�*
�΋w�D��5�ٌ}�+�@��L�ө��O�2C��Lj�-�,�/p
 ��4PrS�����c*g�`��	[>�z�b��r�kS�r[9��K̍�2��S)�9��Sp3�#ȱK�̤.���D�{�Q��&gpb,2�ɟ�n�� L��a ~Z���~�-�``=�;��,�I��Tm
�� "��1Tyj�����`�T$�!����g�{�![
>�Q�$1m ���v"�Q��<�r�I�a�M��Dy+�U�mbg���}�yj�w�鈗�桔�
lS+r�"���%N<MX�'����o|q9�.����2QH��!ˆ$d�Z��)-��2z�ۙ�ļJ'�vpkm�����@��|��L�T
����Ѧ�J$��?f5���TPM����D���8�^��.u(0�*K�����g�H&�\�@(|�!�׺-�6��l�!a�׈0�Z�f���?�#Roiɔ�#����وP��.�(��ꦃ�\aO����W�s��3��L��K�g�8�����S(���RJ��Q,��7�$�*9���	T�V�����|�ÁQcɯEUA�<��[&Q�}� 9�eB"�n����Z"�M���3S�wֿ�i��_���BE���C޺���vsY?��NX}=Φ��"��i/�|�)�'!_n���b�]!Ѽ'��M�$-F��=�}�*QCQ	�şl�l| z~�+)"��d9eh=����e��t��Ť��vS�%�����z�\�݃he�3�`����� �o*���ov]25p�l,A";����L���'�D����zY�'�T�b"냙ԓN�������RK̨p�hA���㙀�zt��+F�/bK��$�c��÷�/o=�pڍ���Zs�If^����m�Gs�HW�������K4۾N�l��X[ �$�Ht2�:U�@�p�{��}^R���V~��]��Ҋ+���7�&N�lͲق9��'�:�`�蜴�-����\�vv)����W����%+9l
�ca�#k.k��n�O�3����/t����XZ��)��o4�"��B� }T���3��e�.-�^p��d{���Ed-�B���.�����!���%"��E�����G���똣�^L�[~ɏQz7o]�A����@�!*��v6?"FB
���Ş�m�P?��찹Vn2��r�������'����W:t��G�1K�7 K^@�������J���b��)����ьK+�v�+��4��TѨ��ڰ�?��$��K/T����|�n�#y0�1��3W�X�I������)&q�� �e~���MH���]��]b�V�2�T5ֲ��O��=��pMQ����w�-��{۽�/�L��kIr���Y3>`)�s�OC���n��]W���Φ�\��Q��O�$�D��5D$B��v��a_^D��Μ����t^kb��)ǘ�챍nh�~)������d4��\ JRHӈ�D��1���ן�؜)��$䉲�"m�6^C�O~��g߭En�3�]��na!���:E�G�)����#[�ˠ�3P�{��+��O/��'�ՉS\�$S0c��'*�&���`f��Fiu:Tq>q�G���q.;-d��+�T6("o����rR��Jd�0H*y�F�웢��"bV�'&��U6/� M��v��j+��wRAG#VG@�h�K�A�I\��@��#a�k�>�6�x�(������<�������(�0���y)��x ��\��|�hl����`�l\����Ve���#��C"۠O�uI'�����Bd3��G{i�U�N	_��\(�d��N�:��x�B�q*��cȮ����$�Z����bŅ�R��H�}d��F��$�p��'<|Za]+��y'�C=����}��*h{���Pkqy "�S��dD�[�{�	�����˝�ς���,��T��U�����c�P&;X� `�Ԙ��8	�sF����Sɾ)2"]c$�e��(�/��|�})S�L���\{�8�9YՋ�� �l�\σ?Z�u]lh��`�Bp�g
���ށ���I��!d��G�8���x��.�+{G��fZc��g�B��Ϙ4m���������\Z�f�u�F�q>S�	�d���@䀚����0A���j9a�x�������h�7����r�$L�l�JO2��BP���~��{��в�ҝ��5��cZ���9];����#,g��_��{Aݐl���,�@�]͞��W��Z
R_���j�daM����Ǖ7�Z�kh���]���|v����},�%8�n W�y'/�5��l6ӭ�9I�ۻ��ş��1h��[t7��~9)60���8��:>��d���	�q���f4��e�((a�va��%.6�߭����[w�FdFa�Ƅ>�ʫ)�ޥrb�&<�i 6D0q=N��"�-�Ɖ�t��_�5�Z���@Ha��
��T����8p*RJ�lkݮqT�{��|U��i����|��Ag��]��2�_�A>���ɦ���J�jw�Jg�(:��}��fh���=�_μ�M��9.ks�̞E�Q�����꒒� ރ'Ƞ
LG�RBo�����)�3G:����|8�9�#����b�[	Q�iMN�����5}��3�G�����3H}<�jF�g�Rt�n>�/�ʠk�Ø���p�:�g\,�0��S����<4@�
�?h�T�o�+���=�e����k�`[�*��D�ĕ���ч}���B����gv����K��[Xo����]�0.Cr:G_NG�	
�倈����?��l7�Y�h�F�i�~��?�!Vs��3�e嘀�roͩu��� ���$��@*3G�_��ҙ���!0L��򋄰��*�مީ�Ѧ8�"ȅ)ųZ�_Q�%�zY�=^F��%���OY��F�,��R��(wy��@D���;֩:��(2��CǸ�f�9� �+���CL�*1௲�����&������FXD7�)����M�|͔������)D�Q�P��#Է�/R%z�I�ͨ9%�Mpu6�N�ս��%	�GU!7 $��"r����҄u���	:����U%�	�Ė�k��(w��{+�٨�o��^bI�&�k��_)�F~�*����ө	�ї���v�����Z�x������
��|�k;2�6|歑�h��T�;?�YC�+���6���؍��d!�5�1�B�)-��Y[��k<
8:�����n��Q�Y#��2&���|�eޑ<;rQOJ�>1�A��-����u<p�ɸ�H�w����97ѫ4��i78��{oR=�
��XEzi�p���\߯R��4��AP������UC��n�m�����k�ި��,p��h��q�w��PԻ���-T���}i��!� wF;�>����/�}�V�5P$=���Y5�Gr�۠�^t�����c��s�Ѿ�_�LΤ��Bg�<T{��S�o��_@�������_ %I�%�<�%*zhD&�|=�a�;��Z� ��um�]�^��,��[:�Q�����T���������햢������0�5i �^�(`���j���a���΋ �>C����0?�
N��a0������sV_�D3��)`4��f�QP��CifC[�z�b�K�&h~0�dT���0�Q�%fP$�kt��d �H�/����14�ޏ��*8z;yq>H��;������;����[�+�)���"&���^։)rOb��#�Ե���;�.������]�ր����2�'�bd�%�a'��veiZȱ��u�+�70���o��(I�'+G��3��ENy/�޼?Y?-�{�c�i�>�d�󿻒����] ��Eڗ��������i9��*���Y�'�txxG�Qa)�>�oCzU� -+���X`�Q�/T��s�ŧQ�^���2+����ѷ��1!������W����Yi�5�����~J*7���!�*cƭ��<`V��ևT-�ʡ ��]葄xG��/7Kк�Q��5��g��u���t٨�tQBlQ�����^�O|O� �x���N5¦'Gc��<]y����_W�? F���Trw<��fìK�M��h24xo��z��/��7sc�o�I�67�mG��2L�}����B�B�C�jح��/�,�Sė�1�hP3�F&z�����e��X!�!�"��\,չ�#O���H=�]��DwI���D�Nn$�ۼQ��b4�T�,�v��Wc4֌�Kܲ��Tkg���n~T���z<(���vU�Wx����W� ����i�U���p���,TD[v6f�%�q�M�q�HL D\C�e�̔Zw�L�q���B�����	D����CМr8D�c��F�9]�����@��F���j�үv���qOz*������N����Jў�x����{ { ���D0�N�����~I�*�%��!�(�2.��q/�aT�FɄ[��w�?���bw�q7=xd)�k���&E�8>	��3�k���l��M���Q��T���nj�֦�"���9�S�疟��M���κ�e9�����iq�I��2�N7��{��m���C�9�	�
LU1N�ɇWc�S�¾4$�<��7m�!XQ��ek&֬�T�4�w��d�|\���,�Äһ�K�$8Ǚ�hBْ���J��H��XL�pcxOO�c��N�$ra�%�&��Aw�A�x�����զ��K4p�0fQ@����ǲ�C��!���'��Q-�ke���חd.���U$��]��ǐ�e&�ʇ��/2%��$O.�%XZG����1��'l㎽�+$��9���6�h�ȣqK��3�.'t�e���ly�N��uQd'�OJ(J�FvB��8�h�n#i���cg0��]��Ro�M9�?I�T��j�ů��ě4K�pr]^�c�33�em<��6��Y��t���HT�k��2�i�Ā����<#�JX>.�T\v��n��n3�N�������t���N�!U�1�v�k5s�!��}������*�V5ڮҢߊ�t�Po4�a�ľ��J�>#Pu|�ha�v
��D�"|�TRp���d�v�+��/�	��9uI	��@u�EZ�P���o=��-6q��������J�d�$�z����G�¤��Lm�1��爎�q��m+�>$A�8doX�P���L�	�|�l�X(Fs�rxIg�Γ�O^��z�h�Z��u:�$�t��=�z�>�׺��eYN�bW��V9�A�-��x���x�*�r)0���� ����Nf<�+��ԵȌ��a�\�RY��3��p�]ۄ��b���pSUk�zMٍ�"�(v���Y"��±�EX��� ^�������J��b܁=��������5KW�4���PH��ii��KtR�Yu4ʀm�J�V3�H�aJ�&�4c v����ԋ���c��&#�8��ҝ��|��KJ����R�v��,�0�
F1v�>V�J^����S��d-�צ��M��a'����&w6]�uzu�r�tX,^�PU���9@��s�%;b�o�'��)`�'C���ܻ	.�B����K�U�Q���FR6������l��3�ϯ@�c�{NN�PF��-Ɏ��.njD��Zql�"12�,��A�SNj��J0��?��i�m\/!0�P�F�p�NoKp4��0�ӎ��!�#g���7�>9�?��"��_��{���%U?�Z�!��C�a�"�G�фc��K��n��qK�r��E)�h��	��ӏ�aF���ZcP�I]���Iur4�zH���,|������K�b�R�'�dדv�B԰x�/�K�ʝ���Q��R�q,G���u흻8�+��~��E��'ĕӰ1�~�Fhն�(�e��oH�QO�迸j)'��
c�~%w���� jU�<�+	�#���^�\�2af�bv���Qm�_3Frv��ΧD�ʗ��%oo�ٞ#�d�0Q�i��G]�F���l�J���us���������F=�c`G�i��m�n����M.|�3'"�7���"��2u�Y�[J�pK�y�����J7�;������/͙�~:wp�&c|�3u'{�Y�Xf8H�`��7���-m�*#�{�Gy?�L5lqs%q�����^! �����[}Ѯt�{��W�I�1u����B��C(o$�`��2fTbqB��N��s�rz�����P�������3��r��� .����s��ei6���2�fI�dK`ې!AP���V�I��Q ����~̔0
FJ)�k���7���
�ѱ�h�r� 0#�{S���l&x�;��w���`����ɕ�X�����DP�<G��Aj�u�� Xf�B`��!�����ف������-+Z¦f�w*TPGQ&��/m�G���i��������G�DX8�W�ł��K��;H~D1��<�١���� J��VK�`4a�O$Ѻ.2�E������IC�"�%h�*�Ǹt"jN���+��Ixi�UΘ5�}1�� ��e�P{:�R�}M
ǧջqc ��V^��������Y�`��H^�HT��T�q���h�/t�)K�c����dP��(Λ����%�����i����L���<���G�m^�����Q�_���w�>��U�l2����wK �X���{��ꩲ���x3�g?��S����1��F`3���U��8�f��C�j�|�}֕�mO2�8�t��˓I���$�ACHVLj(�c��(�%��h��F:�^
����� ��jJ�V�����(�Hw�V�H����(�E
��.q���Tdp��ҪD������@Ꝧb@��Z��;�{	A�p&`� }�'�<
�{�����M{�GB�k}�_�ObҌ�˱�<$v�3C�43�Z���C�_Tu��y��%7ڈ��RYY��))��B1A�KYGF��Em���bn��Z�N��{&SW�wz����A��y�CAl�=a�,����Ԣ��6w������S�>@��޹ )�B�=�^)����	_)�۠_(�Aʙ��'�4�%� �� $3=%�)�,0P��Qz��f8Ka�ض�i�(c�Άsde�����|a˪y�n�J�6	�g�4�wkHo��Ӭ�&7{R����u%E��F,ĥ�s9w�[=�iU���9�=p��C؟����{f���̧���V6���t⿟y�T�E�#�^K��K=(]�����4�/Q0;�)����chF.��!{ kv��E ��K���?ˆ�c��
r�ǻ�*�Y���@�W_3ڹȘ^���25rW�s�r�ASh8{��gs���,�-�	�^�}�b+yzy��@��;�[��2(��v�����u���Z���g�l��"�=�&ix}ٓvʤ��v�Hp��0��?�9�R�ZVW�7
 �	Y"��f얞���P�l{��.����ed"y2	1��h,!�4/�D�^�-��=�w����F����h��Ԃ��Y^ճ}��{�e��@!�9����i^sؤ�\���Ϛ��+��GT�J�&?��c����fi������,�ER��-/4p/�Qb�4~�QYT�����?C���O�K��Q�R�%�3�lw������db��4����
���|?@��P�����C��KbZb�,�j'��vP���(�tO�?����wK�D;�/vDl�v.�rp67�;�c�V#P����R�����X����R����H:��Fg��SH�8y:\&�<�������ooTv>�k�P9�n4k������w� ���k�. 	�?&f5O�f�ױ��}@�9��I�!�<��J�`�DR}좶uE�a}sRV���@�W�[
ɯ��>����'�M�^�H���5����`<j8���&��F�&=�Ad���T�(td��I77�S��ȋ��Fڝm|{:�C�Aο8��Л��v[>�c����qWo���0�i�6!��{�D^TJZ�� >Z�eʙ��L�u��_�$��]����5 ���I�����ᶙ����e��{�N�C&�L���F��~�L)� �u����o=�yQ��r ن��M9K�z\����6�/w����g^sSSsA��)��.S?s6�&T��[�������3Njދ��v�-��in�pde$W���E�t�hN �ÊG)'�J:̓n͎/�����Q����S�����_O~�~D{�~T��݀I�Oߎ(㣯g=�?ay��a*�{�"��X�q\ЊtÄ籷�ySNoU]�U38��͸`&���:B�&'�g�� ���Xe%�#;�$2.l���j��Q�QʩDK�i����^fCU
�!>�ڣ�|�a�	��.�r�K8��_�a��`4�_��e�|�s�ع�ZYЧ�g)�Y&N ?i,�}]�{O^׍x��",IE8���\A�Ѱt�'����#��}a*�;Q=,��S�LI�?�NV(X���=���U��a���P:�8���[nE���g߃fp�����lß��Y��J�������2�mJ0�'4������o&�F�}Y��������08�r(��:H(��hߔ�{"��x�R$�O�7���Lмw:V&l����6�Sڲ3�,���<���dh��c$�b`�
��(E��@b��>*H�8FN�-��="�Dsa�0n�m	57u���	����X�uܒ���',}{�ǼӘ���R���w�Jct�ö���a���Eh�ˈ��e�����ƣ���.�v	���v�P~œzkL��3,qU�A0��]EE�3�4>��yh�Ԙ���s��Y��������A�W��7+4i�X���	�I$�ތ����� ����ᦴ"�g�R1�KsqO��P۳Eۘ��ak��0(���l�-fǐF�){�b���gw��tv`F����	�|k�}��<��7}YQ�f����%	Q��
�f)C��QV |�%D�� ����,n)��7�\����*�kj�%�����t06��QZ�:k�Y @8�lZ���3c���x:e���]M�15���Uy���*$��t�D���q99p\���P�����5-,Sd�UR�AvXF��N�f:!�
j�g�����m�u�'d�}��-�(1�v���!GJYa�B8M�,1;U�TWK.۲"�J޹�.axË'��c����kR��Zd�e���FH<ە�	��X�G5[ ��]PC����t���f`&�s�\}��t"_=eK�}6eC��( j(s�d�r���٥3qS��vtl.�t"�k�����N�"���$�G@@�Q�F�
rq����'��Py
Dn���R�T��5{��+�l㔽q^zPF�h�43\����/u��{.���j�mad͌�{����F��W�Lw��X��9��s�SHc��E�������i`k����ޘ��kRͮ*_b|8�܇�ui�f��3����$�Yΰ b�~.���V�
m���'�BCI�
?�q�z��}0�Nxd'#|g��vSԃ<���ײ6�����V�̌������LW>�D��)i	7��1 �F�"��2�0�U����s�����{`�,���v�@
����ۃf9��8�X4mz2�{6j�(�/�	�������fm:KΞvn�6��XO��7!J� �8�q
sP�)�'Q?�Y;�!����#�o��+fS�V'�N"��3��.�M��ؖ�DCED����-����Yjd��q�[4kM�òhp�JD��J��u|�gpne��6�O����J�n�e30+����sO�f1�	\6�ٖ^�s�l��+.J���ύ������B��W�>%�����s�ݟ��9����A�:�9��|+�*7Av���vA�?�bU�-!�~�fҵ�
D@�lp��O����4�e��$@l�y��n*�o����N"�yCe��-�{�!��)XNK9v�E��5ǃX�լ�����3[F�����aQ��:�Q-CL�X�F$�>%�m����|yE�ㄤcu�5����T��{r�T�k�BYO�	~>��'�9qα�F*��Q�yR��EW��Gy�zr��끽"��#���Y�S�٧L���@�U��tŹ�ѕ��E��Jg?1��o�˷����yr�:8J� ���l�$� �v�����wz��h���սq�gL�������������I��q��;Sd1:Q�qc�����,�}��J� ɔ�. ��yU�����D���	C�A4 n��0�f�	
 �^�MB��e�c����!n0(��0���8k�LK[�ۍ5g �
� ��^f."S�*�x�v���O�Q�@D�\[֐�"�
��s�x��y4ۅ�]Ž���n��ã���-����o�j�SoU�Ϯ>90N*�%���f�����KR� ]%�X�[�n����i�
 �/�;�̅~�Bt�O�{���=�54�(���|?��=k�[��5;L�}Y�_���fj��&+|\X��o����o��;�����W� �/�цoG���B}$v��vj�=����D�X�}��8���m�[?88��&�,F�(��lK�,T1Iv��eKh
�������R��o��h�0,�����2�ZzwCq.�\,�6l���$�<�ݿR�Bx�b����x͵e(cE�R�%ا�Uj���F�̍<�p���$��X6�O�;���^%u�xN��m*��q�$\�b2�IZ�� ?���,�n��{�d��ކ.�S^ LBQ$I/%��4;V�i�qR��Z�E��L���ъ���z��BN��ԁ~-�V$W�I�MLk���DX�З�*����NL"M��j�R�����2�L�ra��]\����:���c���Y.��T��O[���Z0mk�S:��������6_��ɳ����k(r4�
��V�?���/�*�8��f� -�3��E�����Jr���ʮQZ�o'01��1��}��5<'��%n8�����\ܩݦ�wt�����AV�M��7A%}R��+�����
��N"jm;Y'�&i8��˞�q4�[G�ɴu.�(6���P'���kf*g3D�) �dϡ~��L�J�-0d���U���cl��Yg�l�o�/�w-�ZD�2#	�u{�F]P���:�X�;Nx+cF{QY��=ּw�)��ˣ]�	�=��^�H�k��%�sj1���@��E]x� tu&��I��h��J�V�=��_�x��
�V��]v�c�����}���}�ɓ��{����Gє� O������PL�Ad�'[�ȿ�>Am�	�ć�����ǚ�X����%�9�c�o���7�:��B���}2L�,;]VdH�e��dq݋ɚ���l�ypR�`�_5�sG7Ce����}�����`%m7�p[�D}�Cr�G哜��25� & ��(��WX�%�+ _��"|��1 ��-t�M�O<.�Q:�J�+0���I0D1�ub⽥��o���u�y��M@p�A��RB'�<�
-1V��(=1�Kg`[#y������������C�ky��N}�y�N7@���ۿ����?}��#5�oI7Kll(���ԍ���Z�d �{ho�TFW,s+�u���B'�2|9��Rt�cNp�{�{��^��%3|�u��<���xϔ�p�(c���̋�����v�A�:�G��u?h�4�f��O�p�|c�qC_���:ۇyf�lD�N9	l^L�N��X}�S����D�|i���3����>4})ר�zBV�1Z�l��S?�f�Ŷ�D�ݍ	WM�S+w]R�լBY�Ȭ~&P�A~@�e�W��׺�����~�[�|����RO�L��-��6�>��<�cbT���ʏ�������=d��{<��h�=-v�	�����٧�tĜu�Ϩ�֭�o_��i�j̟�ⰶZ�J���|�%L�n)׆��Ᵽ�P�9[3]%��"�5�
����Ⱥ����/S��1!��wmE�]��]UM�vG�Je)fG8��Ƞ��i�����F͏C��x���7��:ym���
i���?Q"&X��.�������@I�@��7Y#=���m�\��/��T������$+�/�X]5|�ւ��� ��^�y��� bt局�[}�N����$��B=��i��L��_���?�l���9V���|�M�o�i�.��^<We|B���� {��,8�z�
�GVo�R=����I|��>��G������5l��#��i�I!rŮ���*i�'Ӗ�����C�Y�?��:�M*8��KӠ.c !������l(�������z�%���AC�S2�h�?b/����qq](+/mĢ��� ,h�.�#�Xw� f�	C�&��7��+&�ڸ0�=C����;m�2��BM:\r`�+X�gr�6>��!o)�Q�Nm���ϼ���5�௺������ԝ-�y[�ڏM����T�Pb�v�Ux��r�/��3�S�<m�d��<ah�!�����X�@�ۘGO7��JGg���\3=أ�����3I�\���;��H�.Y$`�����TF'(�����K������\➷]�>������j��g&�,���v'�wpi�ze�'���� P���l�� A6j>�#;���ITԽJ�^��O�+*ED�L���o�c����Ol8� ]/��j$Y��d��^�;�kc��*�Bw��^o����D�"�� �)N�>�|��2u� �7D��$C�M���b�5fFr���4�2�
��I&�̽�#o��.8o;��b 8� RH=y�WpD�ZpˢK��Ƌ|)�$���������UߡsX�Dg,V�B`\U!��&7��k�.S4ӳ��[���C��!A�k�Z�Bf��������\����ٳ�Q��کv:�.��t.��)IQˠ��q���3b��2�+�b��ؼ��,$�h����أ�ʍ��I4��*[ c�b�AMh�vG������𓾺fAD_NΟ'��=�K��?�e�Rۗ'��ξ���:�Z�<7��AYo�:���h����:j�)-�����h�p�k+[��Ke�	f��x)� ���l�8���!<��C��X�5H�%5�_u����.�wDX����e>�d��w�r<!�����r��_`���qM��8������@:��_�L3�w��J�G�>輏���H��7�6��@@�;�o?��uFZяbp��)�N�ۂm��eV�)a�i�P���F������<3'�tz��>��f�Z8ʜ�"��Q�,:F��+|�.%��4"B��q����w�p{���(�}�!%?�4s����2�5��-#�N��E�ج�z*��ΘL^�&#2l ���w>,vCN,��v�0+�ѡ\�T��r��Um�#�(mi�#})���/W�>�k}��v�]
z��$�w����K���%����t��x�V����d�\��#v$��@�ww"iQ�N�B������E��)�c���V ]9���h0��|H���yVz�1�'��*��a?1B�{嬲�ݷ���@0+���=\��k�{7�m?4���N»h&�#M�Ƨ82R�l�k%�0e1g�3aR.HV;L��C��a���=�iC:|�N�D�}d�5��Á�z�,i�ӄ^�*���H!���3]}B�ђG���`�C�pi9�cS_%C��M0nT�ŅS��.B�z�M��FŸ2ۗ�,�Xѧ�N %����@����hViv�K��M9ї�e��m
S����vX-)W�|�F�P�cCY��ᮽ����	*�1Fdd�Ġƴ�be���+��n~�>����AJ��U�!��Q~&�@N���FIBO;����k�"��Y�҉�����(� �F�P�xƂ��\���HMxTn����1h�w}K^n"9���
��z��B��F��6�I����/��؀�G�L�T-�1��F�;Җw�[J�f|���K?ti�o�y��)���|]�@�k�M�q<W�$��1*S�=g��h�(�GS�<¼9�C��`��Nz_V�FV�������z�u_�Z]Jv��*>Ҭl����wi%;!���}J��0'W�lO�YEI&����fP��X�#�"Ƌϛ�<�7G�!���q��7Q�!#h����������h�=㿔���.��'F�bW���.L*V�V��I��K��zw9oW-F,�'j��BY�@Q���bЮt�	��S�Ʒ"CQe�&U��a,(֬�4��͑TV �%����&��,l>eE����0uB�}��и8�I�-`N9���r'
�m��H���/NL�W0RʑO�5 �}@�; �t��a� �r�w����C�:�G����F�:���P�Na"�i/V�����
;.�2�Em����ٿB�'"4�@�!���{�#m�K*x�Ń��ڴ���?�}N��̈́I�{�C��W������D0FO�ڡFT�����vΣB��V-fi�iQ���S�`:н�է �`��q��u�r�?i}��:R�o��#nt�㳰�E!;F����X���l�0�94r���G\dT��e_k�V�&f����|4�ubF<��N,=N�E�q��8B����.����W;&a38���=ݙY�S���T^�`�)���	��� ��S��M��� 8���l��lnyB�m�A�h��0(j���L�A�2'R��`r�sIP0�0Q�J��(EG��@F�(�m�hVQL�5X�o� n�������S�e�]�#��~~�� 4x]�I�����NrS-��AT
8{��n����?���(��i�g��N�R����3{_����V�����0	҂�X5A�����5Wx՝ߺ�v�:�j�=-��S4��譬�����]����}��&8�M�[H�?�.�K�n�ɠX���~�B��R�}�ժq�F��L�M�K �W��Q �7�t�y����sy��u(��;ï�n%�P�*XR(�uW�C���p�o��8]��FWb�����W�ѳ�����`Q̒��MF���\�V�
�o�dR��=nV%���V�L�뚄+�-��$��Jo4@��\�p1�	_+h���)��j�t6����w!�VB����K�B�P궒�.:�7��m&Q^��nT�T�Of�Ah�J���R��7�(�Ij�ŴS������.PR)��-�8�U`Òyc���L�������c��}��������ݗ-�r���X�����`�x+
�~>@x��V���$%�XU��܃��j�L�HQՅ�ฆ1d�$��]lGD��@g�x�|���Y`�^���,yC.�������Iv��/�y�9������T�O��тsfо��n�c�n�yW1p]�(N�3d� ��X�#��b�_+Ϻ��.��+��B�fv9z�+�m�N��9�E��:"��"Tg�^�0�.��U�c{���zv:�j ����{�1��'=*���MZ�g����yF�)�[+O����K����߲͠�O��\��W4�WKxr�i�۽ K�!fYK�������@J!jK� �;'��T��ZnX����ꀌ	F�*�����f��U�i�8�2���c��o24��ĸ������70A��Z�՞�1sg�Lʦ��
{,o��7��M��[��n��A;���Bh��_
̅oN>���v7��NJ��Cy��k��cǹ�_�i��lC��F��v(j�����d��D�Kڬ>��>@��Խ��g��f�g��J���}-�a�G�#a��(�!��K�mt>}!X�SJ�CAVO�4'V^�����wŤ���}�N܈�m�E��E����gR���3�\GK����Ҥ�e�,1�a9I�F`�,_��0`�}]��Muy}����R�+��\ˠ���[�Yݘa���ӧ���U/�U��b�L����*x>@�Q��۟���e�\\�g�rf�Q�$FP�!�X�yl�ҕhl� �c"%�ɥ��S� ������ä�Q_��R�g�Uk�Cg�Y��Ҿw�0��	����Mʌ�?�c���D,Q���E��!=ڶ�ה���x�<�:�	|�;�I,)�8<}m��hX��q�6��-h)Y�I.������q���psS��u �cw�"c4\2*�5̓�O����^�ud�r�`p�	뉮��&��[�}\x����A��/;����� ���.� QU����92^>�@���k�A�&�n�������!koV�11�| ?�Yr�ŝ��Y�I2���W��y���7'^��N�A;��|a���?�Sx��:���