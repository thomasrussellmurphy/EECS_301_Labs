��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\���V�fnvx��ÍG_;�ȅe�~�>���9�>�#ߦ�����Io��\�X�R-�yr�u���z��`��5C���^��G��/gl)������*�m��<u~^+{J��'|{�V�G���R��E�C��}���Yr?�M���V�ɞQ�8�'^mu�'�m�x�@e�'���C�'L��<��Z�݋���J�|80o�A�n��k��ٓ���j��^�P[͒��҂wG��'覶�<�js/�˥��>FH8i�l3u��܉Z�����}B�.��Y�Ge1.{M����/���Y��p9SW�6w�5SХ��2�� w��\U!��I�:oY0�_�e�N��(��V~�Fy����1�F�L�(O��8?���Fy� F�6�����F�cer�a'��[yk������#O.��{���x)��~�%"^�u����`\�ݠ;>L�a6Gvw�f|��.�Xv�X-Y���[�
�H����L
̻<z�����t��?ѕ;-Z�!�oY>�T�j퀑U� ��@6{��h��5���Y��	kO~��;���u�$�F�du�"�����'�(���7h��R)�E���ס��/L�ʱϤ������A�3�ޤƵg��|P��5	��A�_��=��쏱��5���+���x���L�(���.k~���7���!�w��R��K6+��x,���psy��b��_��	ջ�Ŗ)����8 j�i~!=S��f�C�ZPn��e���#�z,��}���d��7/��<�9i6	oGe�����|A���Tɪ��
�����&4��\G�en�k�o�"�GA���>�~����w�U�`�I	\'6������`�K
ڒ�e]y��$�x��Oo��B�f�l
�]f`'Wm��ںg̮�[�w�{���K����d+n��h�m�4{�F��Ѣ��"��v]�h���S����9~F���p�LP31n�\�-��-�Xzg�&�V\	�YD�R�5��zK���nL���������$?F����p����(�ezX))Ջ���W��,;��z�Lw�k,$���[3	K�a��3l�1_��ԩ��d"����hE{J��l	$9� �rی�4�B��ְأ\˺k�-�#��$P?Qf���Z���%�#ѱ��T�>b�d����T�����.�sIYU_���)��˔�	m���b�D�yt��2?�y��j�g+��u���,�Q�A-;�Ď�Z�:j��޵�Ϡ�!�|��������EV\�� ͹X���Ǫ$����CI�V�S�'��PFٕTjP��@;_{���7�Kb�G
9���[��{�AiR]�0�G������ٍ��.8��1��n�7$!=!��TϬ����(����CRȆS(-)Ly4�Z ��Dt��B�睾>0"J�ڔfW��y	%f���!�n��(F+X�_���pM���m�Y�s1������tIHa�E�J,&b�Dr��Ei���%�����R�sl0�e.��-��l���}�>� �!��L���`��ӛL_�����pr��,�����S���~�a��{� 
�'>^`#D�b�7}�{���%"�]\��S� ��ϫϢ��j�t����K�=�L-L;�ʠY�ש�pt�r����?�YV�CoWZ?J��<G�ֵ���ޭ��`h�^Q��x��Z��&���3��
�����nS6m�3D�������V ��\�?�^Ǥ��V���f�8����}#�0�L��G+��)t�*�vx-H�w'nq�ә�7����s�lx�|C2V�oz��X"QS���auGi����c�rw!$�s��D��UW�(��4�����Ƞ�ƒ�����y+|�
>:�3#����	J�f�7���G�{<�X$����|�O�!�4}(=�տ��Q8r`a��6��lh�D�e��D�S��	�v�L����s�&@��R�B�P��YڇT���Ƣf�ȥ�VP�f_f�i�Zp^+��i�.&`��%���IB��щd�x�|�܀P��(�:�_��%�U\&;-�+:mk�߷��pg�0$��!����Jm���Ȼ�p�Ͳ 8�^9�:m�>�?������S6�3��X3�z@��Ƥ���z����*�a��x��Iz�M�!��>��$�Sa�@Y���W��B�CsB$��m�EK� Ɣt�o�Du�rì��� ϳkJ���2h=����c�v��|Z���<q�F?3or�y]#x���$�����M˹I���:�A'� WU�⮍F�ă�n8�t@1�:P�9��������7}h*ߣ>QQw��ЈKܮK{Y�3�� A�S*����P.����`�������i,aQPL���ȷC؄����K�}yC��h�s?��8�^Desm1��5��@�'�͸ENjQ��K��Ԗi�;���";`�zn��scL��^fqZ̮��"�,Vi�҅C�L^	�I��*ުW)0�u៞�F��B�	�3�������<:��$�7scWZE����$�xIE�}
�~U���]5�{�%����gQ��U�+���0�c9������I�݃�d�V%��wy��IB�Z��3��'�w�g���CР���n�ꔵC����{i�mD�lU�]�$S�H���y�-�A�وfs"[���˥����n����#�^�F8tift���؍U�'�)�ECɎ V��ނ9+�0x���#<�y$nP �yO�4A�|d�vщ�oZ_/�q�! :t�<d�?+|BȐ(�?ע�@�N~�c��q�*,1��6P�6�B;)���d���7����&jiz
���չxn�6�����:; ���Ц��Us �B��$��k	��� A��j���5Dǿ�@�FR`�s�|�M���$���ס�
bʖ M^��f0'TxU����X���9�H�5T�`��8�\������C7.G��:�w�����znļc��#�4-4B�Wpڱ9���H
d��7�gW��w.���H�o50歠��ޜV�Q �4QU�� �}��"�1)�N&��ވ���d��VVƝ�)���eA�l���+��Z�0�'U���P��bn ��L�{��UgI[�ld��;�x��$�u�B-.�a�L,e��H��T�s��IC�P�rt��%V5?�����Q�X�ٜ�#2A��\�Y%/����:��K&F �alI�/���faL�����91�'�_�����缨'����'yo�ڌ4G��f(�
Y�70����a���'SѲ�^�v�Y����U����k�U�	�d���]Yb[�r/�}��՚� �u�I�ٌ��c l����8��@CA�s�x��m!��g�v½{-���R�������cu�A��H!{�rI4��,+'�iU�~Ǿ�Q�S�~@�΁N@���v�Ð�#tM�g�_g�@���(�b��Sc���p�����ԋ5Gm��1������=�s��1�����n=��ks�=oKa,�P?�F2>k�0�pq:��z6���:ӏ���(ᑒ@�u�wA�ŕ@�eԋT ���/�ט��[j���,ވY�R�ţ�NJ|u?�Sxh��r�}L]��b?3_���U�O���Zx�)v��T��d�n��j�L�8���p�!�w�*��p������b�u��e�v{���?�ң �ϗ�~��]�li����Q,t>m~�WK�6�_��-S���*���5�{淪9�8:G���q*���Y��I
,��DYU��kF��@��,�g�Wkg�ƳTu�����܅'x��?��a�w��B�C@j��ߧw�=[Z�� ���d�k�!��~Pk���H6����F�0�=�>9��S��Kbv�Q�
��h2R����� 3���I�5�\����$��� w�9�9� ��A�L4Vf-���֍Z��
ȷ�!d�����$v�yԾ�_4�A��o��|�g������EX��H��M:�E�O>��ji�^]|9rl-�$L�¸>l4���Q^99M�T�
���;׈W�}M��⿧I��S��1�g}����T�飹qu ���Fj6�v�_��%]PÖ6")r7o:�^�D{�E�A����̘^5�o�p�<�8K�&mpl��d	
o|��J����ߟ���R�b3l��>�[�.���޾K�G�@%�''[<���$H�%�(O?|7bzAK��
\F�V[ �>��-Wd	9ܿiI>+h�ٍ����nuN#Ӱ�,-�5�/H71���9~oQ�����#����E��Jsĺ�-�(�%{���9���G���}#/�DiA0Ң�2�زn�@b����/�gE�t�A�<8Ci6:#q\�Z�59�(j'�����Ed��W����·��o �G(@V)�\�:;�f#p�q	�J#�d�޳֢�㒒g��p��"����`]�
X�k��_����s2-:"Gn���i%����_s�{�UJ�����Gm��8�u^�m�ؼrR$砉惣�1,�pʤ�hJP)=5��=@+Q�O��)�c['�����^���6E_�T���%y�_v��o#��bֲ��g�8e4R�Ǧ���0��`4R|RSEChm�����\C�)nu�s��6u
�D6?�3�C���kڌ����}�D�R=�!�ܶD	�cm��
�͇vK:6��nsK���t_a�~���B���!��4�t,���]g��Ѫ�v�ݲ���6�ٝ�H�2`��8%j�VF��aG�RM�l�q�IC!�Rh4�4��Uʟ�z��X��|��{nܩ��4�wX,5ǝ�M�|��t<��Nn����a�����)�mf�P̓p�.�\�%x��Y��D��^�Sk���C�5ӕ&�q�Y6p�w̒���u�am����_�6�������C�k����D�a1zkP:�D��D6:��ǚ�dŚ�yQYr{�ѷZZ��3�G�[ƁU�#+��n	�L�k��P`1�)<b�C,T���̙H�ײ�s-!��~X61k[x\�~���ȳad4k�|N��M J4A�)d��7�n�2���߱E��k�w������:(_l�`�,yW`nd���?��<������e���>��2�U =�U��l=�g[�iצ�|%`��A')}��u1?�N��ku��<E ��q�?���&)��.,.̡�(<Dn߅��Ĭ�3�~�m�EIyT�����	g|nf�gd��T��{��E9a����i���-�P�&Y�����!]S>��Mz#ggq����g�Z<�)ܑ��7�w�cQ��;��P���t.t��Q���Ӳ����e6�
��͜s�CBl��F��z���E����s�@�LM@��ִ�z�v�[�H�vڢ	��,gg[��P���]>r����hT�-��ᰃ�u����_�H{�|�w
^��1��=^F7��H�x�j����:��("��E��������XmZ��g�,�\8"�� ���rY2�OM��F�LW���E<g�慽��B�����ua�q���N�3�DC�8Y�n��e�x ����i����<��"����n@�pĦ�U��Q�]v�J##��uT���qYߺ�Z��Ԃ(��Xk{�<:d�����L.�vܟ�aE������C3w�8͎p��Km#\۪�5�a�ؽ5���d����?�m%\�|�FC�$�~�S0�R_`�Yɚ����bK��ʣy�1u��Pꔂ���L�`��� �i>��9-�W�hNkܹ$q�"ꤌ�����XBN��5�Vx�K�JH/zO�p%��	���g;�l��)N��hӘ��wbr�j��*Q.|3"8�:zػ�躙�a�Lu�:�H	�%�XC��ԅw9��{KG��)<`訡��ɑ2O�+о�<�dvY):|�x՚�&��(}�y�
�T�l�-3Z''��xZ�<�\��/�P[��x���\��o���E�Z������I�Y	���C՟��yVz�F����[O��:~�~�����3�k��ּA����RץV&��WZY	��l�Q�*0�7[Wb�{-�R�X�O@�XLtL�.	u#T�F���]d��Y;c���6�̤1NCJv���X�����v�ߵ:Bu�ۛ��;�ez��hTaGE���}VU���� ����4�a�`��yB���K8�������7�$<�!���� ��M�ȘL�~6Qk/�@M��ˇ$"E$�bB8�޾�j�� �d��dx���K|x�D9���A�5��q��q�}.�<2_K� ���+��Fq�1����TÄ�֚Di�6���Y3��p��p�=�D����(V7q^3ɻw��n@�(������L��G
c���Þ��y�����a����4�a���wʸi��y�㐉�
dn�e'��?����	XU����<��x�=��iC�W:Q����O�1��#���0N�ɾ Y�`�S���F�<�����[��/K��
��%�Q�E@�C��^޲��>����_l��޸�����7)�n��� Do�ߡޓ�r�BKK���cES{��J�I&1��,\XHA��.����c�z�������W�we���^�5ͮH�&�O��d����)���xz2Q�oz���4��[��Չ7m��T�G��4�c:_a>��-���̴d�)���o.�/շWҫSv���7��W��c�������[�m��zNű�<�z-�[��������b[~�Xt�n�V ����ӱ��Dsr���,�`�(
��qh�r�gfJh�Ȗh3Q�د�^^��`MV�(Ԏ^���N0��Qn?9�6� �p,�đ�r�n��fF�'ݶ-Lz�1�L����G3�����}_����8V���3�leS�����a��;ى�p�8S��\�������%�uH6=',f�g�_��|���mi��W�y�o���=��;AF4�����Ras��k�"�	%e��C����9����ӱ��	�I�l��=o���<"���~�8D��[��	e-�+��Šي�F>�؀c��t�	��S�+�ت�lW�w�¬9*3�.+���?v��6�T��o��E	�����}�o񑮁���+C�!�>`���z��|DX�Ɖ^��?��9�*0�f\+ ���{�{�тIh�E,'��dt���0M�����+��aO�!���U��R��^����E�f.ĝ��,(�V��p�E�m��,'�SG��$ܾd���G�V���.�Pȵ��_�`<�'I혃-��D=�hʐP_�N\/���U�	�dbW�8�-Q�gR��%"�	�LS`+�c�f D��<Sƚ�Uu���A�j"�8y<�z�"iw�i�4ܯ;���;��_��F1�!�ޡ]eov@�_q�n���w��Qj#��`4�1d��t��x�H�5����� ���S���" ���7p�w	c�� ��#X���6���B��q�,+�Z��L
�����?�'��4 �&�H[�\xiV6�qm�Gf�����Q��a��O՚ %L���/4Q� >m[��ͣɌ������==�|ߦ����� W�kH�����kI���R6�*@f��u�RLf�*���aF���B��^u��Ź��P�{K��҆���mNS��z D��g!�Z�������<�-?�'z�U��A���K�P�����N������z.?Zl� �
C�f��#����V��U�
�ӭ4 ������aq�җ�'�1�:� ��5�X�׀`A���XI���n��ythDm�gш	Q��z�$�sD�W��;$NI�H�-3wm�w�6��Ʉ��cmG ڟ�&lq<�>kZpvr����Q�z~D�����&������Y<N�BT���[Ʒ��D;������Ӣ��w[/ �z�B�i��@�����eZb��A�K���mv!<�9ǹ�x˟����7Y�Xۑyh��_�#maM@��q͝g� �\�k!X���SA(�fg��̑�J��]VV�Iv����P �0kw8"e!���t��X�xTQ�R0%���V���Ka,�oo�p@wvR���~H��e��rB��bf��*�`����%m��UJ�Y���x�[ĵ"��K
��SM���Y��Ih�,��Ċ��6�S(�
�5W-�"������9]�}��Y�Z��@s!���������V�H���`��3��֔v���pk�e��K�	��%-^l��k>�@�����g��?�{��MYg���Q��������BY���'Z��;$IA[�[D�e���`��jݓ� �t7�ɧ��}�au���1�k�!�4_��@���ͭ�9�
4�v�t�%-#�ϪV2P(�qOPO��,8�(�tj9�r�Z�ʻ�;xC�. �G:�Ǧ��/D�x��w/hs��ڿ1dD�;��V�
��l1�'Y�>�6�̟,H4���cG�ư�k�"�����]bIp���0)��B�B(J�MT;`�ӉCfj*4����WZr�#q������3͎=D*ь[����$x/�e����:��&�A���5I�zGi���|ʐ��%^�Ŗ�EQ���QR� 0_e�)+$���k�a��қS��It�o4n� �[Wv��sm���Ѫ.��w���gY$/+�ҋ
��k��(8�d�����]�p����d*-�#L?+�]A�ZhB{��תlc.�!wl"�2c�X����m* ��b���t�v���;�7r��wKv;����,[���:�_*n4��NF���5�Pz�9 [���v/�[^��EM����_�[��`���g�F����h�aay\�e84��-��!a�<ɥ���ȃ��̙��gw�P~�2��W�h���އ.Ʌ+�X��g ^�WP	��YN�}cU
�D$����Nc�$����r�-�y)l�S�:�F�13"m��3a�Ag}
�8\��O×f+U5?E*�~TJ(6���X�]�ag�V+�!��!� g;��O&��T�5=o���oD��m�t�ݝ(A�`�Pqo0�>��Y ��ķ���r��lA�����L�?Aܐ�[�e�M �=������X��k�>�;���L�M�7  h�s���P�ܤd=�	��
PޥX���c0����wW	�p̔�Z�@G�K��y+��,��D�Y3�N?�.~rM�`�콈6-Ϡ$U�6�~e(2y/7*`��3�3�{����W�qϿ O��}�������:Y��s�T�3%YKi�e�'�x������� c�� ���v�ƒl[�+�v��{�$M7��������O��5:����9�aU��y/~o�md_di����ǷY�q���3�J���s��'k���[�V�H\QO1�����2�`��@H�$W���}�=
u����
 �\{��DӴ���@UR��bg��3�d���Z��Cq,3��.�~Ev<���d�{c�b��*�2d��
��E���y����G��2'��Fkq������GIS����%�zy��3����T5C~��,��� a���U�!��≔��<���2� n�F;=���`��z(�K�(`?�s���K��4h��$�*<�\��p-~t:��Ǣ�K}3M�¦�����>�Wꙛ�@2��z
z-�P��4x!�8���ĭEBuD R0q�P\aDd1}�uN�¦'y�6w��U)�|Y􅒇'��}��x����Ӊb~��B�,ܰ��.:�/��c+W��)���^�25�{��5�WÓ��=B��TQWJsJd��f�ۃ��CMKR���&���eG�.ڤ�����%++t�M�i���:�ꀒi�y���5��ɻk�90jM9��;�K�0�uɡo�}����	����m�2��&N�e�Z�����!I��v�g��J�F�i�!�����u^t���K-�<��x�e�����Ϥ7q�p̌/RU+I�٪Oyol�\\�i�7���f��A�2ǺI�n�?Ğ��i}f�z�Y/?��|͑�:K���D�Xcꃮ-g�����X�QK)"�.��$E0щIU�q.��Ʋڝ�  ����@q%.<�&�Y��)u�T�5}-#N�K�F�-6i�n���qP-�_ߧR>�����~Π�X�������b=d���=�׎?\_1u�M�  �	[ma��&��J9Gs�JrW���B�5��5 Ԫ�|�1��(���o��7C$���CC)��6�0Y�𜤧���iU��V��ū}�]������d�Au��&�5�^b�&ڙ��sю��<�5�^]wO�/'�d��oX�ԟ�������,�V�)v� |��Z`+��9P�I^�N��i�a�hg�Ы�����i�X�qwBW��JJ\'Z�Bٴ��^��1\^h���b���K/4�#��x��� ":�Տ��=;�l�G8c�����h��I�花�%c������
$�'e�h��W�A|X>�τ��:���iH8�U�ު�!�9��Q�Èj���/�j�s1��ޑ�qcC��}l�U�1<�P��j��2�$�Qj����Osp���B�j�Ax3�3G/��u����À�&t�;f5<�w�Y��:�1��
�"Vd1k�&X ��z����X�
�*]��5oO��Ԧ�)�����r�ĝ�]����DW�O�����U��3q�I�X�-�:s��Ù<\�����`O`;Bm���M�rw+w�t�^F��1/�5�������'�w��M\�CH�7:'��!��ð�˛�Y�ח?��������&߲tơ�/��_���o��	߄��A�R��r�8+���W�.�߰Q���@����T��`�H6��Z`v@����=i�=�o':�W�Y+�|�&-�ͼ��L�0�~��������1�w���4�
2z��Us��t����s�q��8���_o�a7> e�/"����
�~@���f������Y;[5���,K��s�ia-!Yv�M1�����Gc#�����E��9�Ư˟�R�va�Q��xiwL;���/��lә~d�1�B�ֽte�I�U׆$$_�^�؁��q�yD[�֝���t��ú47]��,w$�Ρ
&�37��
��b�=� )S�8�$\%zr��T�$rN�A�
������:��#&�K8gm`�CS�~��$���9�k��!G��|
~�<;(�ì�
Ꙛ���j��~����hy����B�4|\A�Z������8��C��|��k�%�� M��t��Y[�%H�	�hh:�Խ�u�P|���� &��˒���CB.���ż�uZ��=��{��{AR��ţg<��Q
�sً
�H~X���Mh�`���}�>^Tu��i�)�3�̈�������F�t$���Ϣ�R"<����ʙ_R�g~�d$���Y����t!0����r`qFVo�F.�?|(�r|	�zR7^&���U��g��R왫�"��ȧt��gh$̆R	�v'�@�] j�ΩHI����Q������_�Æ'��7ֶ(�<`�|�i�9:A�GD�yKy���I=z�E�����B��J�6�[��Ҧܫ�.�:���T�����G��[e�me�P���~'{E����E��G_UZ/��$����3�ޜ=�N�.�&���T���� W�,�,���"�!�!G|��C��$ ��"p�̿��zg�9.��s��1d���'@�#���*U���i���F�� �N���G]�L�+�u��r>���,�l�oi7��C��8Jy�P	��<ڧ^|:32����B�sשjT�m��)�V��p܅U��t�1�5n���:�fz��l$�L��ro	����|���°������S������E�y�.�����@%����ʁ�8,͎�#!���@��>H�,�ذN����c�2@p� �_�����l��� ��Z�y����sh(țĳ7S��曢\9� �!˕J|)&U?���kb��;Q�.����	�dN�j~&g̩*�A�f������kTwuuC{�E� 6�n�2��]$*H����=��L���ge�u��q+)�o[��(��2��S×�q�#�VӴw�w�Z��EyB��<g|Q.�����_7��75X=.Ä�q�q6�C����@&�}���.3�&�;1Hނ����(v\�Z��p����D|I����ݠ8�<)���"����Jmy��}\˪8���ާ~�����}��
y_Z�y��{��2aȸ��>�Cy3�o����p8�E�V���gԾ�*QwN�a��S,�Sjt���Z�����S&����v9���yx)8'�w��������J��5SC�zw1���V;�ݜ6:�1���{���w����;�/b�%��������n�))[�2��=-�5@�����S.������Ǧ���]+�0C&���zsG���1a�&���բ�Ew!?�  �3��X& �?3�Xi{���Q����6kh���� �o%rK��O�QVϬH�����Ŀc@�� ��~��x�K9�UH�);
~5����>��?B�{�+�'����ρ��f�����xւ �����o�Ф���5F+��z1�ǥta��[k�;+�
t��2v��Q��9�����Ht6��.[�|@�dOY�й�a��4E�T��
 ���ؖ�7&���w��6����JּԊ�je������Oa�R�����	)B�{!T
ӷ��ʕ8Cm�o��Cn���L�ϜwR�@���� �ͯ�=.��y�K�1韠$�pABr�s
|��Ꮍ�Bb��Ɂ��Vq
tS�@��2j��Mщ`�t]ׂ�o��I�����
f�� |�9����婫(����h�U'��j�Xʭ<�����&l�u8��4
�m����/u�{D�0�4�eƌ�D��_��g��T$�w�*:ˬ��T�:nܧ2����o�r����nn�h+�'T#8���Ʃ�8�)��$�� 9�"�%ϖ��$NlNt�o�Dv�XH���!)Ij�^���y쿸\h}{L��ՙ��@J�vv\qj	��W1�B���D=�ɍt�q.��%�UL��,�7|i��"WSF�T>�ʛm�b^�E�e}��bt� �^��3���"Zz2�VT�wdR�l�nLw��������~�\�,����&�&!�G��Y��1�sSY���t��l�'"YFr6i����lo
ps^)LN���t��&�;@O_T�^�K�6l��-s�t�@�O��-E���JD�~=2�gK�Os�ன��ņ����]�P.���� LՃ�������s�G,Dv*�
\K��0�ց��w|6#[�ΧGn����ա/�ټ̩W�<�[�+� �?�V�{��=�@"k����~��+y�s F1�5��C=|��^f����e�4k��H���E,�>;�������w{B�J�Ս�|�u��-ä�G�^v��sޯ�Mz	�S۪��d������E.7r���z�F�k G�����[o���YĜy�)�B�h�0��B��a�ɗ:hO�z��PRL��� �k)�_�1F���-\/Z���ޭ�bD5�/�*�F+�ӱ�c^�!Q����ga��=}TuT,�F�v��a�Z)H6,����l�˹��f<p����#r(h��!~l�d��].$���ؔL���F:���8�c2m.{`��z����{�p;�p/Yj�=ѯ&H*�DZX�E4�&��q�݇6ѰA{3�M�� �̭Xd���̼�k����H#�\�wt	�3�=g�:���yC ���:��Th![&#?��Lgwɛ:�7��o��)�9'�i?K*8]�焹��=p�3��I��$�=�km�S�x��[��-��*jY�'?�W�����X�vVoG\�ޢ3�A���#���jz�|�����!,��R���� V�Uj<��y}�=?4�vwČ�?ɶ�u"�;?93殈vJ�Y�0����Du�#��pO��Ɵ�"kxv�y�n���&�uo>��81�=��G��X��Ʈ��|;������xe�$�@��J:я�%�Ԑu�d 
���a�<����u�{c�j��Y����Zp�=�'Jm���ll��R�\L�yYu$> |+��W_��y�c[��'P4�4+���`V������26so�*�+]JY�<�%���z�n�v�H3-�c�����k�-��$Q�^CL��O��4p���wސ&aO�b�����WRN�S\�+���*�ؕ/
�(�A��\=>�j�K�M�W��[L��g�s��1�Vu2����y���@H��I�j�����ONB���wJ!6%�E�;���Z����D�J�	�w|�A@�E����J�&m,�o"�7k�kA��v����JGQy]��'��k/(����xR�1zl���KOp<�w����Z�|}ۥÊ�j�vg�z����̘�(�E�#x��㠪���(�]��%��?�}.b�DUq6�w�:c9Rju�������+5����)!o!�w*�s

��,>�h*}��z�v}9.�W#7i
�N��VhJ̶u�"��,�BG
�Oy(�o�%r(Wd�%�9:���bzb�7!m��;S��Wl�P�4[��vyx�x�j�"\żSE~�B�w�������-���n��F�ޓ&2F���*a:���ˎ�(�YM���$��+N�O�'��0j�R������,��BC�R%���K`n�=؍+L�2d�W�bĪ��-'"��2����W�|��{��>}�?`Ӝ�pd��${&|-G�F9�z��-/�X�x�������Ʈ�|�V��ɾ������[��!�܄i�Ӿ���A!^9��y�j��m��m�ap�up����0JNV~x� ���e>���NM�4�sY3*��N�RF�����-���ר؟�K��[Jڂ���Z�D5GvE�q�z"�hI���ގ����me��sG�a �y�I��&��0�F��۸D��|���Z�h����:=�0z�(�h?�}��e|��0{��{�� ��NP���:���W�:��I0�N�<�"o���倁����q����ea���2��اU?RHR�J��;;,O�uÒ� ���P��;�E��c 7���ƚ���A�bB��e����ŗ:��m�.�g�'Gn6��g�]��;2�J�Z�Z��A�� /�:��/h1�{(:j��cI̥}d���\"L��A�l�u�}�xs�ߐ��G5qS��o*k=Z� LmYBS��I�"(������z��7m��ka-�ya|[�4���_y�8
�/�)?[іǜʛ�ix�kl� ��O�-%zvl;��O��-��c<��Ã7�(�K�/f�]����x�B�B���I�S|¥ɼ܇��uTZ{�U�o�Q�[�7Xz>
�N��=z����^[���G:�J�<�����#��2�ʓl����4�!�#��Sލ�S�dw��BH��D:g<a�i�oMDT��#�s}U��C�i��ho�E�\J�� �-t�(�H�u�+���+9�1S�`z��J|��14�V}>�e��	��I�m��~K��hj�ж�~���@�9e�+�¶Jb��3�`������a� �[w`3�N�yh�|X|�U�������.��P�eЮt{��O��~@_`B��6-�v��*�d}.J�-H4�N#K5��P��m�d��N�O��v�~Oܵ�P�OM0��ZƼ�#��Oԇ�e�(�
Ϲ��Z��)����R�i8b�_�Ț���JJ�m����ޅ��GCb�P�㣈�w���0R��(� 3�'��yA��AF^(�U+?Jq6����l�``�~#+��x����9��Z. f!t���	�tL��$O�*�:�2 ��t ��#S��nI�Gm:kW�D�1:��^$����c�c���k�D�$"@��1b�+�	��x�����V�~�Ƃ�E�D�w�9E$�jU�`+�Wv�J�d9~.T�o�{���u�Du��\e�찝�s��tj���C�Ͳ��(m�][`k�:�  ^��ʏ�Ir�p�,j��6x@��ԁ����A�A�ɨ��e��)�W�x�����%���|Ú�K[��'�oA�����˯���O �"��钔�ӑ���N���@O�%n�{�n� �ey,/�B�Jhӓ��Sc$HۊE������x-?�t�sF�+NȆk�GX����TŻ��$�be�a��S)|eǩ�&̯˛�.Ă^*6��<�L}(F�r��Pg�{gDP��vc�1橖"�v��7<���N^S?k�����pP��܃#ǈ5�]~4�E����Ǽ�t��ڰ��Q����������l����θ+�]^����)�F�!&:EhN�
�`Կ�M�mMd��!ޟ�~��zir/[V�?�
JeoӃD����P�U���.MIg@��!v�liI�o ���}�ZӺk��J�Y�C����~��\�{"�Q�
�9����㒢g�9T����<��o�gqBQ�3�����+�j����Pٺ�X�W��A܌E՗��p)�ѧdA`7%J�&֖Y�k&�ݱ��_�!k��mfR�B�oj
��h��/����������u�D���y������"��h�ԡ�	c�nN�@��`��'v.����	4m�t���x74{���+O7�"$K7]s�i��K
����55e���{>��TjH���ub����D�;O��r�B~c�aL䗡o1z�������e�
V�[#z��>�m�Y��6�3���7UE:��J�{�I�^�|k ��]��%S@SB��^Qh�FUP���|����F�S羇�K�� L��U7DL�rB�����X��7X���N��X�$�+��������̯�r�9�:@�q9Nql�����i���z��n�$-��*-�&D���N���ɗ�:��\7d.P�z�"�M1��=9A�>�|�'E�<�Q��:��6��o��U-�-DI#aL�^*L� ����� �=�'��)�����ۺ����H��T:o �*H�6̾m/�k3P*~�L-�c����ѢIǟ�$�ث�ӓ.h�p��cSё���_��WD+c��h��A�\%v�ź��'w���i@�i��}��-�bD�p���ZM�h�����X���B3Ql0t�y�6Vè�~��%w�Ci.��	Ob�kW\�j�-@�Y�!�����t��V���CfB��Yy5��Nedq�+�-1TvH��+�t]�Dս_z�6��y�K�T���1����o=��iO޵Q\W3u���4�{;��zٱ}=��Wf5[�Q�!+�Ǉ���ij)�U�8�����8љ�:�����-�a�?���45,�/_`���K6�%z����T?�L��5�j������OQM(�R֬���e�(?Q��J`�� I������K��Qʐs4y�V��_NFWm �E��w�F-��W���-�
 ]k��W�g*e��aھ;��j�cש����c��0߲ߙ����rU	���g�!~ީwU�k!�g��{j�=�j%U����?6#��9#�E�*^fC5PN�Z�/F�jj|������"��L;�9M�3����
����wZe���''���扣J �Y����y� =�:Z;�#_e��A��,�Ң��^A\T+9[�HR{"�Y�[Uu������읓�x�ړ��sa �p*6*�����ў���^u=]�楝��2��@?�Ar~}<��6N�L�oRS�� �M,��¤�rTJ#6�Ӥ/���gP�t�����eA�9*����	tJ۵l��2�����ȳ3�2z�4��y,�����,@������ �X�B��3L �V��� bwq�������t�p�c�;��H���n]rX��B�huQ�[�`�u���"�eDr���D�1�g�c2���e�0��_�"�Q���{��l��;v�k`�}��ø��
G�.?Mm6�%��f�W�y������Y��Z=[|�(WB��ײέ,��p3Z�p�ӌ��ֳ-Dx���)���|	��z+M�3�$98���#-��נ/?��=ߵS#�cY0��Œ�uٔ@<���p�7��O�&���Pfۙ�c�=t�%�	2�����ϸ�6=���u�a��O�i֌��@�L�mk$(q��Y�6��
u�:��0I��F2&��ډkkw5�¥X�!@��C�pr+p���{*'ðJ��_
�Ep���w~0N!߼�~�!^z	�AM�ve��#�8�����QBi�������u}v�c���W-�.+�_�J�S*�G����c{uy  <$����dgo��̨,��i�:y�ZE��*o�߻��y�E�v�ކ���N���c��BIJ�#&����m��A���aWn�{�Owlu�K88��O	RT��ٔ:g�\@ߟ:����2)�t6���th��K�)�w���sM����\�џ�@�p<d���[0��H#��k��0�Ɩ���f��(I�2��W{Bp�p.QK�l� ��$�jzDJP�;_���z�'���I��/c�3HHD�K�n<�a�� _s�����߽��ͳ*y����KZ�:�O��I-I�ȶw��Q;ِ�o���OgF0t�S.��@��X�a���Gg�>F�-�Y!�r��j6�<�Bf�0fVp�7���ָ��$q3d��s�}��,���vg�[rSb7J���'kx���U�:����ZR�q #@���fB�)ms�d�W}%e���'�,�E�r����R�Z�@���>�7~��B?Xρ�jM������w�}j��Q}�ZPk����.<��K`�F���ۑ��"���m��3b��n~������`V�Nz��n6�	TV	�8��g��Ծ�@v` ��6����N��R��ldP�'������>�^�R:k i'�.���9�g4�b�J�M#�^�m2��nb8���O灾)�����b��"���~���rS�}Ռ�@uޏEnzV�ٰo���1�0��6�/�D��9�JB�\�@�5&�Ǘ
6 E	G?��پ����Җ{�K_������+��w1I��R�)����:��E�>�\�N��j�*%�pzz8���pu��<��h���.��!�Y�f.��[��`���vNFF;�L���7$�f[F���౲V�O�&H�d}�i�񵜧XX�֡
o�0տ��q��.�jI�-қ�%�qBl��-��叻����s.���G����~�����U�dZ��S7rWY��]=g$_�/�!��6u��Fv)V���3��۟t�ٜ㣜���d*&p��f]U꣏S�E+�>"�x
x/]p�ULj��m��[K����$`��Z�]p��Q���1)�9R}��d�c�~٩���:��+Ll�Xi>�FO1Se��&?�_�a<����@�%{��ILI=�W��|������{�OjY<�-pIذ����K|��L3�uL^'�4?�$aњ<hkc��kE�ϦTH[�Wc��WZ��I�^�\��<���iF��Q���b8��&F�ϸ�#�R���)R�^��ɲj��\g��IP�)����ܽ�D�kT��3��+z��E�AP\>�
�:"�~e4�<X�p{�ZI�����o?C!�T��7�䞼JT���%Y�j:s���l�M��Y�w�U$R��ηݱ��6<�(f)��7�M7�s�n��с�)*f|
�<�ɄDD�U�ed��L�����f)���[�O��z�N�l��ǞbdlCw�{���,��ȗ@�0)�A�9]��D����09��Jn�o��+E�����X�x���~q�FLNi�K`=)[��[<n�����\�%�7+Ⲩ@�����I|B���kD5� �d�ݪ���,&�y����ݗV�|�5�g���u]Nnˬ�QaL׳%)j�J�/Q
CT���c���v�D7��A�|��� �S����T+s�^�❫k	!�N���y	3���B���WՌ���øFHIw�����n�5϶y�,�ʰ$�d�1�3�H�䰧:J_|��q�f*�V*�PO�J.i����_h}l��ي�m�Ϻ��֨��8rۅ�p$%�G��=���X���AS����N�m���7�;�ůE�v9�I/���Q�Ɩ�y�D��ջĈM��3������s��ྸE��i�|pAgG�a���H�e�<0��I��Sud��I��/b�-7��?dR���2����D+��\�c�S
}wD�����3�q�M8|��;l�w��Rה�luD�q]��?����}v��0<���z��������g��V!۵}�8i.�[��� ���١��Dg\�8:��;y����ᷥ|2�+�k�?>1G 0^Cu�?+�%�+֙��4���;�jp��r��JD�Ԣ�7C�e֋�vY}�g� �9�l����5���y� #OEe�(Ђ?p���3�&�Z`/ve��<��!7H�M��t���6���\Uh�w5��� �nW"���.�Ka�y�JB2DR|e4��qJ��m4|cr�&㋹L��������Gj�cv}('�Y���G��Y��:�#@SlJ�y�5�he��g��gsh*��7�;y��X�.c���#�n ^�R�p0 AF	�S8��s0��\�]�-�<X��ʧ����}eV{|>�s�E�;�l=��+���F|���}V�=���F�?k��6�C��[;Pt�뽟�%.���Kއp,�HX����j��(;3�Ч,�]"����8�U�[��ڄLf`R¥�˦`Ҵ�����w�X���}2U��� �a�,	�jzy5��>���f�3	h3ZN��ۏ��Vr��R�.�%Er��&�/d��"��|���ӟ`��R>2����-x�ó �U9���G��fs=����>\��6�ל��v�G�v�i��d������T�;�]卯�ϡ��H���%��LS}����r����HD�M��E"�K�M�#rB����M���2��jS�R@�NǠ���s�����R��Q�;��i5�#A<��>��X�C~�D��X5�&m��-, �F&�6x�zb�"�:�Ȼ�I�]�z<aQ�Ӊ�����'I��q�%���ѝw6d��l��q�;�h�g�9�k��u�`׷�r �R�ݳM�mkj�H����oMe���+�Wx��.�t����gcX�]��m��E�l\_�٨_Nݚ�A�Ǣ�8_��v�hri�:w���8��%,��� ��6(��:��lhq������@C�� �%�6'�I��m�w��~�/8�d ������ܼ:�"�{R���9��{՛�u?&��7��*>_�"�O2����7I��m:�������C���w9��O@���Œ��rړe۵�|�� ��h�`�l���!&�>�~��PtWig�]�~o���9 ���x��%�P�S���<>����7����K?�C�YNB�ԙh�u��APRS�����f[ۢ�_�u��?��b�aF���Y����B�F�M�^!9�y]Θ�"��b�(؃�>�umXr�i�p�.�D]E�S��*��~��$�Z�g[��M��\h7?22&2�Tùu����\:����2_昶�:�!V���^�}����"_.2.&*Z`MCi5K���`�������qƖ�'������y�8�e}!Zw�\R�K}Rf#��m��b�& |P�k �1��&1֌7N\��j��Ws}� &��fi,�q�Ye%d�6G6~c��u"�����A>h��c��ND�t�����+<���N�to�D|�L���B�s.ԡR��P.ь��lf�o�$��6H�����^)�.Nt�`�@��*��'9��k�wZ?��:��p����1$�93�wI�T��^���͔/��ָ8Q;psZ�XT�!3���l�ʨ�������#�S�O��M ��Z��ՀP�e��MT�*Z�c�߹�����.�����ѡ���,��.��mS��v<��=)��]/J�-��vz,��81�I�Q�i�Z������V���x�?E�؝I3�d�d
�ß������^��*�k�U�u��9F�u�
t���D�gW�v-�1��gP�=qE���"�u1cK|����]sc�K�m���\�J�
#Ne!�|j2!�gH����u�9��;�d�BM�W~
2�(/�hriqI'� �dƃX�ꌝ�BZ������g�v�����X��?�q;�b+kN��gV��Vܹ�!&�C t�i����裢��3'Ěq���}P��3���ۃ�zI�Z��4{8�5��	�&���rՒ�����G�3~�-DzX&Q�d����C.��T�"���LQ���H�2�9���f�/�M���1r&l�����k�<����̣�;�5�콨M��R�0�����u�WpQ1�2M��C%l�B����>�.9$?�].X_��T�b$�	�u��:����Vw��7bR�E���L|
�k6]Pe\��4�odյ#����2�~�v7[3ML��Z�i�n���"�~7#���S�$G ���VA�7�\(����7̃g:��z��/0ZĎ4Y�ub+Z�>\y��wy"�(`/��Ô����h��q�!���v{i;�\�����u�����7��-U�0QT���Y6�����mm��y�$%hh&�*E\b��rve�ό�%T�K�75�aNqOe�������~�՚��� ����̀f��Sh={��s�*��k�ܑ�W�<͗����d
����~r��}����򹔤5o��G� �>%��BV� +C��Hp�����V���^�l�5�;-f
H +r��?:»(T߀N�!�ۊ�u��̐�4�� ��76چ�rt��Y�'�����.���X�P�3�+��*ob�|X�I_�K��g�M\͹��S���=��q���Uּf����{b�*H���0W��K�'~Ƕ?@1`��Q��!�
�㻥n1�W�>X~���u��7�`��B��'���x�����������7��w�b����-����q��[`;t
].:ڟo�I^A��ļ;�9�-?vk�"��A|����D��Omt>��I�T4|��wU2��&��5�?���	�I_O
!�Oŷ�֍����-��
k
��p�	t7_[b+�4m 	��~n���s�����I��.��ׅ��@��]�̌gkyH�] F�?79B^��F	��Ab��\3�����+����>6@��{�]n�1x�>r�ڹq�e��ܺ��b֘T�Xv� ��~�`|�R����Uj�U�'=�kf	���;�~^'����-K�q<��r�l�5U��$5-�1v�YY+P�ug]�݌��H�dU�
�����(WU:[��Fٳ.��a`m5��\q��?S����̔�Y�䜙g��_�	�S�i��'9��/X��D�L������N�ܓ
f�sE;����y�\xc��0��8�n��J����n�iM�a�䠥7�2U�0�`@�Û�0��F/�w"f�����������&�w��� �r�"p�+���x5yg�\3�  a���k6�%Z��X����Vx@�����%~+,�?�;�a���{��L�&aZz'�38έ���M��=Z}@ƕ"z>Ǡ��K�h�J�( 5�j4+�n7j,]�X�?��R����TF
?�Fw�'��g�:�(h��:B�ͽ
(�;A��ZQ��F_����h*��r߲�0��Af6isUn��b�N���&�����4&��獄�O̙סA�U�>��y^��/��Ý�O�)v�pR�����2��ڦ��6��T�ԩҦ{�2��P).x�m@O�����ću���dv�?]!����~�3;.@ ��=$|,C�Z��ˑAUא9FPj�5�Y���d�m��M��"�8��?����%��Y����*��r���߆/��q�"�}^���R	Q�A�xY]u8����)C��&�$N�*_^+��g�_-\��'���G��.�f�8Grp'2�Ex@�_��X�nmw7�gR���P9����!=oDa��fS�A�#��$�a:���H�v\��&�?E�b�ltl��$*�a�4h�����R#y��֑��3TM��OW�6A?x��h��ߧ���7�}9)g?�$�8�"D	�|����-��7U�S��h9��c�|hv\�p|(M��b��K�4�*��ꁻ{��	�*.'��*�Y[�	���8��c
�{T}g���O�����rn3Ǘ�ո{��VBb��°2��<���q� ~c�>\��Ou�s�?�C�[��<�M˙�<y�'j9�m�F�=��Y0��CFkh-�?����)+|�p2�{.�ﱁb���R$�z}#�s1���'�v�&��%��	uuj��i��A9�n�oB��nHۀ~�����2	�btRFy�Mĵ1�\���v|��'��Y 
�N�����q�˿�@``^���;�g����|�$�]1�����]۹���Q��6lYtP#@ lT��ev�ɶz�^��K�:#�GhG����N
yi]s�܀L&�Ĭ{&����B!�߾�%4K
2�l
_z��U��-�i�
����c9�+������R�4n���{@Io��(�ZY��}]J�~��5��T ��J�y�xe���Q/�,s=L�����úz�c�D��X�߲o3����C.7������A�|h޾������G_E�%�Q�(��UR�O��z,l*	���_�|�N�d�C���0y�r��lr�&�� _�d���p�����~#>T����7��6�o R��N�]b���w����]�4��d8��V�ض����.�r.��+�柵�{��+m��b�s;w���S����5�Tu���@�Yz�r��͢�wn?�&2�W�n�p��Y�=�|�K&�E�"^_���BU��V�n���.�@Q�+��I�Kp��ث�݁�A��ί�>Κ&�i`i�tv��F2�����<T�X2{p%�dT��8Ֆ�tfߜT��*2��A��r�[׬1Y�-�m�S�s����G��&l��%��&|=�s�UVJ������c%@����2��;[9�9s-"!��}����ɗi7��ӛP�zXD�)��l�ol��y��D5��c�zp�_mE�i�7�,�^��������N2��o��`�WY�@��d�z�A�a��tFr�q�!`18sؠ��f$��[�j@V�\o`p��b��{gq2&3^e��}�Ѻ��'�hNAtIo,űyz��;�3�5��6�� xR�ZO�B���iѭ��m��,�͟|�%9�_�	���۰�n/�� ��F�!(sn����A�?0��9=tM2e��8_55<ɬ//�MV�q(D+��!�"\����K�Y��2V�;�Sx�+ʓ9ظ6gLL �n����F�뱗�2�SRd�ő�gB�Ķ��'|��x�Δ��ACWh ��o<M��vwl�e�^�
v�-�T�\2AŞ��=)��uã�oG��u;&�%n(H���p/�p@�W(̥N�1h�Y�ѿ��2P]bv�8��5������GU�f#�(wm�|]DJO����� ܽ]�<�j�U�ƶ.�9�v�|�b&�$�et�#����/��yT�J����$;�������C��Zd �>X���b�l�ը�e�J�^XP���Y-�0��kw�;���d`P'�� ���$�IA���Y�.T��箾`7#S���`Pɸ
݀$���u�i�J?�tz�3j�:�w���S�q��i�|9׽(��d�1������"�a��-+B�>���I���l�B"`�𹉮B9i�����+�8�� �k��*
nI�Ù�,� ��	��\��E�N�z|�Uh�O�x@k���zf��+��5߇�#�L��W�j�><����[�+�B
:1�d�:b7�&�. ��h���>[c��-���۞�^J�+,��{'*��PaJ�>꼯^dL֌�2�?�������0�x�J�:\�"w�-f!����Y"tQ�y�r��g��!xj�7dͮ���;"wޒg�Oɦ2Y�z�hR�j�Y�ڙ�m��s��$s��s�> �6Ĭ��N7�v�^%f�m�9 �Gdp�)�,��L"V
X�d��Q�%� ?�r�j�XO�Ʋ�,������ּ�������H�׾���s��3M]��"�ZĚ_�����T.����Oi�$E�R����]fQ<xz.V=�<K�ջSk����ݙ��a��j��t�l���?��-�Z ��2m��t��e��Ǉ�U��⦨l�B�M��hom�^�5�"<4+����7�܈�_���Nv �/�O��UzhBV&�O�չ�95�~�#�k�GҎ#������*߿j��<��t��❟��8�!��a_$16$�������K�g�>�y����ہR���I{`�}���0�:��X���ߴ�ӫ�����q�m-�d��{��n%E;�;��O?�T�����Q����`���Ӈ��żƱm'�!@J�&���)���#�?�^���[�F嬸���/9���Z��'��,Pbo@�ӤS�\��oY%��k���u�}�L6�n8���g�g�v��}X\T8'2.�����=L ��ҍg ��k1'z/Ǆ�5�A�}����Ԁ��}�ef���qH�/�4u�g�ŉ?�ξ�������)V$.�1BH���S��.�����~���mI(_`q؆�9bژbN�1+n�I���	�5�LBܿț�����Ԁ�:.�5��n�rH�\=
k�I��gY��#�^��~V+�WLفz>��o������!҅mK}1_�c�j�z6�z��wi$�;�7�V�J�upQ���T�?}����*���Bx>�b߫�+�C<�
?X2��#��R��_k�Z!�%c)�d�i5�s�s+ǂ�?��4-=���$����j6��&�Kn���K?J��:_Ӏ��cNB�'��Q���|�zé/�/��������	/}֐8��k��g"$�d����<-1j�@��"F�4�C�y2e�����6ҋ>��s/eB�v�	b�VԐ'p'�_��6c���g4��LW�<��96�{��e�g��4�d�*��5@VR��`s��=�IU�1-�\�n^[�������m���
l�{�׈��vں>��.��Yք��G8H.l8�H��6y�=���{��H)6�V<2'֪<�{ݢr~�� �5޸�QA��"������R�	)d*<���AVVd0��޾�"yy��_��A���;0�TTXz���Ơ�!Ɣ[XЭImJ21`F��f���>P��Q�M����r�6kL>=*��̒�I�uΎ ���~�,��xR�� �D?5��5���@s���gM��)獪&:��R �ṵ��iֶu�X���d���)�j��P%jx{�9���q���&7"8�*$&�"�y�B��� 6����w�X�Rb�@lڢ���Yr���]��Eӛ���_���>l!
Xݦ�w�Db��}�dг��=Vjӌ2�)�j�H�[�`:8bϗ���+�	�0�(��y%�"M��O�`uY�^6x�j�̾m�\Q�߻���V�q����R���w��u���;P�A���(.�\�2�X�I=a�$��=��u`��d%��$���2������D1|/�� �N/��UjJ=᰻F!�!�߇��{�Ѿ5Ƹ�47�2v���?���xf�5�-�~�R[&eNn�hHȈ7��m/�@_�d�4�ڥ}��_'�f�J���P�5��	�����pf�H �l��콪��м��B��E��D��P��N�VO�]�x�!ŌQ'�u�g9��	�M9?������39�R:w��a_�OL0g c6�9���;��ޜ�="�6�C�?��!0O��`V�q�w�����ȃ��H�ϣ�(�kfN�>�ُ8�k��)�h�K*î��8"�$[�r�^�_�EU䬹�c��4G�t9�m۩��c3��k�����5�"�q_MZaf�+�tdev�)19L~�8��0�x�Y�ꎨg��ɤZ�ރ��xC����R9
��4�+���~�=�/`j�-Kp��v��BoЖ�sP�ՠ�k	��~|�9�?I$�9Aji�-��q�=+�ڸ{p��J�5c4-`]�^����(�p]<<������}�1��k����.�5�,���&��`8�L��J��E�� ���X:�������J;V��Ka�nJ�Y��+J+->�	zڵ&�JH���2��pͲ�MU����0���M*����,�YNۡѦ���	7�l9-u?7鷳���.(:ČN	�k%S;6˻a�r7&:Xu�D����(#S}��C� ���N:�+pVq\�gw�B�G�_i\��G����,'��J!!B�b�w,����vs���ORr����bЊ�y�YNjpؑ�7XjŘ�)E�{TͱD"��j�H�*^����7$���Zj����	�g����(���:����Hi�R����������6�o?���YrǗ.���jn�&�iX�3�����)���3	~�&}^-�RD�t���vGFz�	CX�i8�K]P�8��#�J���ڌ���3�4��i�(=�����c�v��g�Ç¼'�1_��5�Xd�fhn��2��K��_�&�3S�v$����`�}b+���7`�Es7��p����gDs���{J��-6�O�&;��׀�:����� J�xK��l�jާK!�|E��zn"&��������Ikƭ���Y�<�_ec!ʚ=T�]{�M�l�Y�J�k��/������ѕw�y�a�ћ��z����g��IQ�:x��0�)��um�Ց%�な��ѕ�Yݓ�|b"-��ڧ�۬��C4A�*��x��#�vN)�m�Tb����q�C���	跖�H�
޹q���`�4�.��B�i2~��m��そ��E��]g�U ��i��h@zV�W�����R��)+���숺��Fͺ���
3�T����u_��{���??=��۶�H8=%6?J��O7��r�����&����L��4�> ܆v�L۴R#&�H�2����Nw<_:���݊�R�0��.���Nuo�ps�2B<� ��bc7�=��V��`�t��AE�C�I� �XGq0l������Z&4�I�Fz'�%�*�3̓��L��@���$��w���2-d�(���V�GG��v�͘n�C`�0O*�:���`�s
���6@������O�Y�W0�����Cۉ2.A�0O�<�S�3����v��K�W���C�467~�H�\9 �]��`�~����i�{�+��r�d�+6�v���^��K�F[�dx�I�5'p~�!�, ��x)$�����z1Ǌ!޾>�H&K�7����I����\�\&�9DȲ�D*krs���5���C�g����Yw/�y�s���h�'��ڧ,�9-���jq��p��Q&S�<��F��b-z�]�^t�*�\����evZ�q�j�x=<�	���g[��+X��%�J�,HT���t3��[Ѣ("`I��n��V��'>Q��(�z��Т�	Q_�|���!�O8�K����O���&3+)3l��ė	�>�"�v	|靭V1��T�N�9���LT��X�E�M�4�ӹ��i%%��K��)MZ�'^5�{��6��Q�� ���	�c��x\%m�:��� .@Ĵ���l`EX�;KA5�vmL.�?-�$&w�cez\ڢ��K��@�Q��R���j�5��&�A3B�������XIR:�� �0\���w-�&Tc��jo���[�����I��>�0�cu��f'�B�Z9Dy���(��]��y�l��a�u�,Y���ug'���o���*�T!��xؚ� �\���R���*�`���h�5��P�e� 42-�����g"�pܶ�b[��"6��Y�/'���Ǟ�O}sb�w-��_3�<��W�ǂ�4}�gL�"��5$e�� ��xQQh<��z:<S�<�2��RJ��:�'3���3,�h��uP���J;���F�N_|�WمCW�otw.���"�dy�R_c��A����~����q�8wJ�kLF�Ɍ�����x|5%���ɢ ΁�{'g��s��5����q"�!?��v����0�c��?�x��ΝL�䊚��*	+"���Ӵy�9�kF�mb�O$	�_װH�¬�oxT������9��h�����E9�r�� �J�Z���1�X����.�,�U������B�2A����/1K�*�y�>���[���x�|p[��pJ:jd��ѠW" m�Nf[7z-�A��	��t��6�5�
��`q�TPQ�ľ;�]$ P�<'i~�1qe��b$�3�#�"�1��=�Lm�����o9�&'�N�W䑓PM�����%��rL`�KSwS�J��M���/��,\�d�&v�&���w���U�F�8�$�g��3񰘅l����$�f���.�Ʀ�Ed������|��
L� $9��⌇V���R��{І��r�`ʙ.�����9&��jA�o6���MS7�S���o�3�ѾJU ��X��� �-���3)>m/��E� �ʞ�̄?[�{W�x0�T&�J�(6���Z�:���Hg�zCV��s���U��㑟���+g��7�(� (L�Tz����j�$p�������f?W[�w��%��_��<%>�+Oxi$-J߮]�����s��9� y�R�R8.��)�l*��cMm!�����r�����驆'H�V��tȹ�fC��`t�;�x/d6K��Y`�}}�X5���i��-G=qT������n��qS��@�Ν�r?��M���@��_X��>������S��
]���4�!����:b����8ჲ����ʦ���N!�"1,�6i&2�����ҵh���	�;�@����zRG@ԕ�9yBo��
��gdk�:i;R�%����eԵ��l�<ï��iY�ͽ��m�,g�keBC��}4,�h8b�ָS����9�"ؘK7����L�: �X"nl����k�$0�)�z%�<�,�T܀F��(����1dي1�kq	d�ۆ���ɏ/H&�|�~��
j�PB����;K~_0�g�G��0r���R�}��{Ix��Q��Z���7L��׹��Y}be��X�F�s}�7���%˔���!�up�:J���d :���k�5��b���s�C?��p�)e��̄T�{v�C�Y�V��:���	^O��[�����{�Q���TC��?]��yۨ4%Yf�n�D���Qz��(�;�(.y�S���υ�1�����*Y+WM9�� !C�gJ���˼_��-����"�#qm*ᄫ��N=��O+D7��o�W���R���y��ڭΝx!8
y,���}	{Jd$�B-�Ӆ�ଣC�^�z�Hʹ�3�Գ���lG���3.�R�ަ/�e��g�jtR�MMKa|�(��(��v?�'�%��b�a�P��#h�Y�N+�(:�r�T-l����ɩ�� HH�ڐ��.��'(�ib:��N�-Lw�9�����0�Лh ���l��.�+�[�S������/��������a�[(zB^[�D�ٿsOPH�Sҟ����Zav����C\F�����<ւ�xilÍ�/�f�� �VU�d�`S6�e�p[ώ�H5v'������u{W_���)[�,�ގt"��v��k�=���%6t�cv���i�^�~ImG�HX��a����ڞ��>�d�DRv���-�,�zAw���+��B� X�5�Ʀm#Q�Ŏ-*�Y���¦�lN��F���C^��H�+��'�\;�$�EÑ_?�#y�u(��q��^8�q��*���*%-������8�بJ����V��:)y�����N#ʻGF��H�ާaU0e2Jݖ7�F,7߇B�1w��N���Bx~�p6������_	t�@��4Ǭ�;53$�@x1�r�S��O�e�N����w�B���f���E�?S�f?�D�r<�����D�����)��u�!Ʉ�yj��n׭=��ѵ�wÉU�W�� �v����p�"q$����f.E�J+�QBk+����VɎC�����l{b�io�T��ޟO��&�Y*}����+�X�0�!?��9K�5;�}�j�-���{9߾�i[�|�ٮ�*;��x^����S��Z�9r�#���_���'j�����5�2�#�M*}��6�Sp���/k,)����ƣ�zĉ��qD"�#Q_�)����*wF�!�ߤ�PM��f�Y�{:bП����|cB�ԗ#�g21�^�u~b7��،D ��d��R�\�΢��
����c�>��>��Q�����,�,! 5_�sQ�Su��K�Q�D��Aω��b!/��/6$6WqN�1�����3� \�6���c��8�ٛ�z�-�B:u�3搢�&p���~߀��hDۻ�T�߭l6��Ji�]��gd���A��g��舻/�L�Z۲8�´��g�z���&�Ba��Y�i�����\K&�f�m�<���k9ʰECf�G%�l��fTk�L<*T��(���2���׿	�r��	��H�*O��֍����}�xG�p;*Q�w��ˤB��W�?�J���b]�37�\ �jq�>�pA�,��0���t�)�l�gQ��ۛ��RE��l^���*t����D`��e�� G��$�Cs�N��VrH]V}��&8S���m0Z.���~�gKr���(�qa����Q/��1sJ��I��� �k���XdJ��4!&)��l���+c�7Ζ� @Vh
�ɭ%ș�٨������A7iX�ai,�` ��=�9io��^`]ߥKALq�#Q��3�����j�0���gd[c,�K�����בE3:�O�}��YT1I/�'P�<�ᇠ7�_�����F�掆[���eG�w�_}B	JKPߛ��+�DK���{ω�6��q�:���V���)O�� �	��.���H�[��b���[��Ԓ]�V&�J(]Z[g�I�҉^��P9��e]6C�2��E�%�ᦠ1��[|��v�@ꘗ��
�>��2�χl`�:�X��S
X�1XnImV�9sk��v|�@;^&n����&����mc���W;�W~���<�k$%p/yC��\.����i�}�����Sx������K�l��:�d�"́��[8��w��z~�t�5\F#{�pz!nѤo-�nױ�����|�� l���^������m�E2���ky;]��
�%~�!/R�����\[�`�O��#5`JH8�lk���|���*�e%ݺC�5�G��gQ��
�U��`8�F��0R2J�-j���%�Hcc��1��(�a�~Je7��\������?a[@_�S<�`�7���<NxC��:4���(��hT��w'�Xu&i�R���)�g�Jȓ9��Ah�(V���b�v�������)u�9ߵ"����aG9��&J\��w��i$��sH��d�Ѹ?|RGy^O5�ղ�#ݎ��U��t8ی�������T�@��l�;��X0���/
�O�]!)v�p�4����趐�md�_a���C�[O�Σ�6�E��AZ@�r"��Mt&˞E�t�?*\�^��5���VM�z�v�t��~;$w�������7ɧ�������q&

be�IbK��{fa�����*㞶�^��2M�=��}Q���1T�%3ML�=�U?fl�2���܏������5�8����R���,������b3LF)�r��,L�{�ؾ�&?�{��y3!Z4m.�=9r���B{N���IXRt��3��l��i���|56޴�}�W*�>��G?�� #�@�\�,x�蟜�(>�H8�-
}]-|�������1���?f���� m��&�ATŕ���O,S�9�ݛO����#c�Rݟ_�js�-�7G_e����!¾�%��@���*���7��x���h>�F�<�Y�N;H�̹���$x�SR"��$�(w���N���>]��0Ɋ;�Si�j [�W2_���<�����Tn�X�'5�A[lbv��{��;�t���|	"8�-�����`�z�/�V2���UQV�5�Q�
�:��N�p���ò�v".�=���U_�� s�o�k��i6�#��*�2-�~�f���$�a*Lr�n*ω}\FE�a[�:)Ā�6����4�x��	�(�P�2���~hs"�,Q�}>$&��.�b�܃�?���"�#
#$W��_D6$���/��7�r���!�`�d����334�H,�@��ꐃ#���y���V�VRo�(T�a�x�e�4c��	e�4���U�����k�)�44|f�g��M�*���(鹝��M�9��>Ӣ&����%��#��a�|����+7�a���$ρ;��rT�I���SƀצU��s$����nU1�E�X p��P����%H!h�|�&mI�CzH�yu�t8w0��L����x�h	q$��l�a-vi������
���Dk]�����?��K'�eE�9ήh��P�� >��۪9����"�Z�i��?��-��e������ǟi��������`�HL�X�h����n�"B����쏧<�5����lF��+h�{��m/����"���/����3�Wf�D����e�%� ��]:	�cDZ}&�^��)��6>	���U�Y�����U�?ºT5i<��`=��!��hs��q_N�uj�.	%�!@�Zi��5��s����m�d���i)�vm��,2ٝ���$�u��nL��o�G*<>�3������&��|˄��Z�P�����@��¿�s�\*�5{P��瀳l\e���i6�j�w�ڨ��ÁG����|eR&�vo��3n��Zr��1���u�D��֕�]Pe���˛�,���!J9�g�jtv�o%�-�';$?	۷����95��x>!![��9b�rV�Ƨ E�?P����R}�F��d݃���	= @� ����h,�<hv��E��J��k��iKe� ��ˋ}/�?�3���N���/5n#8J����?�»���Ӯ􀵆��;���=�Ry�5")�'V� 4b�s��~��A����r���[�W��js���+a���� �1#,��>����۷�lUg�_%K����F��U��wv�y	J�x�Y?�9d3�5�D�����ۼS�E�1
�v2N�>�ݻ�j�]5�]8 ;5��r8(�W�ܥ?��d�b�B��T��mp�}�Ho�^�Hk��q�$zȘ�=7�o�������<�~��������N�u+\�g��4��Hw�/:�1��E�3]��Y��A=:|q��<EStR| uJܤv%���*5�WG�&��6KSlE7���9��G�e�6x��_7Q�a��$/l:�I�O,ۡ�0R��}$��+"'nۭ�% ��#�ᬿ�@�m�	�D��AFuT��	�W2Sl�̪�EN��~/=2	GR<��֝wB뽱�e�\��I �h�7e����:��͏,)��E��E�
�Xq��)e��KarX���;�a(2��J�R\��9\�x���;���ˊ��Ȥ����It�x�ݙ�"�srO6��M8/D�K	����4v'e���@�:�8w�gk�[���D����WW�����/��5��c��	E��\�1gQv���㚞�v�?��]���C����>����Ao*#J
v�l�ɾ��p�����o/6�E���;|L���n�O�wy�m��>W�1�������}��=�F60xx��CT43��R���p.��Oۈ�4Q�e�\>�������c�1z���b�8�S���{��PE$�����O|Qx���]ɜ1m*xw�6��~c�0��򬯼U?s�7ZzmxA��Vwk��X�ӃQ�.ls�r�ё�r�Ap�"A�Q�<=+l��r�|�q a�h�<g���GU������ ���� �u��2╂�f�Vm�����o�_�H�r�as��}w$--�V ������^#�o(;����؜�Fy\�oS��J�kS�5	'<�c�V����@�d��kI�	o���ܲ���] ��}Ւ�;����nh���W�Z_K�2���p�ES��8Sa�v>���Ɂ�RPm��L�7���5���]��J�+`�ԄV!���������f2�eM�~�p6���j'����Q����-�;�_8`b�E^�U��#1���s/�I�2�����Oæ�
����/[^��*������Zܹ h\�$R�K	^\v
lrK�~"�����2e:pq��,H]8�g�N����ņ7������u��E�8}fB[1��_�MI�>l9~�>W��C{��3F]4�I�'��	�����Eb5�^��{���P�p��m"����-�vo]�DL�y��>9�;�aO�.}	����x���72������CEګ�5�a�Y��	�dPR�N8"ds��݀K^6c<u��Ě���o�����?�F��=@��{�� �y��c�?����
A��-�e���`*U��O��p���wgZ#Nt�)�U[/�(���5���\�ZV�+7��y��LD\Oݷ�������QUu�)����5����2#,u�6�D��siV4���LL��1'6
?�s���ː�s��	}�W.G��N{���e?ڋ�6폐҆�M��b� �L��b�7>t"3Xǰ�.�M #�ey~�y�8
d۔���
����9�RW��4J��縊z�
Q���[���J�[��v�|x1�r#.)(�ʼ>�C]�r/_m��$	�d����Sg�vK�r/Y��.�"��z���3���%S����<�\��U�#Ĉ5�"�S�"�w��H�n�~�©�o��;��х��d�J:b(U���
w�%G�0lVS7r_=���`9N/�q;0��o�I�!
wھ�O�� a~ S��$&�q�n?6�#����Gk4EW�lT��+c�M\�{�?hj/����A�a�����ag�ԇS*��}�|,�燶��L���'��WL���1S3�\��>�Цy4�P�ɥC�67W�1������M�Q֩�L}��|�i8�)3+�{SoS�O�H�j�#d��wtt�S#�[[yb�����؂����aD5w����#�vj��&�q6{���7�0���=�]����k�[���VMO :�)��8���0DtF���;D��6��Pv�K��T
fte����΀�}�������p� �qx�ըy�^������p�K�l�븘�ň����K�7K?Z\pB�u�T�&�����	���(C�_g\%��L%U�wlz�͏Լnk�K_h�i)�����E���' �X���������W��2^�9p���o2>����J�����\3����SR.�(|��e�KQ�7�����W"���r{H��AF�;��p-�I�U�nR�-���e=�#�K��(\�g�ϛ ^>bi���.1gp!s3��5�Y��Z���0���ӂ��iI*AH[��1C44�r'�N�Qe+�[T˯�p�h�`�_��Lk��8 ���iԃ���@q�6�ƕ Ί�?W��m����\�dm�^R�=��T���Y8�<��G�����e�ڪ�	mA� �F�(�פO�J���<{��9ѳ����Ͳ�[O����|.�qZ�`T7kEtK�|�6;IS�]q��r�DA&T�@���������s:#�����ϔ�|�麡 �\+qh���7-e%Z9Κ�-�ڟ|�����Y�%��_JBc���~s% @�����#�e���g�-� ���>����j���u5��R��^i��B.���O�d��>/Gؿ r���&;V���r^�_*}e�A3�.�Y��Υ͒w�W0&�'�n�������l��=� �s��{���o˕;s;�����/�������4 
۠3���,e��{1��hNTʊ�9?�D�GMO�����z0	��t��߳�t�����
k��{���tQ�^Oҷ��%��9�F���(\�~�같�%\�ۀ�Lw��x�>uK����D�K�lb�H���´Y��3�G`g޺�Ym
�LF�А�K��l��q��^�P�����{�~|W����S���U$�ꎏ�^x?ƼNa��Q§��H���&!����q�Q#��*�Q�@'�S��t�D�Uˡ�Bh{!�'�Gy�*�-�r���f��/p�O�ـ���̥���-Mˇ�{��Pҿ�c��_��$�t�&��͸��bW�x h��8���#K}��R<�4�j��D)�t��R�a���G?	I�M='.�~������fW�)�d����Go| ���}B��^�'����Y4�tОW���V�T��hGm�����*$��l�¥�p�.��=@�S6�ک��-5�"�4;ZVc8j������N��s�a���M�頸�~Ѿ�Fb���.�Zw�/�\԰���O߇�����1�5W(&d�<L ��y��d4�Ԓ�)��	(�9�3}�#P��5�R?7X&����s\�A�[V�25�M��B�}0A�&�טЩ�ǥ�>p�Y�:I�Sm��e�3"AzT�����o�j��R}�H�
����!��O���UgH>����W���R_��I/������~����p��A�o��^6�$�t��o{+�H�T/��7O��Mz�N�|X�e�/c��?u��xs����E���4�h���p���{DX�T!Ǿy��X����Ei�R5��p=<p���]2�����m����dL;_�ίE���қ�����oJ���^V����F�Y����/y�B�����#I^�		[��
	��,�d4���%7o��÷ f����Z�R�-E����#�;఍B���Or4��Nw.�V�ڼ���:莮4��W�#���M�J�U��j�Im���u"�n��n����`D�+�nw�O������AGrRfP��b۬n'2Ǟu��f�CO@F^|�K�E����>�S�an7�FO�:��<�G7�9�r�{%�HZ4��o��Yqg�o�@�΃:�3��h�5{�����m�B�.(��Y�jI��b��]�6	M�o9c ���U�N�N��#P,��2�^�_��F'��'v9�Z�=�M&ARuMxh�����+�D+��nKq��d�*x���$1I�dr��TR8~G��wm �0g��	L���l����'e��OJ�z.O���,Ǯ�C�&����*�:(�'~O:fF\Y����[Z"�6h�WKu�C�5����.�m��$�9���N���@P�#���^�����-%ZT���<����lq/��H���nn"��g��i"�.Z;��S�K�!�ԙ\�%a����I�!c��GT��?�y��]���.8y{n����!/�M���@�hb_}_��0�D��+�7m���j��GJ d\ń�S������C���h,3�6����K��/�u�遖/ l�[>lW�b�p��8�'0��[���dKJ���\�9?�c��r�קWƯ�E$^�|}yfZ�M
�__X-�W�� ������|�}	(_%�rz�o��x3�o������m�ʘ��gKM�@R���Ó�=L
�6i���Ms(̏���O)3�MW#�(+�=bT��;+;���/�ұ�
�D�q`�d���������1m.����BY�#��� �JO���
�o.����m�]<�y�5��O�׮:�Ǥ2�h��I0Ԍk�߸���SS��qC��Z�6ov^���v��UەZ�c�ƨtå�N<��k���{U�yп�z���̹ۯTi�X$�r��9�L�E3��I����ոMdz� ��nM=hZV
��h�S��kK��D��p ���=�4b�,���Db�ᆩ
����XKg��rn&x�9�1����}�x�h�4 ���y��`����kԼ����w����	�N�j���s�;���.2��2���"{��ŗ|U�Y��F
��*�GY0<Y��7U�l���ێ�3�fD{�M!>� �ì�YX뒭�����s74�i��Ai��y��I'�E�$Un.��zN��xVpM�����4��h����e���I������@U?JPޒ���h�,�Ŋ��À?����j�,/�,^/U�?��r�mA�X�e��F /�x8���mm�۽�C�Y_�e�ٙD�	 ��*n��
P�Tqr���^�����e���'�Iq��t�G�K�2l �4"�����;f��!�e�m�6Ͳ`�/ٻ�!,���,�|�l���x-�R�)�4Ed<n.��ڐ�`�T�ܤ�;��E�H��><N[���Fo ��)!�w�̴q����ۛ�-e4�}���q�*��cKه4�q�x��y��(�F<��t�>C�7Ƴ���a��D��J��1Y}$���=�#�If���������eBTH��n)�Ὺ��	�H���eD��.G�6�F8U�"�����~_~��	���F�.]��[X�1����������Y��?��T������i�]�9���x�:*��c�Jt�"�BsNx[��r}�
�mn^/`�r="�0x���@�3b^���i���H����H'�'=�F#�Z�z�rG�B�1l�,�:9�r�|Ĝ{�ry1A�U�/D��|�V�8����~���<�׷��$�и�p�8E������l��=TcV���}����KzJl�]�/��1��
T?6���l��J��̞�vj�/�����N0��$<W��Z��X�t!A�)l�2D_և�`��$�5ٶ���{Y�.@�u��cg�׻�.��q����q�S����B"�/bJ���Zژu���1��s���e��hZ��R�ڶ��eȷ��� �u�e�b�c�b�|�⤗���k����(5�A�D1��ǒ_n��J1��
D;�DRd�
���{JM&��8��U��{�p���)���'v�|a���h��	Ӊl)�;���&8Z�9/�M�������c��%�/�������@��tʐA���q�z���*�������i���tGN��E�� z�/�NY���i�����uƥf/)~o��?)4�����!�R(�C��x���X>�zi#~�wj@݈ۋ]�T�� G�N@4���tok+Q�N�w�ﺸ�������A3�h'���H(�B�Cxu*5�>)aLU=[���,:�}��ZΦnu�&	jy[��E(,�>�_1bE�
�@�[�[�2aA��i��X3�J�U�Q�;���ݵ�^��;_�Şjc+��r-�j���f�?��U �k�N%�4���$�߸��|2�V�\�O�%L��o����YoQ@q�K����%�E]������-ݖ�.�+�ræ[=G6�:^�T-�MV���Py��:�s�$N������-�P��Xz�^ۘ�y~7;�dMx�F�����X���O��C(�<���ΆA�#��X��#]�!,ݟG��:$�����Y>�T�&�8:u��Hd#+M��.r�H;8���Kî�������o� 5L��Z�p�pK���v[Vm� �����M�o���J�r��KTN��\��%{��7 ��cӚ;�}m���	Rw\�#d+����IK�[�:�������e�-5�ӽ����$I�@,f��l�rmV���Mn����E�s�Ɣ��S���x� B�f5;0�AdO��<�l8)�cF�{|�6���>��+�ZiuRb��䱐�6}��-CD�0V�2�a�it��5xo��5�d��X=#E��U	՚��]�TI����;�ʏ#��h?�|}�z΅@ۣ��h��ݛ�I׉ܼd�ZJqۤ�Q4[3�_[b��!��g���s�D.��r-W�'& �T2�D�Cg��8�oX|����d�E�$�<����#[��;pgԒ�UG�hܱ_�4�l���%�v�ƅ���<p�v�4@ߋX��ݾ�4P�7~���lhnX ����V1�	���~.w�[����O�%as6�Х#���gF8�Q�|�ѤF��㭭*ca �̺�11h�*�,�E�=�N�ޣ��
U𣤞O�f�>����0��D�XN'�um�Ix	u0��p�4��v�f5yĲ�{�U�%��oC#�Mc���I��w�H�:�"�7�������S��7K��o_e�.��"�(�;`���ز���*��U{�#���#�7ή�6��C%m���!TF�2��rh7����n^�����q9ƌ�f���K �8�}
���QT�$�M�Ԛz�X�s�9�>�6mPx��#�u�fU�x.#$�BC]G���		ͧx�m���5-���[�=tj7�2
�a�M�� w�=���d�^H^	�7��i�����ppD������0��1 	�-�O�(�������d(���U�C7^7�8���|�i߾�=��HeEv@���t�Iƶl̺�e�+e"��%�l�E�x�������sg/�.p��5���-!�r���C��U��n�Q��s��w����� 9��'^	�7� 4{i^M M4�L!U��|
:[�m�"֓j��6�����ү;^uE @a���OZS:�n&)��6�9A��7��,�����J)�i"�*]/�&���<�ë��1eǦJa9�L��KVH��C��y�Qc���y�K_�76<j
4"�dz;;~Lt���	ZO
���ӮOOB��;��R���V�0kB��?uɈn�k�&SȞ�r=*P���yK`��O~�gޛ�hł���Є��h�����.��<��F}h?C���$'�~�7|��^#��\v"�a$�nf�� �V@0�C��[����_�]-װ���g6�s?�`��T+ᬧ��ʹ�n�ȯ�yH����歜?��.��>���iQ�.@�.�nd}:X,<-�p 2֣���o�����B?_Q����˵����1]0Iz8���ǽC���&l�aC�!c��D
r�;�+����z��4C�����ō��A�2�nE%)��7����k��{F��7�a�<�ҏ��g�@���A�	���b1@cx9� l��
��(Ror�:�lQϧu��� ^�G�8+e잆0��5����=i��2W<�7�Y�TΤ[A��
����Ņ��x9��J���9���2F��@v�K�(F&�W�>$���A�'��!*�
h�IYO�Z���q��]BY]����=O� �m^�+���y����l��p������<>�b'��+с����Ŭr3�pE!������Q������KK1�@Գ��5��f7�w��jmV��1��s��ovh��(�O�j���jS�C4������Π��E�g�^|�P�[��4#���aO�JI�{r��N�����RI/HD�#�X�+�8��B
��qp6q������^?kE����.̙J�w���G�D�*=}q�?hH�RC/�Sy{�����"har��x���&]��C��%v���"JR��̫���ݿky��� 7�q���n#>ۮ{����U
��7��z�3�E�>�'�+o�w��=N��!f�<팇�I;S`Yꣻ+K��f�*;-)B%>�>�sm�7(HV��)�T����ӧ�4�l�JHm�e�kapE�r�S�v�)�:�҈ҷ�起�@��%��l�]�.���^�̗~��n;�Z{y�� �,���3�u�X:ј	�m8�{(��Fk�W
��ň��q�jC �a�n�O���*�C�!>S:̝؄5D��'��o�6I!y~�")��@�P�d�0t����w�k!�8��/vq��#�R�A��`8N�c�WS$���~B�����o���"m��tQ�-<i�$Փ�9���[IW�bd�V�`�%�*M�����8,|��3+4�Y���%��3W��kBVH���&ZTЍ���VVp�҄�?����������?�-F���0%D"[�~S]QB�QY���X4W��z�J≥����٥�%�xp�m-����˽Ǯ݃�F@"W�Z�s)J3�2f2r�]��
��T| qRU �����Bp��e�$�\mS�4ݞ����x�Uy�&�ޛyoݗX n�N����̶��@*wL�l��;}�D���ٺ2����ﻃu̴ru�-Hl��D�Fv����d���
�v*��K ݍ"�j�ި��5�� �?i��YJ�0���,�AzM��a�-`��x�!��s8�T���@+k����|�ֱS��,=e!m�8�c�H��k"HN���Q�<`�2W��WY�P�<KF����*�6œ���O\g�߇c������v���(�}F��bÃpovi)��B���l�S4{c�?�w�U�&���@3G����U�}�S�Zֹ���J=9�8Ƕ�V�
���� �t�W�9�!4���Wn���T��ז�|{փ�e:Uk)�KM+���DS^�%� �2ë/�q��g�k�Gᅷۓ��ߤ�cFa�j�o����苏1N��U�=5��)�p9�5�d �����:��N��a@k�?>�_ �@���k��p��<��"_����Sj
����.��B!e�'���,f�֬�8o�j�u����p"KZ#�"-��?SF�ם��:9r_	�����b�N8b��� /��W�j�g%�\n���A6#O��A�F)B��:.A�6���=�����M;�B��
���d��I����S.{g��%Is��H̴�BN ���v�6���ش�D�����R��Ĝ�r�Ғ^j�ǳ!%�����i��ئ~���F���\��t�Mj6h
���҉*�5/��[o���I@����ȟ���x���q-�^C��ʾ @�dR(Q��]��1*����濚�NT���� tU8����.k#c��B`��ʾ̆��56���p���/za%4��z��u�Me �3�|��ں�V�k�E�x�}@u��Q�6�)']��pvrm�}Q�jY�)�٘��?"vs�^����8 홚�O�X&��p�VT�f-9a[�˃@���!7����=;K���Nj���5?1��T��R�.��{�B�whU��U��-�U�ha��>��3�)��)��I��%Տki��� �5:v��P�^�lYk'���"g�{��IJ�g���f���Q]TC�h�e��pxB~�h��Qy/N����m��6w�JfK��ѻ�<#l� Ɇ�8B����1xC$�4h?T�=���E�*�$��^"�:�$��03KM-8��K�0[��Wc���t�6���:��/W*n��/�6T�\f�݊4�7�3	p���+�py�-Z�ɭ��h��P?�)I�pV��)���ש���	��c��Q(���z��cױ��	�Y�������ۅM�y�t���s�ɒ L�Z�6&z:7s���o�[��Rk)��(H$X�ؚn0��) �Q
+�,�Ti:�y�p�fC��'���(��
u� fu����niV���g~O2�6%��r�ST1pF����t ���Q�U���d�O�f[ 0�w�R���19U��>﮹���S�pj9�Mb�����1�/��~6�!���1|e���%9�(m�r	D��$�������e��m.���i�!�G{� X�X�ts����#���ܶ�r�6I���ßkBL;������H@t\T�*��e��⠏~��	�H�x,@�O�m?M�p9r��6���%*�
F?%0��>��;�I����K̙c�b����Te���E..V;q8ޏ����o*�4@�a��V��+i�:F� j `�:x|�|��^� ��^ ��x���*�.����Z�J-Co^X�*"�K���F����X,UZ�H�a��s�d`5�˷���X��"*���i��}
s5`�"5�?����?* P��&��#jF$��B����li�An�,�$oW{{�)�WPgx���is
KA���@��T("4N���f�C ��%
1��\�dT�eT*w_N�%��Dg�oZ�,��<�YRC�o ��E�M�}��Dad��D$�}�^�]Ւ�[���;3
�A���Rf'�?��qO����=�>���<�@�j��I\�V�V�0�A���)��K�c�h]��͍6-����Eٜ�d�2L
�[�=���s�V���- ��3�aoْ�v��^+���Ӑ]��x��I��}<���k8��'��o���!U*��B��FL����X`��vҳ]+Ɗ"[(�ӢGLK��	��`L��w�Ê���֭`�r�	����)�>�u�!Y%BZ���p�M*�T��x�xTXP6���Q�s�{��bN�V�I���H���aG���5$ͪ���m��O��'�1A��7yx�F TJ��"m7�5��TSXs��J��yx�ƇF�ȼn�n�'YD��G�;󨹒1Z�"9r��D���l��G��}����.����_j�QyĢh�� Pm����۔HNJ(�z�.m6��:���!6��&�3{��j<�+-D�G~�q|������`�l��*b��ؽZbb������5�~l��iYRb(tfI�"���໻y�v�# ���_�X �]ZF�>.�"�?L��L�/^�M]������W��*�����މ��A��x������U�]��;tu�q�$�Wʊ p89&�KA��k >�����_��oXL#���3���qn������:�����XM:�z��ֆۖ�n��29�;mF�l,���Z/����s\��*�gf�-��x���z��~\���:�荱�]U�K�t�8���*-R���Ѽeߘ7���:��X�)�r@�����'5��9��f#�x�8�]K�Y9��ϟ�A��I�HAG���xx�F�����.���4����[�9��J���z�G�O��;�b��oU��L��-�����)[濰bT+���������eC5ct�`����<�s)�qt49E�~t�?�7�yV�Mfϓ��%�~���L��Lg�Y����x���N�.���\�C�W�����?���쨒/�+ G΂��ܽ�炓�I3��N�N�ޚh
z�eq� ���`�͙��ߛ����������k���b"O�a7�s��N�h�����[��s�)�$�W�~%�����D'%v��6�?�=6��� ]����i2�Z؏��fF1 _�/��5(�N�}Fl�;,Ɣ�dUk��6I=l�]����������C�b�fڠ6�!� ��eM�{)�@�|9Q�w�t狼b�A��v�X��7�����U""6�e ���������TC4d��*��B!Vݷ�p�ìg�A�=�+Z����E�־\��l���E�F�� ��9q�5(h������`�B6;�N�K�y��}$8/\4��+t�������B�"���ɼZN��j6�)�ml��|'����rE�� �� ��,T�p�n}0i��!���OAL�CrQO6��i\����u4�/t#�K�C�J��B���/��&Q�m��<Vl�y���U�}�9�N����fdJ�y��|�Cn�2�A�ָN�W���I�	=��d��a���2a����5�砺\�۔����{�`.z��5a�j<�ԣ��Ť�T������y+��=$��H��@�R�a�QW^�V��n$v6#1�y���/Q�?<$�n�H's`�XR/�O��T��+ݚ~�1����H�9�d)F������I�ާ �L�3���,��hz��))d�L���1�`��`�}�6���A�%R9H>L�k,���.K_(�$��f	d���уV�<�0�V���|P��樶������O�/���޲),��ԷӪN]ݶ�+>���l�5F8nV�\�f�IE�X
>�]�W,`uѣ<?�
��3��P�|���#�5\����R>� ��2����*�n�b7C�O��H�����Ð,��$ާ39���F]�g֘DSm��F�x�~�s���B�q�E�/�/�����y��Ā�&���$C��u���۵x�0�ozZ��}��f��_�v(����dl9�-r��%n��A�����TB �I�Z	I�����&�@�P �@���NH]8SP��-�HH;�b�TkȢ�44�t=��LbpZ�V�C���E4e��J���)�����u�AgŇ�eC5c�< ����,��#�1.�Huc��O��U�
�C��\�u~�=9�%��Oj>3��@�va�Y���I��k��#9���`٢�r�
P-���0�����6aLȺ�/���.l�}��ۍ^{م�by|5�'n3Q�$I�a��{\��Z�'�kK�����~�R�1Ɩ8��ڶ��əa�S*�>����2�����8�\�I'�*JX�M������e<j�f�[������ٚז��1F%��w�ֵ�"~ů��A`0��ϑg��3S��u�l��qMΣ�����*{֧�=?Pw_iĜ��?���o�aBc3�VH����D����Eh���f}�����OE�m�9<T�o����͑�Q���#б\�3�qQL�l�]�ۀU&a:�z;՜�� +þ�ii�~�+��;�Yw��1
K6E�O2J����-�B�vE�=:����Ⓠr���兠�TF��h��߳9$	�;��.����o@��,�=���/4��@�b>�C�W���&���6��$EI<
�p� �l��{ʛ�v�uO���T<j!}��〜@�H���혵���ɹ�P�m��P�a[�l��$������
;�,R�$��{*����v��░��*|�NE*��0�Srv�D8��T��ac�&�E3�^0T@;����?�����;8#�NC�P�
�W*��!h 9��c}N�
� C�Ӂ��O����|�4l�0�>6A�ݷ��M�/����+�j�v|;��AC��Y���b�ٝJ�a�]lY3�8)���I����e+�D�n^A��xO��v����r�^�bc�c��,YV�|jGj9���z׺;݄����,6�ݞ]�^�{�A1g�zЃ�]:������X?]%'�<e�cFقw��)��qi���b�0����9���R[��	K�R�lIB��1��iI�ę\�eX"�A��S"�x��G���F3�p�=��Y��֡V��C����K�6��-�Ӡ� P�X��j���m�n�y�92���c�:�H�x��T܌�Ex�L�Rn0�@�c�Q$������"�/C�q��L�*�ڔh�f�4�:F���X����S��������%�, �%���ɶ0j�a�����Hp$�#Ȕ �1*���#��{�e���M%<�N�p��˸lW����d�Z�W��\��QX�=Z�MwX�A�	�{v��%����m��[s������������USS���_.�ޱ�r;�8��7�^�XY���[��%������`�UI�,��\#���E��%%m3Uk���t�����I��;�P��H�`3�f' y��H���G:{R ��;�@�.g�����A��l�1�|�C�r}�x3�Z.BI`!�s+=��Y�\e��G��p����0�h�Q&L 9Ǐ�%`T�^t���[�'os�3�|e�T:��-v2��c����$��E��4.�_ )\g����CJ͇� �Y�)g�Zgw�[F�A��]��,����쾽�;�N[�+��
�J;<���YZ��ڼ���3#��D�gRw��N�S�dj|У T�!R�ѭ^A^yP�V��,������o2�1�>����p4�?�y3�)�sL��;p�M�N�?&#��q�$�P�.���K���C�6HpcäO*k*m�2}|y����1�N
�Vs-���G_�o��B����~E��|��}qG$u0��0v�����8��sz�':��hy?`'�H�f�E��+Xg�z;?^�2��J�ѕ5;�CF��+J�xFx���4���N>҇
��U'�I�%d��Jԉ���3p�%bB]#d�tR)��t�!tKCa�ɬլ�h�&|��T�^/���,��RWV>]��櫶,3Уˊ�S>n�v�cMÁ� 3T��B��v���7V� kf]{0*��1�l����h�@�^������D��!�iM6���'�,W�q�#�������j�Q��N@�����A������^?_�A��$���$o�[*H���C�"��2#̕4�(TH'���$��'Rj���Dxc���{�V���%�����$����e�Umz��q��Dz���D,�X�7���H�i�4
��g�4�ب�km�FFΧ;3�ǝT:i(����֥�(�� �����4ڗwW���!zP~�������=��D�ѡh 'BF��akx�_���X�ǃ	f�t���{"c��0�����Ɍ����Eb��ϑ��,ŏP'���>K8}�IE��7�ě�3�9�`go��ē��������H��x�����R踍�^o?�4���=��<=-� T�ԡTU�9��ٍ�:�����jb�[fS�'�] ҋ��n��`_���E�:v���ֆ𔅗���6p��w��4ra-2��|�CZ���-�N�XĖ)�� e�(x�j�W^/|u�Z���,h�J��K��I�DQ�ޏu#��Y����z&�g�����u����"���/��Eަq������Wnv���z��}��4�;����3��~�9��V��k��Yd
ډ9)�x�$�;u�: �dGwf��H�i)6��)(��Έa_���%�P��ٌ�l�����tf�:�\��������֢�������=��ƒk�jG�q+ɑ���d^�?̿�[-��N$$�#�u�\��ݲ���E��q�����±��EΛ��Y��y��h4ۊ�C|�o�}d��2x� )&�P9���(}+N;]�gU���=d�u:��LO�$���ZX�kFSʹ��Ԗ�8���41����(�@�Ih����9���rq�H�!��L����i�p��^&�R������_��mtg|�8�=�u�n������T^s���J���h|4�.b�&[�L�1�Ls(��m��%C��V#2R������J��ϢyN�� ;��u�-���[\�M�.�N�m,��|o�v��\�#��MAU����������2�o��gU^��� h�uA~��2�_�hT�'�z��G��#TKP�,�"�XY�Ҭ=����u���k�>�u����;�{%iMtW6B~�8%���M�ax���.��ķ;h���X!ɮo�-�J�����g���Q����,iE%g�m�R'�x/�qkƞH�7M	�"��e����Bc�Ӌ�e\t�}1���N�mnį�><Y��R�Y?�#\��(��Dʎ"���'OYj�B4�K�A��&��t�c��;���F�ۂ�@�����%V
�B�1�q�v��uw��>虚�p��/?<\�w]hZ�l�+�މ+�V��<��%�PNe���ؘ����`X�:m�L4�3y�~l>�c��8��e,oF�)y�I�jc,��m�
�Au���?����l�V���w�om������0���ʲ���U��A��tL�_�5�h�d	�v^�rX�`�0%�FCl[���$R���Ш��<���zv�"�a�I�o �%�%�b@�z<���O^	n�s�m����VQ9%��
�����+��>�tT�^οO�4�_t�o�$8�@��㐙렞V` �v�eHɠ&���>N��r��6}�����/���2��H%_���~���~DN/Tu�R?Ih�,B便\B�c[X�����+d8yt�!�������Έ���m
�D�`��7��;�
BW[��A�%�"�%���� �DW��C0�\��[�G�M���o=l�o\���0��9��#u�[`{�V��~f�ͧdk;��7�A��f�j'H�ίS�*���J�q��JB��S:|V�H���.��ݓ���H���t6�i����9FV�"���@ӧ\t߬*��w��;�Wؾ�Ņ6�K�x��N�s��ж:�jD�pYzE��Q�ȩW?<$���D՗1
K�,B���k���z�:�ʃ�	nV�o�c���"Ң��O�"_"�+(���͉�pE�k�S�gkU)9V��-�U-R��6"�3�2��^���o�F��D�\��-���,��Sȷ�x�\s�?�%��\�l�@�`cf=	�o)�m�����Z]L�:���+ S��ߙ��˃�Yܛ�3�L��/���<��.��O�l�OZ qRm�����qV.��k�=��rq��dy{l���1����ő�'M3�� 7��hN�#
�>��i��8�J�h(h�'h�-0p۷�R�sN�ܜ�`I�<�ƫ�)���Wg�m �](��e\[��&iT��y�;M�뇤�$#���G�P�	�
 �����0�0�)̙g���_:�������n�b<w`�j������/ ���MZ���ػ}:�$ܝ���}���'"[F����X����{�(��:��~�,��2�����-.T��u9L�3TR�ڠ|Фt���� ��	���ܦue��&2X�T�����E���m�*�k�#����N�� ]�_���"�F���ZSOޑ�ye���N�����EЊV����%|�}�)F��5i ��HWƆ����t]E�>͙�oޢ|� ���ߪ�(��K�� ;�NK҅�g���1 ���B$�x*�N�E��j�0S�/��q�dܿ��^<&�Xp�K�t^(��B�6��)QK��|{��RN�G8��X^����CԤm�M~C�8Y�1X���;���2�A�FFs��F�8�mu��!�S����$��8O ӊ���T��[�Y82�@�ٳv8�i�9���̆:�$HD���k,:�U�}� ��&�N�Nk�=ck�߳@� Dq�`���`��g?М�h'�]py����-��Wշ|��61���Iw�w=��D,�*�*ܷ�/����Xṿȡ�("�6���ծ $�V���5-�wz��u��������_7q��m��=�[�A!�;�׆3x_�����YzO5�g�������-7�\�`w�)p�o�G�Mǭ�{�O:�?c���)�Υiqi���,q�AA�c

pd~�-�Gͺm@�cqS5�`^]�!MW�r��j����(���v�b�#� =0V�u�u�����G�>}�yLpq[v���I�\^�=�d�����
_0)|l@�p�o�"��/_�������^�U@��>
�]����B����,ص�һ^]��<�涸"\�R����= �l�$��o8�ǋ�����\N�sei��t�
��?��WfYț'�tC=t>�4�N@�>&\%���}��,��#�C��5�(�2�|�6c�m�Q֬k;��S�؇�!Z�J�El��o���i��G�J ����ȽSw�Bt\k	}#����:;-F�)y��G �q�	?b2�чBi7�F�$�+g�Tÿ�7���B����xK��:�L	_�IQ��\�����u�'��w8n֡[_�G�C�q�y�
D�]�y�~\�j�q췬�S�T�
����K
T�g��=zb���r/泆w&l����v\�.�{�-�fƎ1��:t���`��a/�M��S6JoN��r渎-���p�B��ԥ����e�b�b|�� ��k���S]�2Q%c��[A�5��?��i+L��n%�#��h�x�S'$�Q$A����1�ķW��o�{eH���X����:����]������/ȉ	�1� |#"��G0
������ �#�|TiU�W�S�x3܀q�^�Oe��1!�;�R����z4~����l4G�˒��s����'c'Hӏ�V}iC�9h"�I�/	�y��ʤd���r��"6�f���⧖ʨq&4�@��������.|;�|���X3����!~C��B�H.x4���[Q�*ǲ�r�eױ��8�3��X}���A�ŃfT��!�#�n�����������K���N�VY��3YJgI��մv/\L\q�΀ɬ8�����Dr�hnM�7�H��t[�錹�U��0<v��}���RY�¾���0����E#i�[72�Ac�K@�㵰H7RLGv�7���l`��A��L�� �"�Y[Q���y�e7���G��bu��ZE��k����������_��/;�=��0=�5I��j���갘���SL�!]*`�߹oH$�Z�[}�۪�G���@�?�J*���p���6�w�  !�Dى*ߌ �QjX!p}�lb�R�{���Y�u���J�ɡ��T�������O��5OB���GE��\>hͭ��g]b���\ü�R�&���4�D��46�X&9X.������B�4n��+b�E	cS��׬�X<�&���DO�9����˔x<�w��W�������'��2 B1*���EX������,����� x�F6�l���'L��^��i��.���~�_�����8����߯�B���`����^AuV��U"�^�
=�>#4�9�Q ��K�h���x#_NH�X�++�Fs�I�a֩%���
�D��F��iB��'j_��߆$o"�-�{�������k/��'/V��:��W�P����N�:_/�B�h�V\��s~�u1;�^�u�������j�G��<�P���:_�y�H��9P�@q��t��{/FD�{:7�̀h��w��s]��ʍԄt�|int�RS�]<��33ɾtJ�YqF� X���}u]��IN�BՎ)�ư�t�.�s5���v�&Lv<�j���9[_���:��wɍ�"	��MC-<!G���U� ;�G�f�R`A���(:�*���p	�I:�Y�V|6~�Tvv+{9��.���~�^5��3�jM���aǎv��.~?�Ԍ/���bpiCޫX������-�j/3=0e^\Y(]�!v��g�!u�ͭ�E6:ĜJUE0��̫8��e�.����`���,`;�ed�X���,d�7)y���󳉻�H����FՎ�����LѦφ�[:МO&�j��)�~��'@��δ��q�|�������G|g�A��-�w%�'�bW�Pv���ab=�%�<�t������j��R��X�d	���-�&Q�Q"l�E�����U�v��@�����,�r�_�x�k��U:��u��R��8F�x�9�!eۃ����0�L�����P?sH;�A�V�$�u�qO1��tO��Ki��Ә��<�n:їd��5��
����s9�m��3½���q��
�������֐L��Zsg���84f�k���P �Fx��k/���$.���簋���~l:`��6C�E�cX����{���[����zG9n�r��+��:;=��A����Y6��Y�(�����D�D]���j�ns��B&���W�봧��+�["�zo�)Z"��I�r׍�����!�B���N��vE��q�CE��8ݱ/�\(ե"|��_�j��Դ;�6��]T;��^�*��m���-%� �b�Oq�?;Xml#c�x�+^�ʫ�Gp6��"��a�2��|[nZ����}7#��X��|/h}����+�Ɍ0=n#>��`.DG�]�1�􆼓t:|f ����'1iY�8���5����c��&s�hp�����-���"S'����&jz#����D6����Ց�������$Yʮn4{���5�&�7;ߒ^Q�nz�ɾ�Z�Fli9����h��N�C*@#�4m��(��o����ۺ���(0�X>��e��:�z����-G�$f��8.��f���k#c���k��~:�z{�\g鸇�HxP�\�5,��>�h��"ޚ���/
.W�����ۛ��Yc�� ���/o���)ѫRY5�WD��ScNnv��k}T�eUT���+kFjj������צRFm�l×i����\����=o��@�����<#fy6�:��j�Y����Cn���m�V}y���dҪ�=&���6{�q��M	[D�\ڑ��q����뷳7�������"�IE�� /�a?�2��(�I�{����,�6���7ЯƼ/�7�-��E����T�8�_)!�£�:���%�R����>*9M��Vh�ψS}|�M����>1�<����B�ׅ>�|��n7��J�EP? ��-�U?eNPp"W�ra �wA���ބƅNwJB�1T�a�S��Qtc�n��\H�BF���VJ%�]q�ղ�M-f�7�i���WT�xo@���|m��Rڄ��n�.c�+nJj��"5�ӷ٧B�Z.՗cv�<$�t��$��d
�:����O��[u���֋{v-X"��}����kRz��D]���F&�.�u�r��]�9(�]m5	1A��y5*d�aykpl��l��I�f��}�F������׷=��'
�cp�f�C�Y����}��4$r� ����3ә��ȽA�4�lM��6���ČbB�C�߅%��ܯw�p;��ȶ�{��8*Q�����\����95�� �����C��.�W���;�ٙ�/�M��������n�r`�J�c�#�OQ�
=baez�9 �A�O�u?ƐOI-M�}e����=@&;�2 ��<m��c�,�sC|��1+��e ��CN(���KYCr�Q��<�R�.�H�Uvs{����RVOAƑ�8S�,�e�k���Q�::��[�6ܦ"c����;i�ozk�At��$��S{7��w W#����貰<#DI�A��̛LP�v�`zwK	��Z�׸���}3���Ǩ$
�[�ɂ����}>?+cÞAumbp���]�q(h#���� �u�7��8}��Ql��3NgtgT��f�-%]6�14I����Ƶ�Z3y*N^��p�6�I�Wo޿�K�}�5�Oݶ�[���<��6�J�j���;�8�nuHe�=��J��3pܷR��0�(i���w(�G�s��ֿ�R7����ㄧ@!V�."X,����3��Z��W���z�� Û���o_ �ŕxf�ͻ�����9�#!U�����$���	黏�8���a����2T����T:|,�
�܊e������X��ƬաW��)�L����+�sK�L$��C�m�_2X��|�"�p&�&��l���*�V��j������ O�[]�?�
]�M�-H����2�F �����MCزd�)�7f[(��q�r���w��ш~s���qz)	��9#�LL���A2.���o�Q X��}�Φ�IRZem�I6�7�ͮE���tm-> ��*$Eeꇶ�]w?��C��GK%�A����6��Y�a�{r5��!��6`��C���=�:�������$mG\��r��>cmv��&)����|N:�>����I��$�k���D���9��?|)w�ܮ�Lx ������}X۟�-���9Jƭ�T��3��)ʄ���P�K9�w��r�t�H���+�j������Z�6.�0�7������.�Z;��_<�:��,���q+]��p����.�C��K�w���G'�����r�,!�
p�y˝�n'lր�lN�P�:JP�559	�F�E�Lo����DS۲������A"Q�6铰Ww�h�(� ��9 �E\�_�(L�,sm�A�f�y�-�3��9��8B'r앗(<_K���5�%���βO��ݸ�����褱t��G�&�(C�w7v�Ȫ�dӉ�<y}4N�qV�̧���km��B�bO���8p���4�����X��M�A��_���A�-T�A����[Xk�/��P�2�J^I�L55q���t���EFjO���Q$X��,C6�y1oE끰H��\���j��]���$����_�&5���G���CL��JFHa���f5��m��+�F&�\z��ۚ�4>D �|�7��^2%���/qdcV*`��������E�(ZBD�K��D����D��o<��Q��
��!�Cyk� �K̓�k��s�*���u�~��]1$��@p�$�2�zca�Ԧ�_4<ao$nV�:���[�6�w)�84�Ӓ��FdqeA"�ZJ�I^g���J~���Fʘo��Gty�0%`�3q�a?���q>/x"�z��la�;�3��D=$L��4�r�E����
�D���4HaZ}BE���L~�����|J7�C�}�Q�s����]��Bb^DuK�d��|d�9���#�����c�;�~�S�ȨB�.�C�N��ʤQ&��Q��r��r@��N��p��1.?�?�f֭إ@�^�sfT�I��6�zNf��%�FT�������
�z�i��"M�8��y��F�q�M��.T[M�\z�;��V3�X,��%G7�&�z�f���3���#����l�-�����Yh��9��J���/�&~I�tyCjbr���9�} G.�\�R)n��:!
�i��)��.'xwl)V���?Y��
��gj��`���)VX�s�k�b�'�O��03�_U{�фx���֌_�&����̚���n�p'`N���Ś�ӛB�� P�tE�r�f����˫?^Bl��:h6G�(]5jƒ%��t����s�)��l8�l�Ǟfi�Nׯ�ɹ�� �+�^�RJq����U�k��0� ���.,y�Z�?2�����8�c���9yd�Ώ�꒙���.�,�u%�`��c(5�0����\��
h�*0l�;�����#���;�|�܊������|gI����{�H0i�MU}D�s��%<��w�yJ�Mn�3��{�(��̕1{��~��űfy�2�#*����H�5U������@��#x�I}����$,z(JG��߮��;(�Q#�YiW�Q\�X�TS'��a0�˟a3���l�²_�l�~����t��w{����.��8��&���K�Yi���9���H�$���-U��R�l����J��G0=��<T���?�&gσ]�MOP����}���C��3��>B"��WAy�H|��~��4,seM�[h[Q��EjvZ�����0F�����Ц��۩o�k�ڑe����D���w/�O�g��Rq��	pV�Hə��b��{j�G�FEbo��^l���i�pM_T5\~UU�~��v�q �f�E��3v�����%BN�e�y����mO��28>2ڤ�2�0�Rn�ea4	fnT-���� f
)��j�ƀ������Ɉ����G��#�g,�h�X�J���щ��{��t<lp�q��Д�6��h'BKZ�
�W�F$,;/n_��Y;�2�}$��-_�:�A����o&s�⦖ �	j�eT���w�rƛ��N���0�\������,�2k���s�I�4A�ր���E��b#}�)*��&�L
��$6���$wu�I\�n���JtcfҸ�=�."9�<�G�[Cс[�M�ݘ��7Y�t��D�Tg�{o(���~V.�7�Q<�]��8�����~�Xq�<�掌f�c��m���E�ԫ!0��_4ԚiJ��v-�T{��'OA���i��r����a�Q]�)����@n�"u�K"�a�\�~&�{4"Ϝ��`RIDSX�O�`��!;����A��e"�\)U='���%�%��^��^n�]?L�~�r�gg]��/���½ߏi���G&kƷQ� ǃ������M����×5�}�p�`��R�[Y���b|Y�ި����Jew����a����SiJx�v ��;O�>/�e���y�ۣ�ڑ�Td(�F[��x��5�zFE��C%88@��>��3��P�hOl�`6K��ĸ5K�E�OO�7�<�cm�\�!�	��,[M&����E��5�Q`	hae�����[q$:�;����,=o��Q*iۑ]��w��K�>*�|=O�:a�a�u���s����esVY�EW?���<��*�r܊�	�9�G�{��}�6��9�;�%��c��� �c�{��O�7���ݘJ�9Z�|9�"���0~�#b8�JM�T{-��,�:F�ՇH@���_�x��k���Se��<��P�-v�-��XȆc�1��oR0�6Y���z�e5U�4V�75�V.FV��6�,X-��(�h����7q�.=����*��|(��#У@Zq5ʂ�Dx�Y7�n���X���}����5�?C��8��p͎Z�T2N=;6E�}F�g���vyH=�0�ʁ��3f�Q��8�ˍ��J�m0,�� ~U��T���	J���P05X#�����6��n��OL�u�#q�@(+/k+�z�q�d�[����/t�*g[w�J�t3�?���r'��zk� )��/�^Ԩ?FJ}��uC@�:��h��N��,	��\/SJ/u֡���Jh!�Ҁq�:(}Ф��� ��������y=�u畧�/� 6H���t$��0�K�5.id�G"�t�(	۶N_־4�0}���9�"�f�����=�PtB�.6�J;??��a�����0�f���@Żt���
��#d��_v�^�}�m���+j�}���Q�3Ϊ ����m���b8��d}���9ڠ�46�D+�qL���cwAn��]2�q}Ï%�����d�E�Q9�ֆy�M��$
�LTI���4V��R	K:��x��s�j\ac�J>��{���ՠF%g'�2��+��;�"v�?c�P!$�<���B1J����r�=3���V��i�O��aK	�.Q�r|<^�v�r�݈�[�������3ed<�J�`��	PLw�&�$zI�����8�`�Z�c?1}�ahI����:��\�H}䠎u2[-��z#&����(O��"�suw��PdhW��V�z��M��$��O�*w��BsĦ�P��:�V��UK�k����X8��D�5n��x�U-9ʚ��[	SEWqN�׍�g�}
��8(<�i�L����n&�@b,U��']Hg������
0:�A.�����;(Yz ���ST�>v�L�̽�b9k��5ф���0Q�0݂S�j�Ӥx��t�q΂�;)�W N�X�l}��W��G�I��.4��a�Y\�9��l��%���H�X�H)0[3<�eҎ��p��Ѽ	��UM&rG��2�u��J��Oj�%�M�Y�w3�,�x�Ў����.���T�����!i���� �ŧl&�`&�����H�
�0�.������GQFA�h��8�!�80~x����I.���`i7u.���wd]e��iVV��x���zr��z�"jI�,k
��8n�`�`�����,xŗ�@�^;�@�>��nb�ƙYI
t��ں�]�k�;��!v��X�v�Cs�Q�{�����z�z���R1��	��l�5�MT���_I��յ�N)���)��j/ǥ�!s,ؐHu����2�~F<�;��W��k9�JM��-=IJ��W0�� �d��g�@�,��>)��7ļ��!���XJ��F��� ��m&�������Ç�(:]u��J���4MA��z7���wJjtB��1��	��s��T�(�"�)B��3r'=L4)��_ ǚIDJk3⩪:�4��S�BB��=5<�R�z��y��T��2n�\̚'��OR��R�#"��&;��� ȈK���b#�Y�F�]f.k���)Qg��].�eH1�f:��>]r���z@�����P;��=��Z�}���/�|�^��?�^Y�~��rNX�tƔZ\aU@�W7q�/���e�4Ba���as����,ӂO���v\,��g�?w���?��7_���<� ��:,>:b-tR��^3�g�W�0|�Tۡ^�@ևβ�{����+G�[��A|9i�{]�!xhќ�}�&�eq�`�	��Pk��I%��3�q�M@&�&�΃��A�O�!��/~�
ƨ�V�dzۏ5��G��ј�?$���%9_�R����tP��mu$f�!j���F$�W:�^�6[{͟�[�w�m��%>|��̨|��9I<�$��l�S�=�"/;��ǈ������hR��)�<jr%�_9�S��\i���cg�oX`��(�A		����Pv_xo��e�+ʏ ���*L!��r2����~��p���-���U����o�g*�5��P�l�n,k����p��K��Mo+Rx�"���OTb*���4T�����[bp(�h�	<
S�+��]�+PH�<�r坥��%'w�y����L�=�"LZv�9����Z��?�[��]�d�u|N��e�������()��gnp?˸�2u�cdb�˞фZ=·ӕ���5�sIZ�7��pA��\%����Tσ[�O"�T�Ycr��:���cM�/t�	����!�s�63Y��p�y =�0��2K�}�y��?	Ȟ���S@��/� �ؘ0��,B�4��L���؆�w�Z��ň5�Yf
\N��=�#L��-����n8�_��ZK���5���z�m�ٙ�����&5|���=j^M�׸�*����2�n��э�aY�$
n�TL�߷M�^M��q���(��}}�P��h���01�B�Tc��p���'�NjL�xK�N�� �q=���(�a��]���Eμ;�t�	�F�ѐ'��9pI����~���i{��.����]�����QƜ���<������`%�sq��n��)��Z]�~Ɠ�&}P-�8P���������ף�6 �D'�2���[	�jz�k咤�z��j�B�i{a|N�E�mP��K�����4��k�E�w;Z&�vX���������%M���H����2����^6�e%�S��L<;-f����{�fMk�λ�y�[p_no�D�%�=iݗ	q*P�����Gu���]�~�<Ǟ�j����&y_B�zt�W}:JLI��!���|�C}ே%�۹�업��}�fJ����]ێ�#����쳓���}�Z�ٖ�a���!_�պH�\a�I��BJY)��c��?!���I���b����c�"\���8��;+k���*)e��G-yu5��%�yE|N�n�����z>�545�'
�Ot��0��R���n�U{>@���M��3���ѓ,��W�����Ň��.�\�U�	{�h*�i%�����7r���qjDQ+��b_�p|�(��.�� �1pG��񲟔G�ܫ�x��,$�ӡ2@��\����r2��e5�m��z;a���@?���:;��p sˉ�x�}�¡�l���L8�<m��C�V��)��N�yp��T��>[���\7~�ad�$�KbKL���3�;��(�h6�U��nk����17A�gD����� Y���,�䣋3�� 1�^@��(wQZ��̍j��BlA&7�\nّ�q�h9j9��U�W��c��=��QO̦�ߩ�Lf����ܢKHgT�W�#VVw�s��{4�,~�����cG����ZA� �Jn� ����TY�M?	 ya��tN �2�5j�q�<�V�ш#�K3�/&��-	sk��������V7fzW��p��8*�}VZ��'mDƣ����d���K{n90=�l��� �~����{�x%��Q�M��8�\��P�M�(,�3�\���1Հ �;�{o/3�!���H�&�A?��|wo%���h�]�۩֯u
!gi��$C�(�6�����ਰ2�O��.k�6�S�A
`{%\7��VfE��ڷO�m�h#�J��B����4�i�kŖSn�6�ÞO)���f�v����-ef�pBa6���r@�ջ�o�� �DaG�G���v�z)ߞ������M��w�T�yg�n����Z�W�}�����'@l ��'b�g�/Y34��Mݺ@?�0{Ĕ0��9π��5n���h��g��¾�U��M�y��ЧEۦz�dy&�׭;z��f�F�`��1�)KŐ��xZ��w�"2N�����:�x%P8܉��x� ����� ]�˴0`�H@�K�������kh�ҁ�����t����f��;�$<����7P�i(S|�خ��c'!�hƨ\[���"�\,�Մ(r�-`��J��c��EJ�͋m,3�r(��o�Z�X|Ƌ��G��V <�����TLt3�l���;
�[UQ��V�j��!��a��p�|O+�z`Bf喅���/M�wv��Ҋ���Þ�;���'Ce˞A��8J������P�´'א��l�b'���&�)��,%�3�8jl�]T��/�oZ{��D�t_���]��Y6�n3N��g��_92����UU� +��޿K���i�g�����YH�auc��IurM�\$�-Ey�]���o��N�Nx�A���x�\���
������� _�]���q�qf��`N �+�,.�����ߴ�/�?5����v���K��YB����N�E�!%=�T/x�U��?w�Mv}7e��"�T��I���
�L���J�D��L�C��Q�ާZ}���v�^�P�;<� g�R��*��<�?��LE��ß�dԪf'h�f���⃠������:�a)�i��hȤ
(~���͒\��vΦ�D����$�O;7��-�$���h��8�Hʦ@�F8�s��긓n�KCJ6mRǈST,���.�ȷQ�}3�*ݝ��5���I���b�S�0����ArQD0xf�@-��3l��t|B�	�01��E��*���e�o�(�� t�k����/|��:�%�����`#"|J�����D����!��=�w�cS�e�Z"!�3�p��c�B*A��-�oCy��?ekp&%6`�~.<���X�+8`5W�Ly�p�7 �_Q�8)(��7��v�4j�Ʈ�8̀}��졢�G�f�n]�H'������m$�`��ѱ6�y��z�Y�H���?����A�|WӂVEUվ��:ZB������� �Ƭ9u��W����=���K��� ;\F���}���ۦ8�H��q�eo��2��$��Ә��o/,�%3���$n*����\}݅�*M���@�M���wz8f˭G���qPMֶ��/�o�I�z�K3`���j�v2�J����1�\��5JK"�O�x�ʪLo聑�^I��O/���Rq�FvL]�+e���$ܜ|�A�&ޱJ~��?���3c�iM�����խt*���Sd�a����J>Ӹ"��D��*�k{:*l�4Sm�y�^1/�_#/@s2�!���tY3�1|�Ϋ��85��0ƍq�dY�$2��~{�#n��{��Ff��@:�w	����z���f�8��;�#��N��=�=��$���{�1h�y�����W�^PəATeR�3V�W�r[w�T��+�5�/s]�*Xˑ�q�C�aY�& ��$:�@}l��;G����7�P�y�>Ņ������ �Z�WQ��^m���"��ɶ�*,5�_Ib�u]���<^��3�rT��a��GN��XX~���1o�o,XT�&��#O�f{�\r��8q"���M�N3��TW���+�D�S_9��1PJ)v�R�{�7�k˞��6Rm�}4���FVN�:��lobn�����R,��0�'�����ų<��Ma�|�L�Y��"k�1�r�7�&�k�ڢr(؅�^�|o`���e�P"I`�-si%(V�I�`{ծXw�p[���7�.!j�Cx��y!+vpx��1�4���+J�sZ�*S�9��EP��T"9�ۢB���g��x�X�k������X!G5d�X"��v+ҟ�jU)���� ��M�.XP��EεG���2���#� l`��}R�yh�
x q=6��QV�K�x_Ʒ��d�w+�E�s�[��&�^7�t���(��
��<d�6��/�Qp�\*�PFQ�����r=��I��2�����uWit��Z��K8o�7��պX���J��Ud�����Y��C����o3��<�{�-V�M���턦w�������Va>Nx#|dƝ���,���ƅ�Yj㳚>�?�݃��K�Oɶ��e�xqQ`\���O��9�-����%$�'�������8W�D`���Yn�z}]1�S�X�Á�����f0m�_uH9s�=@��4zr�I5Y�v�;�4��ĺ�!��@E]��IsB����@����-��J�f���h �S)9oS
�3�����R�\����6ʚ���Z!�r庮+/��[$F�y�@�5s�1�|H��"g A"��ɑv��- ��G��q�Ddc�S?A{�s�s���<1����T�>H�3�&��La�(~nqk��=z)E�2b�W�쉬@��c1����xR)��x+�|�<:�*`B�Y6��r?eDZ�u��~�C�Y���p� o�`�~�j������z�=c�-#��z:��}��=/U���3���-��zN�+��j�=��T},��"NV���y����y2�\�ER[V�M��t��<�&e�:�h�Ы�=�\OՎC园�\b��R�6�����˒H�Ⱥ���n��qm�\x;l�&g>���L��^�9D�J,�9�]����AԱ��tw����3�m�N%���mȂ�&����z������LϔeC�Ʈο(ւ'+,|:�y�W&�Yr�����rεH�k�W�����6 	ZU�AenN��$�e��ԻuP�����a$��Ӽ�^��������%���Ǆ��R7'{Zsֽ�%%�U	ȕI/��F��Ǯ�JI��|���הw;g�`��>�~$����On�t0c
���7�?��
V�d���L�%e!������A@�FЯT��j���$ vxM=' �<����OF��g膴S֒!������r��b��chVĖ���0�N��3�XT~OVʡ��*d�Q�,���Z�!X@TDv�
���_88�]�����t)@<8=t�2<̝���ٚ˱����P�u���ƀ)O߄} ���\z�$��~F
�^b�żf��*�l�D����E��ː~�2�0\�w���S�>d���>T&�Gl��-!�{���7�R�j�d-�b�*3�L������9bc��,�6�ib����`H�@��s�pP��js��~:[�1��Xr�}(�����,�@=�=�(d^ǲ� R�����ؤ��]��
j��&�1�56-}U��~/n``Vm�V��#����pⲇ�����d��O�u���y^�N0Y��!|%/��c1XqJ�'�ҏ�PIϡ$\Nu��r�����!=���H��Xɀ��J����	�gx,0V+bL��tv\JÁ�:���f �$2����"��?.�qD�<��o c�nG�Ng`Y&�u4��?7�)�-_����-�l�ὒa������|zLe�2��"�+�G�[���=-��L,��w�Ά��ZDN�Y�d�=r^��U�l S���*ь]3-DA+07�9~jc���e�=U��ǥڙn3* ��S�:����YZ��q-�^�~Vx57�Ed�/��"Z��"'?1�n�r���8�M�q1����g�9Y�I�0[f���$~\3G|R4-X��,;>�u�pc��D�#$�)�u�qe��~���%^���p���O�J��,�!*G���Ȗ�o#�C,1_�[�p0x�pkـv|;Z�D����8�_���ʪ>.�B<
�� ����N]ʈ��ܓ:_ ▉P�����2('KH!�ջF$@��s��3�(5�w�˯/kf�P����5O�ޜ��%��M�,�Z��ܶP�ن����0"�:KU�|���C[��M�f�Ɉ��������;�րG�D�+��r�N��c�$���ֳ�e���ys�t���LT�᜙t����f̶_&�SW	6�^�n��F�R��n ˦:�.I�=�@������wx� ;7X��u1z0R���V��!EԶ����$>XA8m.s�sE���`�--��a��������LK��E(�<���s�媄�,�@̔� ��Qn��j�v|�5�2����d��Z�rM�v��hl8��X�E�΂)�@H^�|�2��N��8�`�礏�V��Mpj&c#U(U�63�o'|T<\
��6ɘy�s͏��6Ϫ��r{:����\'=	i�u: �汬G�ű䍯���o�B/�1ö��K1F��fhm$_� ���~�}5��.\���;@0�OsD���˻x�DG�vL���:C �+�z�-[Qu#3����cdwrD���<|���FP���\��9�w�'yc_����D�?CH2�Y��nNԖ�Z
��GU=������X�}����4�\oh�ETsQe�YI�&�`hی��ܬ@��n�"H;�G����@�����7}�e8�m*	I+R.��%�=S��Su��pT�`rL=�7��y���BG�����C��>�9 ��eN\~�)���&��'ǫU��*��e�Ν�Vyi=����t�k�-��΀U��.`��9�6Z`g$Y���ʩ�]���	�ؠ9#�q����|��q�)�H=���>�&�s���_ �a��W,^�ϝ�lꃫ�>����u%G��n����G���-5*l����C _���������NE����ʜg�誛�(��[���0'��һ����U��~J��ُH"�.�Oz[��+�:�F:#y��[�|�)y��o�̀體���[�	�o���GK�k4!�{�i�g����K�~�s$L���9����E%Dy�	��r"9�"�Z�<�v4�k�������x밼_*WPD�H�NT#&|mu�8�;uۂg�G�D���FMq�V��}	$:J*I3R^ڭ<Cd��~�&2��}H)��Ķxqq��7v�<�ز$�oNO؍w��հ9���Q���d��L,i�)n�M٤*n��$"�:cq�	��o��C����I$ &��J��@7K�h�p-eiTF�F��`T�djGӒ�b��Q�d�`���㖳�����@�.��y���D������Ǻ�ܽ^�J�:�D��I�%�׃�
�|�|���|z�_�y!$����c��Ü�,��-��+�+z-iV���CC�:i��� z��DܣK�J���2�u����2�&�J�'�O�V H�<�����;S9�>��6u]��� ������+Xp����������e�O��j���������ʘ���ή��{+��ps@2����%����Kȣ�x��<��|�`;��	���Qs]��ؗ"�P�Dp���\qw-�hEY�mF����~�A��~��Y[Q�R��~���	��5W7�%!z}�<���!@�jk)/����d}�n�tB����5�\W�A雒��J8�x�L`�]P�&,����TC�����H�����t�tYҳTU9�܎A�4�\'H��;3~/����J�#j�=���6|�Y����#�I�'���P(}�W3bI���/@�F���FJӝ���s.,u������>�ĵ�n�Zp5I�>��L�S��i��m> c�9�g�� P�ձm�ȕ�z�	�!����p�D
�$VK���M�M:�&[h���ܶ&���w?7s��Sīeo�����K?�'�b�ދʭX8�cW�'��s�_�L��L�����%2�8����f��]�]��ǛS�'����sf�O4���t�^��;)�1�\���{_�i��9{x���R@�<GG��T�Ei��.��W�i⎱�v�".$����#��0$�� �l<� ��%�AYI>f؍}z�o���P5:5�Oo��8�f��
b��M�RT{dˡ�tP�t��騖ΠL��+R��Ym����)�O#��J����!�Y��hWt��m����7O�����a;���n�2�?P�G��cʞ�mG���ܺ��8�P����}.l��>��#1M崉����hk��@C�ӌ�����<�~�����1��2s��z �=�t��}��c�l�� 
���0پ.��~&���"��������كT�젰�%�G����"��C�c��}{�|���v�ǳ����ұ�Ԃ���Zs����,��m��.��XD��[�k�o��sL��r�.>����5U�q����/�kH6炏L�Ay~�N&]�&���D�Ɛ�:%Z�{DV�
�޿��ը��="��J��b7_W�NH��AY|���va(\��&C*C>X�7����� j׉��٧�_�7O((����@\U�υ>���Q?y����y�ɾ��d��>#�R�T���ѷ!�eUH=m4��Qꏎ�%t
�=�s�4{3]�"lF�L*�(���/~9�񒮸,֍ i�*˟�Ӝ#�������}D�T�[���n+�:�x��p�(���U��r9Q�EZ�@�,�mO{��%> M���M��	�ȱ�ԷN&�7��{��e���$��c���v�|G2�C����teDƮ�Z�u#��W���f����,��\ӎ��Tt�P�?��9���;��[|DY
�Ŝ���t_(��R�П�(-����+^�^�¾;��������4Y�M藊�U�2rX�J9Od��>Ri-���?��0���xJA��Q#�Wu:&��u��~g������1��H,��J��+ �sa/;ʟ�G�`���a�1)D�UQ�A+z���m��I��Gͻ~Ey���������x�T��	��у
�A}Yң�*�� ����m2�W�^�'�&)0���?7���5J�$�Z�X�#Nv`�u��LE|�9�C@M�کDZP3�GaL����N�����O�8�Y���ܑJF�>	�5k����2]�"�$��}��g�VQ�3�k������Qb�w�d��N�Y�^�����)���@[tD9�q�o�I�J��b�+S��PH��"-��k[O�\k�u6�ǒG�'�C#�[��a��7��Zz���%���{���(-�UU��,r�3�F�Q�̏�']B5����Ra�ů���@cRO[��
ݙCܼT0"����������W��q��g�v��(�ĥ�rr�/0��ќ���hǉ5�l����C�te�9"�g�P\�ϗ�6% �ۙ�WK�sC���S�<�����md�7�9�[��R�OG�9��ØՂ�sܚCtR��������H~�Wۇ����ƻ�����Y�
$�S_]��u�EM�4��p�r^����M��6K'f�lc�=ikI�&N�l�^)���JV�����c�b"7�H�e �Z&�]�T#8��ګişRǟ���7��k+<�[G�7�ݟ�V����	�>�s�L��+$�}��o��Ӌ����0�G[�
�ת�4\o�ҁ�ƟQj��d�`�a�֤�#e�����W�����&n��ў��8E�ɇ�j' ^QORW�^?�HNH�:��ծ��&G���KoY9�������4M吲��gbD�d^ �
�6;}�ip@�/�#��c;�~�sTZ&y�y�ECއ���`�<;����k�O��9�^m|�eA��)��ߊ��ܜ�1rX,t9���U���ul�~����C�i6+�8�mf��@����Τ�H�Kغ�[��J�s�AK�{�?��0ǥ/H�pl���/RE����`дB��#���
�
�QN{\�e���S��*����q#Cs�o�-�BV{�gQ(�TfN^�����s'U�f/_!��s��9�RvM��>;��Nt�lܵ����6.�W;�"y�{��x=c���>�;_�Bb�J.�T��vK�3E?��a�zL������_Eӆu�Q�+���/���1̈	�$�������|v�Ϣ�N�q�G pf{�<	�r��֍#{,���S��f�pv=E.�_�sIHaT9��*U����J$��6���^�J�["�3��aS:�	@�	Z�Y.|ʺ�P��7i���B�`�{�[�
�(X�`-۸ү����[�~���|1�S?gOF�{`u����Ўr�?c�Z��R�rv�STs�[!�/<��q���*�#:�t����*����,ڶ6h����Sm'r!�^g+��Ol8�S�?�F�?�}�N���E�P�FYV�r`�rTmk|*�ዏq6����ki`���Ѷ#����.oBi#�������};�5oI����t��n�&�YS����$����U�<ykf���:Gd�����:�R5"�]�ء�]Urܣ)�c�1����S������w#��EE�t�@��:6�`��t��o3
��igE�{�dD��\��	k�0�9�I$�R&��BM����ɒ=C��1���DR�z�/��HJ0kUu,�k�k���A���<���S{'�9;�	��S�Nq��~GT���Q1��Zzb�,�Jw�����[��k��΄���A��������R�t)���1���e�~��0��e���������9�ߣ���h���g,F����G8�|	ǶA;
���5u�/g�_b�b��Vc2c�!��u�@:��~�yn bRS����h�a���hDm'�(4�θ�D+�G��rҭZ��c]����,�EuP�X�tk̨���妾P1L}��S�U)e��X�C�~N���j��'��1�9Py��=,�98�&9��:$����r����рl�J2E��	f(�դ4Qx��=���S ����7
հ@薥ʾU��
��+����c�@]%^��)�&��T���Gt{��}�6ٴ�����"XG��fٝ �z8�� /��]B_?���e6>�+α����8���a]cm�:�2��ϭ,*�`X9��tJ_�ORS��Kgʍd�!)��� `�u���V�eCj���?w����:�hPV΀rq�f�t��y� CU+�Q(��F��Q��q��;�+KQ���x��9�йh Z)�fo�S��|���<��T�?{$p`��}��]aX�1��H�Hͭ�5�B�e�i�B��b��I����Q�d�	���Mݤ�|�+���y�H
��w�E��s���Ze;T���#2�����R��]`��N,ѷ�����B�-`%�h4Wׁȟ��Q)�r��@���5C60����g�UR%����a��l꤫u��1s����]6��n#nu��{2��檦��x9�� "+�ǈey�s��P�N/�,4�H�t���(���0giG&����>�J	-7��Tɿ�Jd�.��7����T���n�X,�4�ZJL���!�'�lc|�����h�V(2�%A@�3�o����6dZFᤎ����������s���K������7ץ�b��9\\�/5$�?�<#h�B���&�v�2�X)�A�ȸ�z�-�E�`��nP���-.����ǟs1C-0�P k�-��  hf����z�^M�kF�qA���}�bSxb����B���NP�|:*l�ߺ�����ʥB`pR�yj�q�*<��K��C�.P��w�����m���_x�a�͂��r����1�5�e-�I<�7o|�佛�2���c�P?.���v!e������Y��{%h8�������c#�����~~Y8(can/��u2mƪ� X�Z�P�jj>9���9�[@
|�M%%.�	�e2V�X�ɯy�a?��+eO:�Pz��gv��;��8�4CrH*�L!��/�����6�^*�	��R�m��@��SG>+3�f+�@f���4D�`��=�[�?�QU#r^�8�d@U�ĤÉS˜Ν=������Y{�_��F�fh�!��vQ�r������9����5rxo-O\L@E،��a�w;$�D��n�6�ak��_.�|3
��/��q+r⏶�
l��ͤ�|��@CY�C>b���*ߊP5������e�e��
����D����͵���*���g��h�iV���{�q����,���+�JMG���(�st(x'�x2��c#����� ��;�6�Q#��.�+��!پ\���_����8�Q�؊�C����`m��|)
Q�!jD(v���-$S�w�,_�e���vY�~̪���_
���N�	P1H��M�>�Ë��E�����c���y׾i{h�6�-0�z���u��IG�u3|�^-�Q��^�D�Z�k���:�䐡�ȁOW��H)m��|eP�v�-pM�I�oE'�`�� p@�.>;�HH(�0&�gK|���v�T����8�}�1�_b ȡ	W�����Đ���=��E?@@+9��Z �*���${G��>e��h-�Ab D�42�v�����Ny��	���,65�N����˰'<̃�q��̑?-�����c�柼B�E�"��v����^�Vc0�ho��:
K��K�J��O�O�N�,6R�[��!�*�[`n͹�S;��c�b�U!�k#߮��PUI�x�6΀Zq?�Tv��Q�������2''M���?Fg�T�E�O������3t�@%�E^,�q��ێV���	����#޲�/�:'��R,m|�jZH�B�q�����h�h�]P����Ne�7a0��ˍ���"��&�FA�r���nI�Y�Y�c-��%�'���Hy��.��B�%i#�����q����\��z�u_���;�@�P<�t2��#���9q4)^�#�Y`��~5���9�߷�$�3�,kH?���T-N���'k���1gz��W1�O��̽|��{�c'f`Σ#�s'��p�C�[�4��I�Ka�bY(����ɏ�s�0��u#��90zUo�����"t�H�u�/�xƠ�db.L(cn��s��6�e;�4�*�~>/|Z���΍=#���9}�1�?�=��-1��I��z�Wv�tZ�i� N��T�g^��n�!��ZCv�k�6 r)�����+�ʌ�F��L�3�`����$���cwI����h(��'�Y�U:x�:�#�2���M�o#���ZL{��fG������������]|�3)�qs$���"�'�r2��y9���k�X��yT)(�FC���D>p����q�`*�\Rㄝ�9�rԛް�VX$�bnEo�Q��6j�\�OX�}�j���3��#�Ք+F�}�)JI��bvb�~������9�F��C�$L$r��dfݪ>3ib?�� �F���o˴�e���v��fˤ!����ut~r��}1yR1��a,�,iI�`y�dORgp4�aT�}��<���z��?��}{�w&�u'nf��b��x⤧A�A�$�݄�%9ʆ����8������T��D��s���#�g߯��`=��{�wd�˷6�r���aӬ�9�(�9?8�l��e��)��<s�3����c�#ZF�q+��oF�
A2��4"e��KA(T�����L`h���rmQ�h�XZ��(�1���袂�]��\`;ȝy�va����O�(��xP۟J"��J?��Y��#��#03W!�������^���ν$T=L4�f�f���!�C����)n�x�[[����º�C�!���Z��M-'z�+���1�ݱ�ե���g�.4;Z}�/D�|$-:����2��|%���R��iG��f���9 ws�:A�U���%�rW1�N�i=# _9�gJ"T�*�j���� ��q��3�����5�뷯}p���p�S�Y,V�b�p��pd �<�����otT���:����/2�#�rو�"VJh�\:M�xr��8��E����&�����*�R�q����P��.1pD.����	fgF��6C�{@�Nͥu�P�c��y�pyH`s#�WU�Upn��{ҧ2��*۱��M��x�kSr�o���"re���yu�)(��!����lRJ���:��%�����^��p��E�da-��O�qkim�h�T�Wh�Zne�t��J4�����ת�?�=UI�BBZ���.M|�z>��d5���"��th'.i�t��?@<	�F�Fܽ���"�i%��A�rek�!��f��L�����1�I�%'p��د�� �Х�m�c v	`�")�K�9<�kۧ��؏�x�~�� x�GH�- x9��%��0��daiW[���R&�j��	.�l�;�CY�������T�ǆ9����MG�5;<-�7��E5��h=�x��H5T�p��Bן��f�5H��v�I)����1t�Oe���t����"e�������4�!��lS��zh�@1��k��Y��R6$7�3S��1C�m�In�\�J�pf`�#�� qg;�F�$WҫMK��R	�c��Fomu&�P8�Z�,|��Q���q��[=������C��r?F�\�ۨ�vX�⯰�a��b�%d*,B�`���(c��>���7t��s�g�i����_�(��d�����g�����R�Y珩a��!zY�m��}�xEqEڦ���c7�Ҋ)��*Mms�Q���7+[�mŘ\?h�w�!�`�0E�rŎ����Hs�j%���x��,�@�y[��dT<R��K蔟�YI�Cc��
nr��繑�����^fȗ3��� �C�z�;�
������=U�*���B ��H!-��B�v	'�>�SH36�Z�� 	����Q��o���o������	��mlj�R�=�N:�:ˬ���*��kp~n��eDc�#;����0�XE��=�����{�L�|�[F�2�m�U3-�N��	�H�S!��d#o�Gْ,XӺ��*$89�N��X{ B��OR�+�U�L��T*��A�*�R`���@3l� �J:�%���j�8��Q�}� ��,!'�CV}�Y��yL*u0�$�،��;�h��X>�DD��Aġu��&�zl�K��E ��5�]eG�s����o�"%�asR��uK�ƲPuAb����P"�-"�Z� v�ش		��}2��2�y�Ё�49�`����Q�Hؕ:pe��Y^I5t�jc�2�2��^�)~��1�>]�,.&��mX��M&?)��5﫪���Kt֞ca�c�G�֤c��7��j�K~b5�"J��|_�Dc���Й�s�@ p�B����e�@����n�d!�Qɳ륔�#�w�QAb3$��8j$uBAAV��Tn3��p��!~�4ƿr���Í��-�J����v8�N��t�@�t0}�k���w���_���=���I����K�ıe���O�Vx{W(
��Y�~E��P
�$:���x�mO��R��~�QڌP��<�
�Y�@J�d�s���Xu���b"`)��X��ϡ�%��D����\�oq���:��ڔ�Y�E��aׄ�_c�o�.�}eS(D��ۯ[8�ٔ�1|ˑN��!*��|ea/$@�G�{9�gZ�.���)"Qd�vw�^p��.?�#e��r�1$�+d|��(�C30�5r��,'���vX�Rz����H����M�M�@�t"%("���{�ʲ�=���`{���,?�������B;4@��>��P�yfX��!Q��Vn���N�-C�Je�3X7�*�r�kC����7�(��� �㈂��!O���I���ca�#egQ�]�����:W����nX$�:^�뱌�
@�uQ�f*�#�H���RS��pN�k�u(96��9�o]u�����8�,�v��Y )G6��w�:�l�����Ʊ��:G���r7�t�6��~�RH����%��0�[�{z�;ۇ�H+'ۯ��4�wΦkY�<F����J���b�y��aךG���!qn�R`frS�Xu4y�<�Z�*A�&U��Л>���1�kꯎ�P�A(���X�qS���bQ�����A�����}�#�D���L�G�x���밣��)$K�Cf)#?20B�<��>�dleC����W��p���9FX�aK�ή�ۦk:Tܧ��M�^n��D�@��"��^)�wq����8m�	�%�%�v*��w����myqGq���w�o��G��^"^�k�M�X0��Z�:RP���ͥ�]��م^D�xN#�![��WV�\����$�p���;�0�a����S�.`g�{�FzP�]�?�;�V�ch4��Qn��&X�e�;�:ol��>�1`P����+�����%��Z'��4���SC��%L��mo662죡�]���ާ�顂��f���Q�1j�7&}�M��������A+ְٜ��^�%|C.ZMr|󉑹��(�/�j[<m��|����.'�D���Bʑ,ک������sM�8��r͹aKK���g�B,���)�0ϩf�[1�/�A���1$���i�X�{=?��\���+!�2����|����l4~�У�V�\p�hbrHX����� ��]!����V�ix�L̰�>v �/��>�����a!�\�kiu�#?��-_��~�d�I�Z۫��]��>2�������h�	\�䫓�×��Ñc_�cV�|��ֵOר��eT��^��_�0'�膯�u��}+s�V۳�����2u�w`4�Z��K^���W7dL��ف�z��#��N7IX-U������A��O��|�@k����Lp=W�Ѡ;��^ݢ��1�'�$����-%J����'h�yY�|�I�Pr�p�����G�r���H��@Qɝ��|�pK����:-$�+Z��,m�ET�Fȭ��b����O21�т�[��+*�9>H�S{'����R���P��LV_;�8F��T}�09;,��N@ﷀ��ZM�
� q2MdX�^ڧ���+�������(����]��t��<]ȕF�hugHhX�-�0%��w�Xo!��:JC29=��D�P�h�.NU��2�3����i�[��٦�cA>�qj>%�=�% =�XY�3�ctUX���A��4pf36� �O6\
P��� � ͘�8s !-��y	��B��Ҽ��V�p�������J�k�M�]��r'�L�m�u:Z�H�q]A�R�)���O�sޯ~"�����!� "*�Z���R����/A�|D�v6ޮ?ɷ//h��%�9���3�@�L�6߽�D�[�ݑJ�O1�������3�;���C�Ce,&�P���c<q���[N[zm��)vg0�0�4t'���I'&���jż$�!,|���������;��:\�?���w価�<,�����I�~w{E������Q̒�>�1uL��qd��s.F�~}�������$���Gt����3�4�8I�r�7?��ּR�]�Bw�!7�μ����}"]n��H�#���3��\_�<H �fN�݀��@`P��g�����4�)2E�z��/#$�;�2Q8�@�b��ڞ]�Z��,8�Kc^����\ ��΄���s�;���&��ؚ��1{S�b$�Ӕ�����@��Ky�k���mObl ���"�q��U���
t
l|M���W��}��+Ϗ��b�-��<��
v��9���Õ?G+4UE��<�$k	��:���
�l=2�:!��"i��
��!����%X�����n�6�:n[���[^^�`��C���x�I�b�G����+��MpL�F�f��w���l�∴�Ǌ�+�V�>���r���-H�Ҏ��$SE���S܍�J�9�x"��J[CK)�x�P���}���|�2����5���Ζ!
-���;�+!wL&�{���?�`��Q&��h�CU7.�Wl$�O���F��]ͨ���)�=;�$�+��栴����D�nu��ձbv�v�8O� �>87(7� .L���6����k��$��=q	��� z��_/��ܺ�&��s��G���
� �7�N  �2��S.� d����V3=t�*1��٦M$�7Vdq��~��a?�9�y������9	�}�d_4�3�b@"�~�O]@x2[�o�,$S�Pg�����2Ԋ�|qB�YH�|�I�xv����A��˿�[�y��k˽�|�l���e�-�cV�4N�$y|o���e���~[��}��sl��/ߦ�����mI�������j&���ps����%	n�!�ZU��e�:#�z�I^nY_�iG-�#�y�Ep����f�I����H�S�|���j�h�qL�V"�����O�[u�w'�x! 6N��shڙ��m��}bA�8�X���=o���H
գ��'����Q�Ps��'	y-tq����uC#��!����W�gK�5�k��`�-KZ$0$����B��$7��-�E
�7���.���<D�q187�|�_hl��DJ�y׊)a���65��eG��̆X�f;�w�i�}�O��l23~��l��S�1�Ε-z�2�W�G޾t����J���c�Kh>Q�r�e��<#�{�5l��4�N��Wp��oi���a���Zʋ����	đ�&�b�1Η��oj�j��M����G'��B�o�K�梉?�ŭ(@Rz���=�<�}�?T9�z#	�G@��r|JJ5`5{��9>f�}f^���n��\w��7��E���{��-[g�u��/%���r�s(g0���@o������Z�;_�K���F���[
ܜ	r��YN�a�.S� a���o�@ǆ?�l�}Pz��<Xᚿ��� �X�˛{٩�b���g<!���Z>��~�7Jͬ�ΐXͷ�LC��&Y���eP>��,��?E����X
��嚪���p�df�Y�LX���)Qk�D��`�^�[y@��dF��YF���`�[�;l��of��`�ʰ�X���k�:B��=��O>(���؎iY���C��q�,���;�<���q~`�`��e����ņ��_�#��yzϙS�mփ��
�����l�]/p&yqS�����2�)��"��X� J�̓˶k6W������ęg�<���k��h-��X��_-C#u�k
r�5<��Nǚ�NM������r`�r�$��ߤr�%,����Pr�&��9;X�=崂r=D�=Ѫ���/��z|F�ފ�X�uڰ3I� T��	z�q
��?�<���7�0�n��o2uȈD�5L�bvGX5��dZ���!�bG����Rء�魆�W�hi�&Jor/}Ys�y�YJ֗��Pb:��%*��������qN�tZ;���Kʎ}6OJ���n��x��C���^�W�H��ND"w��/~���؆"��d�"���LG��Ũ~(�E�r�ճX��	��4q-C5i�)p���i�U���1҆IL�_4�g�����xa�-��y�K�2��4���9��	^A1B̉C@�l'í�����"�q�8b���,�dSX��j�U�1�'j��֑QEGx,�v0Ń����m4���df�vˠ����\Q��xf"��c��z�O	�6I%��r�d)V_B��{|����h�v�2. ��\>��N����U�Rca�t����2|�+Ş	��K�C�Ko2���0
Ot�i��q�9o?cZ�1��z}�|��I"�`������G4�����
���*��}��W��UcmBw9v/W����0j��y�i$Ղ���T��eʱ#�2tlW�{C$�7IY�` �w�� �kʛ��+�aK�0,��4��a���%��٧:^���1:t�[fy����Z���A�D����?���ۭ����p�z�A��p'Gz֧|j<	� ��|��+�+|)*���!��+LLh�w�Kh�1���B�hoW r����t�kw�Z���17�(f����� ���Z,<.\�:��z{*0�91@������o��!|x�C�l���n�SQ���YIk��$���G��u��~��q�����-�������x����j@���	��wu����9
���CMk�3 ^X �Ϋ��U'�S�A�f�0�R�p�6JT<+ND�����1���vs�3��߀OCٜ�zC�@|]���,$꜆��)��Qk6�2U�+�'-9w�s������Bu�j�k�.j�,r����H;�%#��+B|#�"���0�����;��R�k��(�g]��F���^�Gu~�E�R�)3��������-�6
��!$#mc}�N,35��a��BR�G;���QGy����Q���i�A�pI�(�~G��n@��&�(D/m��@�s���l�=<w��<�`�8gP\�b{G���b��H�t[����b���:=��%L���pe?�x�k����3�s9��@�k�ky�L9��>h'�,R�`Hfp�0;�#���Hz�R��ZZp��aI�o�Z�q챋����U^|��%~��8}��~�B{��S����Bڞl�evgs��-h�S��JP�H�������1MiV�pذǖ��^�kx��g�ǅ��X���@Utv���J~�,�`�W�#e��҃��8c�0����\���flv����*�*��[qL���u�4��u�*���Z����?��D��3�+��X���Q����@��w���v��(��
%���*���PѦ�r�(��i;��yY�{4��U������L�M���T�☾W��va��!{>��uj���\�Ӷ��٭�s@õ���#<�h�A��"�>Ƽ!ѹ[��}m��I�D��f_�1�^�g�e���&M.^��F3]�fE���0��%��5'%�)}"ͧ}ؘ��ݐ�1ӓ/#�U8h�2$
��H\хx�����>�P=ĭ��K��
��� ՟���9$ko�A:���49>}^TU�Pq�����U���z{Dc��t�>!��c@�����^��(�$���E��|��uί�S�r�~\�F=6�.]Q��X@+=�xH8�r��N�������b�7�`����[�I.`���uh��]�M�Զ$$;w� �ʦ�9���
�꛶IQ��C�g��=4���ՃG�v_MX������!��/�j�j�8a#��}�ϔ�4�,z!EG�O;hF�,}v�`�ov���'GC���7l�,�A�-c>�gr]�}�*j	�Fǃ�1[�I���+.g����)y��7�������ʦ��z >���s�������0X�u�5�9h�ۥ��;d��5��F�>���b����r(u�	]�ƣ�fOt� D��Ȇ�V��5~�{w�x�G������jJ�4w����K�
�.ڤ
�3��)�"+Q�rs�Ƣ���
��xԮk�h�:#�Dn��	�t��Fb��]����1e�`ѷ{���n�����OYut!�>�y8�˶CSH�ߪa�z�b�NJ���C��d`U�D�6TCA��,�ػ�����\������Q�0���x_�����	b-�V�y~M�
v�]g$�a����+�ȇ�L����:��%��h��_��7p%oݻ�5㗪gO�z �7�0"�û�e���=�&�y�ܾE_�@��)MU1]2�)e����v� �U���'�+zCD��^z�y�̜��oȓ_t~���B���8����E_���s�u`L;�O���jB$Y�q�r���^��u�b����e��K[=%��]�Gts'��{J���\�&N���&��Ϲk� Z�䉊���H���~�@��Gj�α"���a����f��|Z����wI>��_X��]�Q�>��"��#�X`OJ��+? f	�=�{�$��`��x�>)<ȝ\��L{��LvӒݵ�M\��9��>>�&F��:3�`�$����6@�b����T�s�<?2�#�͸�jE�P���G6�0ӆ��QOC����!q(?����f�aoS1��$>�����
d�^��$�����]rox��YP���og�\�H��>�=��`�XN���6�����c�FpN�a�8��E=��Ъ��i}�8i�$�8�*q���P.<�Z�H�� ���b􃂜�H6pI��?&��q�HY^�<:W|6�(ۉ��@¬�8�$Ñ7&vP���I����I� P�BPƌ��,L	4�@�Ҡ �u_%�����Ґ�b7+�J�|5���B�������T<���L��R\���{
(%n݌W�c�%���:��4%brE6_�l�-fΣ�~�v=O7��'��������?�j���݋fэ'Z�T��z���I������w�����p��8�F<תּ,���F�6S|�aK ��݊m�i���0�5���&߸S��� w m,T%�vtudh��|��XLb2��Ӈ�6�æ�2!������4Ƞ���B��;�G	�"憈u�;MvP	Ħ�	�/}�l��e�O(D ��^�¥ �8�kD�����o4���=���1Q^�tR�|�u��V�HkL�����0�퓷w���N��G�T�}pZE���"Y��&����p�W_����1%Z3������!�.]�Ӷ���U/h'D)x)H�˰$��c�)e+��
d4�`Z��s���n0��	
 �׮͞�p�t���9�֢C�z�N(����FH|��V[�Q��}�'i��ܡZ�2�x��]Q�ݔ$;��jf�/ ��U��y�y��v�7#]SL�
���Hz?��~�7쇡6[�b�ML%:�cu��=T�"�҂�1!ල�6v0��S�����(o��程�4 .������_t]��'��#g�S�n�n.�����`_Ju�S�'g�iM5��O6���7�_�S���~��9��z�̷��Z6�{�������t$D�ODk��⏰�����<���S}�!��C�����S��{�NBTʼ.0�k'�� �V~I�=Ԝb�mc��H@}�)�z�U=��#<k��f�q��,�lW��L>d*Y��Vۇx�g��#�o��yE� e?͞�g��%1�
�5b�%��:�AYMFU(���R`$8l&�Vw8�*�r�Q���X���x��{��ӶJ��?-v�҅&�O�#�<�s�42���g�j�.˫�s��!A�-t��&�6遲�H�x�l�E�o��/C�T��l��[�F�B�1��S��o�����b�����ߴ_��ŝ/���_��f�'�.� ~����d��-i�E㟫	�U��;b��OX����7P��E)�=Tuz|c��<*'����I�m����@�s���=|z�h�����N�&��n{!��ׯFb��o��O9flr���\��O��l�'�"\��q����jT W6~����;h_ΑBz������3?��1�\��6uH���������>�u���C�\����O�5AT��'kWJ�׾�/ݙX`l��Hc�:��n�Si��Gt	���6zTd�q+�:]�w׉���E�� �g8�7m�U+J}<�лu��o��߶��^�kJ����MG/�5��D�=R9Y�_H�~���!@��!j��OoU
��>b،!��r�6�>P��
�	C.�&1$�%�E�.�q����CH�G�!��m(	�\54��?Ur3��:L`P�b��� k�@��x*�����Ď�jC<Dq'�h�	O��9m���P��}og�@)��O�c�0���FÈ�hv�U���ڭ�����0�_}7�@�~<�u���I�MHy�lk�Y�O�T1Xb�0���<&�s��L��ǮN��b��_�w�bYmQ��%$�s�w�E=_&��b,�T	)�u�>��Qk�@����\d}G�B+3���Y�Kj��!���a���F��XOR���4�5(f�,�S�O;'r��5����᠐w5�h���	��(�W��Ud2r)>I�ssx(GdV��z�T�z�ܩc�,2~n�p�ۂE.ru��`rD�v�����vݢ$u9�!���'#���#I��lȿAЊ���ai��)%�e�.R��߀�'�S��A����-�}��q!/�Ђ�W��_��(W�}���5��o�b��>*�����*GH�'X��#>����P�L8��MXp���q��1�:�b�B�'�!FЪ�D.+E�mD����:3��,�_Fx�8�D�0����)����"�K�`@9Qk�|���d�
+#�i�^���	�Р.
N����X�O�5D��wRZLF���m�|��ӝl�"^�m��+[e?�[Al�P|=�;�$��V� �f��y�!��o�"���%�ʠ�{mYP9"�{�G*�SS���H�2����U��Ƕ���t�[+�F��N9�\Օ��t��'��MA�&Vfd!��Ξ)�1[!��^�g"����_��F����Uڔ_{�����Ì����Z�}a$A��n��7%�b*KG<I��ý�M��Q؈���Ř�ό�В�L��