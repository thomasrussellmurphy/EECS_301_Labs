��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�i��a
Α1S%� �uj?�L�3��TLei-3^5]E�$����/ԄDa�ZO�۩��僧O6䃱Cg�L՟�m�g8v�TSZ�WS��a���j�1��j��,Z����ȭMsW7�wZ1a����FX�T�Ʒ�V�	i��+�@FT�%�������eэ��a�����~L�+80�S�(IFt�ޫc?R���H��TO�{~�\��i�WV�����X�OG8�5��kj��CQ3���VK{��(�u9��ņi�XP��T�dt���RB�h��5xWѷ��{�C�����4��p�g�!g����h�J(~�;��"�5 ��w*'1ޙ`�z䂯��ߩ�X�Cަ&�0���/�W�����]�VlfIbb:�#ƈk���Q�~��%�0����K��{Q�����x{ָ"槅�q�#�p�]zg�D�9ݨ(���w��ߟ�Π��Ll�dAn����wS��+*Z�����(������
��HQޯ��n���݉�R��G��ި��ԟ��GJ��Xr�q,��{� �6�۶w:#��n*�h�j�s�sv�Г':�O���c��Y�T2��a.�=#cD���\+���<)��.�/ͱOnn���> �Ŭn%�J��Y�XF;��ot�u�E-��W��s�{`�����e�i��y�?^6��f�L���m	��U�a�������%xx�9D�.�{����j��^�����&f�q�6�00�}4�e��������&�\������e�ə�S&��G��b&���*�����ųq0�J�r3��o��6g������G#�L7iÐ�	bwx��P�8�0��@�����;����G�X>vap��,�Φa�!��/� T�r�J{?�����
M�F�74�5�=}`j�3"��U{Gm�Jv�|�>50j Μ{ʒ��m�ٿ^��5Xc�ʻ>�_I��7���P['�������0}g�0��Ĉ�Ȭ��h�<��9h� �1�i��'χ�����೴W�p]�L��h!nps��E����`Q��@q�P�����ш�`1�i�>K�
���f�U���F1�i�����"�0�Ǡ�TG��1:�oּ��ԋ�*jpں�?�
|��42:c
��B�i�[�6-���4����q�8:�k3�P�Z0����g	�=�����õ��׿}��}7@in��uj1�E�[O�7����$ ��(g:����p��շ[*T���׵�-�u-!�ÙE��-TW&�|0�k�{x�j���X�)Q)��(3��>Q^�tfg`��A��}	.��K3�1��ҿ�%��|C�5o����1y%�?laRR`���*#�7�-���г3F���(�P���n�pB秹;��Ao}��~e��~�^�D� qV�9q�7�mt�8V��2��|�
�7'9[e5e�}<t�y˛�}�9G19����8������Aǁ�,r����	=�M�r��́ނ�g��kR.�F��������5�3�~�K�q�`s�0L@�]Gd��4����AM��/�e�J�nN�w���o�ҎL�r�B�($���?-@\�
����_^+��ێI��Q[�G8�O�§\,Q��E^�ǇO��L��,�O�^��[e<���!,�����r�&�!J7'>���/�^�!S�ez���w�"�A�b������	I&%@��H��4s���eU��g���!��F�i�;�}U��YC,��MX.�v:�iV�j���G�J[�"��}�Lw,>���gdF�.�xR�؜U�1���ܶ��L�2(�͒�vQ�*D����\�+f�M�T9հ�L��=�Gc*)��~;d��]0�t��b+������\�|�րo�q�2@Cy,��+lt%ؐ�.��U�w\�Zh��ގ��H1��u]�cҞ2��M�K(�Wp�@]zh@���D�5�YħSq�L�uf��m6BwX��22td�49�R>*&�]E}p;�X�r~��U)?�:R1��uVkd:���&����=��ā6��ɳ������PO?�Ъl��p�[G%����E��������2pk����=FMQ�_�8Y�����cC��䔺󈋤���` �F�ize��g��&<��}�~䃡�kζ�Y�@�KG8ޔ%$B�<��C*��������{����l���z;������:����nڞ�*I���m$)4�h_I?;��`P�j����EF�Z��x�e���T�@ ���^)ԛwm����Y1*�vquُ�IZm���"�O�d�O�'g\��`if[�/Be��C�����/3����,�����a>t�XUV�@��A�殮l8�2e5�;�FS	ڜ���f�VSa��]�W�$'y�rW�Vڇ84/=�)��Xp쿦3r3|(1%���@�5h�_����f��|˗����q����*����'%P1Y��s��}�j8��'����k���9�v ��`Rt��,[~���,�7(~ ݸ^�o��E�j���t��{X@}����Lܮ^dr�tXb]����nʕE���%������z_:��@���˰z�}���5����8���&�h��C%Պ�/��&��[8������j���P�)�{�̈�#�k(^�4������8�:��b	��t���tǂW����K���4"�:DAW@���F$,Z���ھ��EvO4��Ց�(LB��6n��l�iK��tzÄ����oJ����2��S�`%��r;,lˀ<�d�)ЃJe
y�A�&#��?9-�/�`�U�Pb�ĭGnT�=b��ҥY�)O�}2��M��Q�k�4����>4FN}�Kf�
ҁ�#�j��+���
��*~��,�`/J�n�����q��A����/{�N>�Ќ&����Џ�8Y�����V�)-͏͎��o17����r0��OG��|�kF9�|O`v�j<'Zu�!�!�aS�Ŀ��뭣�韱h��Ro`��xX�����hؔ�����RE)�A��MĻJ�����I@����h{�6�,	Tɋ�ʀ��/h�P��. �!@�|Ķ�����v嚺��05�޳M���s��P�qBM����M���N/A�ˀZ`^��F�y F�E�_0�v*��1�t/Ǉ];�cNM��r~�+�hK5^���Cи ���B�W����Е��i�V��d�'hIL/28�ѷ�5(�ߡ����sK��G�����%� �9�r�I<� ͺ9Za)���HZ+��+�̧,=͐2,�!i�	n7`<��vy��<�־U;#���9�:������m�� �>0��J@���rJ�bE(w��rH��*��ڼL}���z�2�=���r̡j2�/���Ա'�ZO�����|{��@�x�8�K
���^PA���'����&����a�/�(\���#��l�7��6Bk��Њ�u=�|%��p"D,�q�%�d/Q^*�����\�?FʒP���#J���T���ZlK�K5^Ħ��Z�����S�l�>�{|�ր4P$Xb��2<�� ��S:9��2-��Ӻ"#�n;�X]�ލ}Y'D�'�_�w�A-Q�. ��0���dmC�iF���!�ۮ�b�<����GW;�d���m��L�7�s� !G�"��+@!�����T�0�xmP^�N{���]N���}�H�V+�P,3��2�S�EFJ�|�8�#B�eE���8Lֶ��F�
��{�l43{B�� '�%2"KFK�QA�����7��j�h3�Q��B�nJ����)�M=�pDq�1�]x�&#�w� �FH����Ԥ��{G��7�b����	���ӆ�/�Oo$�|.��D8rK�����_�;�����ݺo��0/�4K٬��6S��DЌ��;Mk�n�àCI4���G�N��g,�R�d��b���؇��g��}���;�y]���Ý��r#��_�TP~.aL}t�������a~�<���M)�|�G)��~��G��&]��ݠʐ\L�{��D0m�LJ8���[Ar�"?-!��q���q�����[#E�����������1%��f|η����epxQ�QW+M�T�EVD;q30��J#3����G
�;�C�e�N��G��P�u~|����ok�%~v����b���SH��S��Ҥa���&���!=�jlHN��(�Sro�V݈Q�V�t�*��<��4�b�G�}��G���#Ib_0��(f>�aE��k�,��>{����g�Twh�c����͇�v���Y�L��a�^M]�ykB%�O[gvBvG{@wV-��%�J^J��Z��W��$�9�|�HBh^�t�S��Y�p#6�+	iFK���QI%�����{(Q ��Eܙ���,D�7+���w{D�d���B�E���2����k��Mn���KZ�`yi����(��qX�m`�;Qi��g� ��wSRR��NK���g��K���j,�Q�p�
.�d�����8�#V���O��VJQ1M��cFǤhGx&�r�fv���f�����!]�:'�p��Ӌ7R��~B+��Gע�yk�&2}��5�[�&L�ϰ�iC�}��Ey��S�hZR���nq� z��%�����p<�~��jă9!g��e˓WI���P��$Y�`2b+��X~؆�pw^p���E��)�Q}���3����XaAi���Q}~Th�e�j���KnO�	��r�y˵��K����H���g���������E���eş��^�]P-~`�C;�����B-�$�<	5۪+�-w���r�����\^��]��gH�g����*ԫpA\P7�:zUWY�+�zUc��w��Dv�1����i�Kt^��r�o	u3����O�pr_�0�)�Ic	+hk����R�_�E����1_Ǆ'���|
!����;��8G��{�vp����,	�1'��u�2�ھ�I*��a�9�6�<*Ix�Dbԥnl��3zՅj��mc�=�D�1CX���"�QA���Ù�������3Tů���btd������۲���+�)hQ�W�z���-�'v��o!gùn��ZTG��0x��^=������S���^X���
e �E'�9�tс.7H��`M����W0yo\��7�]~�<�f5��K�"̤f�q�f��L�w=v���O�iv�~�����o.L�A\�����đ+�Joy\l���s��q��JTV�P�`��O��q��G�2�m��Ư�'�5�|�0� ��fS�uΥ�#?k9�?�o[�
�#	���q��=Mk���SN~ܽ��MGp�K�{@eK����U�FɈ@����q[���0��{���ruǚ��Ln~��+��yI��ĭL���pt�HK�>�|��ч2�xtfU�e&�\�CC@`I�[!^C36���S���dJ��gآ����ڊ5.������W .5B��K��HE��$d\T�I΅�a��8Z�DC���Ĉ�M�B��k��L ��{��6�4��d#Z"wJ�`���yZh��n~��\�=�G W�\i
�-�s����D��48,�������y4�J������"��H{�3�X2���f�6�?�}YQ�8�I��n����Z�+ۈXV:�=�q:u�x��C��,H���xT�o�c��KGJ>5�8�!����-BQ�ƙ!g�kd��f�$�k�o���-7�Z�U�����K��v�#�y����@�pH�8����Su!��K�h�5	�`4�_0�����Ǵ1i�&�E���X��v��l&��>�gA�Q�Dvzt�G�*��]l��Dc��o���t����)�L ����I�]��[ZD�$��n^�$O���(87(t��ib2��3Ȑ�x�]n|���4�_�fZ�Q�t���x�IZ!V�$��:�"-��|>���	��+�㻯�9i'Ul}
mE�J����9՛�Vnx���F`m���a~�?}�J;4�'s���o�K���8��x9��nA���f�%�J�q�|*�(�|h�j9M�G�a�5m�OmQ��?S�@���&�s;^�	��������6�M4ʍ�j&�5!��?Ϗ����/����e��b�h鼈k��T�V��G����.X��91IG��{l�m���p+ j�d�A��"�!���)�iJ��
�������I�
Ȭ�y�zwdM��#Ϛ�����ɏr!^��s�3яz�4-$��h�it�u~q2L�3SC���������{$�2ه�����Ȁ�r��j��~�5�.J���~!ۙ�C�Rl\��tM�F<�%��v��W8������p9�J�o����f]9��PjJT�<�X�jS��p���Ɗ�YӚ�N��^v8��oB��Z�E��f���1�X���!�\ʉ��!��#�x��C���<��G�oj�ʟ�Q�����1�d�QM�W�<��(�FU��n�YO�X2;V�PD��wBe��c�����yVPw��X/��tF�����K��K��N�e'w��?����� ���y���nT���$�R>5�5��/���qH���	Aԯ��3~���sH��F��t#4jR�� p�5"@�c�)&�����N�	9̃.q�o5ʧ%�v��c_�I������Qs�_,Rm��J1!��
X#�jh��b���9x��Ꜿm\
c`}�)V�*���_.�m�u�2d�q�b����}/��� VuZ`QK�	��� �g#YP���~D���K��3z�#��.0�`�F��_����&dr��kW���ݎ�774�׷k�����t����3�]�U�CF��X���*<oS�����]ޡ]\�9�A�GG�+��J�O��CA�t��r�g�U�'{��ŅYT��TQ���!_a�gS�����n��п+��kE��;���"=ީ�p撘�$[B%'6�dN9���ʒ�e�y���i�T>��""��Z��YO��I"�'$��E��%��})fn[*�)��Z�=Jram�M�ދ85hR�p~Y%�39�v |-V\řl��q����+k�
C��3j���@�W��<�(�=����lv��R���o� ��#�/�m��e�^��T�0ڟ����Gׅ�UtA���`	��� ��&W3~M6!2����9�珕rp�/�����;�����ߌ����_`Iz����I�; ʂm)*^�+�ȭ���Ϟ�v}S��*և���� ^��y$`��%�];V��a����F�+E�F@Q^v����~�}0IT��u�l���6� F���{��Š�Cc*W,Gu��ش��ʏ��YT�,_K��'�vC+Zi��0� �M(�U���Be�	��]�ԁ�YP	5u�����Z���г�w�s�o.�u��M�Ǉ!ҧ����������*!�`�C�nǾ���^7W)d�J�2�֝M��l�����O�%������=�R#٫+����Ɓ��t.�����4{U��$&,�$T��KT"�ZaT�j$���M�Sr�_�k�Ov-XƋ��Ż��L��kK�6������\@G���kd6�$�n��c��ƹ�@����/ �!c\vu�"k b�d�(�#�;2��D��nm��=��������-u��B�C�f�%W������8�J9Ӕ­��}U�r곱_0O�=�RH��.��ç"�c�B��S���uJ�^��U�ٸ� �%�`�Q~R��8c��p=��N}��'�{����{!�o����l�M��Tкz��	�Jߛ�vp��_I8�)�	���=��
�����!��X��`ΓP�fX�)�m�$���Ō��w=y(L\H�	~`ظ� {�yϸy}�he��+���+��i��K%�P����/�$��m.�3�SZ���V�6-1���c��kKv�>#���2#1sגּ����(��)d~&�/��ސ��
{M���c���QQ�T��Q%�%�Pg� �"i�����G_<;,�I��O���:Fd�Q���w�@.���v-D`����=uw.\�rی)��{�Ik���GB��'������agG��ETc}?��x��35��]�5���qU�g1�m*ԗx)X��}�1f7]��F���-�.���?K  ����&�Lp�ٟ�Ê�G�?A����	.�A۟�q�X�` ����oF�E��n�c�k����N�F�'&�&r���2�]� �t��^Z�7�*�$�bJA���� ���[	-*n����wR�5���I�8��Q�|F�-/�둿=����	.��%��yhgz�q-,�Mga��է-� r��w�6�D��c��s�����8hx6V�pə�;�|�G�)�pԑ���3
�	��vWM$�̿\if�t,�dCfQY��g$We��n����F2��qadqu��Ү'w4����r�&^�}E&R��5J��o5$��z��99�sX
Q�X�5sQhȳIVXOHE����r���>7�7����m�����_[r���~�����AڧL�N���e��ß-�u���z�e}c��i6�Vb�����sI�B��G����D��|��0���̑��m;xV��Mw���&���&�;�-���W4C�}���>D�ǔ�	�z3k׻�7�֡�|�c� ���z9��J0�H���][��WgC-��ZN�w5��^&�m�� ��ۜ��0���U������*s#$�;�K�����O��u�D�~2�=��gy{A6��(�&aQT�o�,��O��L\]����I&�u�B�	.beF���W>�7�)�}��U�>�|�F�%#W��K@�X�4��#"�+��M(�@C�spX��@���6���������Z�,���_m�E���<�5��� �WafL���,��3��Ν�����Q��9P����pX=��t���0�
�iˈ6��s��� ��C�p�֪�@u'�X��(�dA��"R����/PN?�{���{-�-��0Dh߱1ٷZ�N?�`�`= �0{ޔ��m�r�J:70s4&KY���xށ�JS��eܪXa���MQ�:�m;B2#|�^���c���w�� ����j��t��݁�<�G�\x��ZqT��v@=�Ê�.�A�BfQ䳳�\8�������e�ݨ߷-d�����i�`Vu_�Q�o攻<X�����9<�T*�-��تR�ɑT�	cBN��~�����HJm�cѭ�����{�s�����˾P�'�C&�i���/�=j��2������%3�5Lv��ׄ�-b*eѪ��-��i�?�>1�r;������:˗*��c���,���~I�f,@@�$<��
P����R�.����Q�����D��Nnx�22Ϩ�'�G"��q7���6���7�ER��v���i�CF�&#b��k6����<#ö�4� �{1�KS�պ��Dw6��<@�VL�3oj����O��z?S����ЈCC�c��h����Z�UR̥�Y�)��d�Ë�����m�H����	��N���ͤ�8.���边�:����5�	g(�=(W 5��_>���Dz���9
��#�,�O���S%�%K�"G���5�d�Y�Tg{Is�<5����kt�̎��ұ@))�/���*jI�zQ�	w
���,��|�ǒ0,��%�x�Y�@*?��w�:���M��h0���iU�`%��@�%&V3��۝�:\�G��~K'�p;aL�(,���er2�>�%!C������~6K:�p�r��q��`}��!�y[���O?5B��nmt�����e"��0�����LEX�bn\g�K`�g�1nL����|՛��a���Q�������j(�v��6G�GBG���(�̬}�="�Ν���%U������F�ojދ5BI+�uI�T�s����� ?P}Z��W	zV���Q�4�}�|�%��L�"���1V�d
������p�Ûd��c�,��O���h^���!����YU-V\>�������0�I��n�Fb+N/J��'v~�*�(ʯ	C9$��o�ed�"��a��* ��cP�Y`,T�B9����	�I�@c�A�����ZT��uub��t�qOqP���4;iP�W-lؓed�x>z�d'q0�1>��_�� Wb�����Ĵ�ҽ*a���<��
^)�	U�:19��8e>0�w�}&�JP���\IF!.�����7�1�ԢJ�%UW�Zg�����)�7aR�_z��:"]�xh8ѧ3Q����l��Mu�E���l�Mg\���2iLrN�<�@<�޶�g{3���?�=P���9����ޖ�0֦��ʕ�ݼ�R1y����U���z\�Zfև�X�H����_�AGkHg��	��d�n�b8��\D^2f\?+�p2�UI��i��]钛;���1����I���q�K��6�Y6h�$���6pߪ'���?�Ԍā�KYz!��p��x�?��5ـ�6?�������Rg��nIw0����2w�,����,�.*ئϯ.��/�^��x�b��)�q��R%ȟ����0�_4�E���p�v��0��]���j�L��q/�� �'��������5m��g��Y(hA������K=I)r�У��ׅwW���ud%����$�u`c��(�kݙ�ꎡ�!p��s��В�^�{�Fb�mA��Ѫ�uJ4ƌUo��<�8��q�$=cA�p�}�nd�V�U���� b���8,��]S(ѓ#'%��je�ToҦ=��A̔�7�F~g��tm��5��,׍�������o�o!���P�D}���ln����×� dU��ާ�/�b�����ǟv���.���:��������[� S����;��WP���~{7����UE�G�b�#WY��M����fZ���`\�ѦG��!�8���S `}TN,&Pc�;y�v���:c����bU��SvO��H.ȍ��g�s��N94R��"�V$�i����w#(���M�Ѽ���Z�(	\�|�E��D`�f��[�N�Z�Ab�>��&���T�����X�Qj�
�T���1#�Ap���93� �����1�^�����j���]-�g�g�?t�� Re4ĲD��ի�O����#���������"B�6\xZI�TB��eĔ��Nn��欜.��{S`�*�[�bzo��TR���xES/�g �o$�k��[Yta���g??{�� \;�+J���O.#5�ܰ� 6-��2�����q�Xf�	�Q��l�F� w��J"),x��G�P�P�f�6 x�y�; ��v�
�88$'w?�HFF�6�Rly�Q����߷�KB�� bb�:�ߴ���Aj^����W6���~d���/d�)��R�Iө�I���$L�W�B���Q�zrof��m�Q�C�0��b��,�g^#�g��0�'m?���q^M�4E�o��G�C��\�)ΙD�`��8E&���D��^i���p����*�;�w�dI�0�Y�qt�SP�	��N&��2^pƑ�C���]�yS �8�B����t:��ϕ����Ҽ�w��'p�f��r�(J�7������'תU�L(ϻ���:�"�QMI�h�F�3*����.�C(���p�@n���8&IB�M`�����j-4,lH��*"s�������v�֪��w�E;]�A5A�N;��M�ЫyӴK��;�<c'$�Do��wps�����+��F8B9�o!�0X�g�&Z ![�ـ��	�����|.>#��
8��#��D@+�!aٵ=��0�>Ѝ�imM#���\��w!V��`�ܰ@����K����D�����if��X{���?�)���˽#��A�bw�̆�J�\�"�2u�7$Ds�
�w=�w��&2��U�O�#��a0輩R@�˖�+�Z�����Hpˠ�������s(��}%�Pi����RΫ����4���M�9��8o
s�������`%��E߾}�'g����,���f�,��o%D$��\�L{�@���������Z�����M�:8U㢝��Y��l���8�j)��]�^����h�E�6�;o����K��ڄ
:�������8���[�{,��|��a��c(���)+X��.�|޾G�
�y�W@L#�M�O�U�M���؍p2�����X M%f{w�9����f�X�9�
��!�3fh�5�j(Ɖ�s1����I������ƷZ��\�����9p�N�Ӎ�[��C��j
��.}�>���������3ם�dM7�[J�gi�_�:�8��)~|p�Ý��T.qn��|j&~�7z�*:T�UG�ե��b8u����EpG�����o��m+vq����bܸ1��B�s&w@j}�e�*�zjZk.�w�]d��3&�%fs�ZI�;�E#>�v��ӫ�}Ʒ�����x`*B��^�}�<dw?r[�c��h�p����Ò�z�%��D[6���}����_�7SѲGĬ�^�/� %�ս���]&G�F����"~��X}M�
�bpf���q3��&�c�߂�[0�R4�#�F�ُfW�(�^� ~���JJ�廿!=^@���^􂗞?��ahL�2=�[ɚ[p"�������M�KS�k0;e��%-�� %��P����C�>��|�9�+ё]�l��<)�!4���x9������C!a�;h~_�/�	�m��@%�/�`MG�٨|� A���������B	
F^f� ��F�?�>�*���oϚCUR���K�4o�󐇋���~������K~�_��Z�
����k������l	T�j'���SE1��a����V� �.�KV���������ӳ�_�.ݰ��1(d)��.��� �X�m0��7-��Q�tG��`wz�A�sQĎ%��N����^�c-��,|&땠1��\[��e�_��<g)�K�4q��⌆]���I�ą�Ia��^�Ґ��9�2/�F8N�(�� ������T58>0�$]M�>�ƈ���t�d:�F�ۄu
�3w7S;�z^��i��(��ÎU9�}J���bht��N
^�6.g�%e��X9d�d���!�Mb�i⼃[ͩuI�K&�TBy��yfY���v��f2qH!=)ES�,~�mtzCϧk�|gd�RWcِdf}ѵUu��H���}p��8��q�Xz��=
��Gu�Q�Ju�[{<ȭ�<� {"�.�"P�NӲ��4�� (�b塐��O�Jő��8�|P{��ՙ|o���g$9�0����ui犞-�#�/����3Ms�3X��j���;����U"�Ϳ��g�n�Yyk���gĥ�� uα��	�fA���l��?id�v�<�!���u��)��x��E���#d�Zz��A8_)s�P-'Sa�ŧρ�m������}�K�l�/5���eƽ���)*�Q��!;��rA�bm:����ғg�����֫�ѥ��b	 ��+�0M��5gg����qU]��]ZҾ+{P��t7�G]���E�`�����|�u\,�;n��(ľT��9���+,��p�.�0�����#w�l�{��z�#ر�
�GWВ�؆��@�"�$z��'����g�=�e�`w´�b��ߦ�PU��u3K l;�Y�����J��v��+b�&4}�� �P}:rGm�L��A��*
���Ci�i�;F(9i�G���Z�Y�{�_�j�1*������ټ�:�7�Q
�FJ��{�����Uu�(H���[�ƈJ��-�,,7�߄�6��pF:�� oz�oyu�/�A ����U���ø��fB�����ؕ)�*y}�0B����/C������D;�˘���H&�.�v�d(��M�p0��9̃��s���[zQ6z����b+�Ȏ��jO��[�]�BLM����.תҝ��Y�5I�A��ћy�8�Y'c�_>P �8q��3�do�����"�\�����Y�R1�4�p�K:���,`Ny�ff`�[��R0�C�Ԉ�ّ��)|��<w
_je�z�X�Hƞ��pԢ,"����Z���k������!S���	�QF�뫎k����(�%,\Z��6�Fx��z��ή�A��� �q�p���=�N���{R`���CW��+���V
TQ_ޙGE���f����[6*Ϟ�s�V�.O�K�\S�0Tè�;�KP�d)�ݙ^E�.������-R q�W��
[�2͹X?N��z�������#��B�W��`��á���}ս]n��<��A��n��,/<k��k�!��q�0��*��#�;Mt�X;�9�`�S)���.���~��@i��&�y���0��Agc��#̧�y�2Ay����NiM�P}�1�]�+Uш���m{	:������u����S��#�35
��ި��h����&0������8�a,�_溹�e��&ϕ�5F�D[\��	�Y�&�(B��k�!-����G��!�}�S.Pk'��ƛo&�;[ z�O�65��\�~{}.�a��P�������<*���WG���c�-Gf���)`Ÿ�On9bt8%=..��Q�Đ�f�SAt�J�x��]i�tD�&�����}���:�D$@v}/��iI��t�v�%m2lB��Q��n��m���N/��׾E�,�3j���Q��� ?��O��N��_�r�48^@����2X6E�D��?�g�Ê^����9�������N�j�sXPQ2�R�b!��
)c��b�K���S�ev'-��Q'�[�uk|��>?� C�U7Z�� ��o"�nQ��Ҳ��,��jɚg脒X,Qb��u%�1D�I4�� j�$ͻ��E�N�����wcb����y.2JZ��,E�q~�3�l�د%HX?����h9`$�ĳS�	�]�}{�1,��펨<�.����k#�50o�	;K�
s�������J��F���q�g��e+�9�9WP��7�r"���az�/�j��O;?�1>��[}��\�8K3-FJp9y�Hl#�dP�UbL��;#�rf(6^��/f�z�0x�A���~��m��w���kɧ	Z_�گ�QB�f�����Hǵ��f8������}(�$Y/t���O��T�I(�u��~���l�
r~�������������-��O������|�?G+����'[O��f/���W�b@��-+�`�H�<`E+���:K��k�̒���鸷E#ĝj6��/N�ғ\�6/�I�X��!79���ss�l%�r�p�R.yQ�k�����1��g͆0�{�L�JۣiC�fbź� ��(��	X�{���,�U}t��{m3��3<#��
�O���
C����	�(tp�|�${��<s�2{��_�?UwK7:/k
(�]��AwK�ɢ?��[�N��`Ǖ#H�'��J��) ��qy�_/���iΩ*f�!���!��b�K����;�y@��Ŵ
���D�Z洒��U��qX�S���n�M�wß���V�����9����%��Q.�a<vO1I� E�^����H���7��6 �7��j�����形ބ�S���l�����@�[�J�$t>&���6蟽'f���dH�~��C=T,�@nŵ�ޯ[�ƅ���-|�@0I>g!�/nA��]��"��vI���2	Ba;�}:|-�vt�A�.��墊5��"=	z׽lC�&���t�J��rd0A��ybr�AL�ͅ�n��i������2��v�5��+����)���~Ʋ����nS;e�y�%G"Q�����.K��-�>��4�[�v���7��${���5�̕��e�jx��x�����N�?��Z#��;��Le=����$O���=_�B��[G����b��D��Eb7�x(ǌ�W����e2�}����O��f��k	����R��Z����F�[�h�S�&A� �M���ٸ�A?c�bH��=XS2%��j����[��Wb��7�o�y�ݰI$JH��yat9��l����*ᯔ�זr��E��	T.v��˖ȍ���{j��z�Y�-�Հf͛���l40e�q9�6q��	c��h�;��;~$�K����J��)�v�̨ �gS��tX��
�G,�S��a<H���g�T���,��v���;���>��&R�B��W��A�g2:�&�X�[i���u(��[����B�J���tԅ(����z�������ϣ�߮U�I��]���4~_��O���� ��@�ҍ������b�?���"�Շ룇�����~)�ʝ�b�A�]W�^-�=�c�|��6�V�9�'�z*��������/k&�
AX�[��&�ʔ-
�άx�Vl�t�$s��e�[���/�yN����B?�aI���>(�
�4l)2�lPr��p)%R�'/��A�e9�W�O�_�������s] �P3)�H�B�;(^U?�wc
@n]���L?�2�vMA��v��Y�Ⱥ���U�"���MJ
B��#���ԝ�]�dx�H��u#;$�U=�4�3�8@'o�ӵS� ����J�c�������OKiRƅ�TA��ʤS4��4鱑2������<�r��V����Ya,����|CN?W�-�N~Ue�e��k�"T�路�a���w��'��ID����3���g �џ�<�0���4�=���K�ۑ��������m���
dU��kW8�1΃��j��8aǞ\b���hk��u�zU˩V��I ׮��Ύ�%�	dJeL���~��-�G���
��ߡ���)���`�]��2����'�#����w�k���dQ�?|3(��MH�Oj�3Z=�Eb�`^y��*��<�nhD7�ji�<�pù��֪�R0�aP�R�i���^;�S�����x�2˺��O	~����%���o��W���M��ZT_���O˔({��hj�O�B�d�,I��D�sX�Æ�@K��i�}���Y��נ���E�P�����幩
B��}*!�Έ�
Q�_/ߋ�hm�oQ�*���	3�D���&����j}���H����[;�`;��`{	+s&憺���Ln)�H�*EH�
|�];�M�5�����CL�,��ڗ1��W����8GC���^�7�WEd4����0N�0�f�W%�K40�h���^�3d��	�{�j��0�`z�&��6�<)q�pu�z������t�)�~�J�.`vJ�\� �N��5EgO��'��S���yy\��l�a�\��$|�g�:�r��p~�$K���������A=��Ob��[��!��:[� ����4K��G�	��+?B*�J��;�K=�[���V�TSZ��b����Z�����d;�Ne�1�q\e��̶m�T>u(��܂���Z��̸�xH���/�-�R�I��}!7����$�tr�j���T^�����A���	C� ��ѽ�����x�׶��E�������z�vk�E�N���f�M��zU
2�v��<Q�����l\o�xGvk�{�T�^�%iF��s��|�Y�f<	oHw���R����Ar\|�Ʋ1A{�4s�^�|�ã�ZF�dq�^r'S�D�X�����R_�{J�l��`P���w�1z��U�	��3�4���*T�V"J��N�|�z�6�|����
�=� �nt�+J@@���
�z�����������#�,�/dK��wlN����t�1Ϲs?N�V��i��sb,[(0�8�`T%!]銘�V,=9�����&6.Y�a|Kqc��y���z_IEW�(������UV��a��I�)�D&%I��A��f�4J2�f�%������J�{D3�{�(���ȣR���-A�������4}̓��y�����M�H�����vM��WJ�]�t�fm���y`/�Df]���gRL�Eل�ln\�w�;c�8'ra�)��,�k݀��w;L ���&#kX� e����S�^�E�����4>o�d���qW1<�v�d���&���0svd�G�Ct��hX�v7$�)���Gs����Ť��w����#0��M�!me?���%Q�k}��0�`,�[q 
�0��Z;Bu��zʨ�#r�N�������4y1��t��H}ұ�y>��|Ǚl��j�X?,��<�e�ܬ����x� �O7��P�2�sť}����W��x����	/���˨,-���C'C�,щ����z��ԼQu�p�����tr>4ߎDHh�ȳu�� [g
�}i��8E���g�%��кW���>:L�:G��em xxt�+�u�$�ڀ;RJ&"p���$����	�W��P^Vϰ���^���^��6��ǻ3F�sp�7�LZc E~�8�7�R���������~��_�`�d�Dp��Gu5ܴ�PL|�k�����x���|�#d
N�����J�/:!�y��8`�#�A��Pg<�Z�tP��m��Eƛlc`�H�T}[���<E��8�J�O�Y�a�-�'ɭ|��<֎[��6��Xj.�`�@�^٣���V툱4���΃N�ݘ���L1 3����[(O��>`0?N�AE�o0��9��x����ݘ(`F��9�]xr�wK_$�RHɸ�