��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\���V�fnvx��ÍG_;�ȅe�~�>���9�>��Y;�0GP�5������~	D}��tx��i�0*� y��j����{��5~xf�2Zs��Z��ܣW�S�1�JFJ�ջ�8#PI�W���k�<��R>.-����:6�<0SÜ&�n��)�*tG����g�5�NC�me�)���|O��χ�>��>O����K�ʚ�̞�I.�T4Ht�*x�X�=����O���\T	���:��:��_��_f� a�!d����̉]b:�_��肩�@�MǠJvI�Vj�����4�2m=��]"��&G��T��Y��<����}A����c�^ GT'j*Ph���XflЮpח���P�b(�?��(�]������{�3�PLw�����H���G6�В�)���K��}�����A����&�Ȓu}����y�)����u>�'�]��-$jmƘv��Ъ��\��:s|j%�sޘK��Zl-�����A���n.�6}"��@%��]��m#����� j(�z�����7�:1x���(�r�xP"�V-M_�U�D77?��;lBK�|������mп)8�����qg�l�E)h�%������ڢ��M	t���M��*�t�����/�o- ��ú�ҙ�{�*��rׇ��ܚ�>�O�i/� �ĸ��kl����$P���$x�8�򞧇��^;K$`�?U�z�"����1u�Z&��5�)jd����f��}��xGZx̟��A�^<�gl����ݱ���2�	H��d�-Y�zs]K�}�]x���Lӳ�L����p0�8��ȼ\��J�[���g�C�ѡ�G,,|�W�@ʭ�Eǿ��#��{��cׇy"u��0'�~��pT�S��i�:����0I	.��M~��5�g�b�,:j���S'��]^t�ʜ���\���ت����]���HH&JN;��0�@�0����Ɛ(�&B�t���rn��7�f9��+%3,��i �8C��cs����"�ɮ���=W�'�]��*��?ﾯ~<=4���+�"����
���Z���"y:$�?8b�m���M�D�x,e��F!�bWxXL���K>��E
�o떲��k/��_���D����l�S�����C�2����1��(��������tsL�%|!�_��4��R��b�(���(6B�����E������u�"��$�!É��E���2�g���P�I�=D��{�Oa(_��G��ח3~��e~���c��]/`DU� 4�I��������#+o֏Iw���8+�3�-��4Dn�X�P���ǫ8fӒ+X=Τ��Wdv�}��2<��{2����F�:.�o�"�p���p� v���^%}�ս�=��y/�GbAѭ	���k�TGM0F���c��u&�il0=�X��`1;��^�N�@t������7�W�%ٟ�3E��`�EY��!鼰=o�Yl���N��ʺ��/�s+|�*��G���'��8MuZ�^� ��X)o�;4�2�7�\o��o,��#��M*��\/c��E������@KRt����ϑl4�y�*����	��(_�=J7�8!_qPSs�ҲNUXr��F��{	��u{멅��i����Ɔﮣ�����Zyl�����.��׽Dz��7��|kː�Uo�P*���og��5*w?�w\rQ�LdmB����h�a�X�t^�� ��N�99ܜ�	q�gZ)���Sĳc��(�m`M�J/RA�5��� k�3��<����vB!���xח�o�v�!��b�����Q��c�p��j�z���dff�ì��_��T��`S�~���7��G��K����H��� ���$[��3 EV�I.�ت�qC���u�f>$"��J�L�]GjeC���ќ����C��\*Z?����|o�H�b�r�t{M,���)����i�t�m��IPkL�Um��5(�R�[|�W�{��]v*T-�4;�����s{>6XK��Pȭ���2u��dhϬ[���Ff�����v�����nz��Ԓ�m����6yj���4�$�\��w7"�"6�w����&Q��X�]�^~�/g���7TzU��߶A0��N#]cJ�N��������o��Le�ǜ��t�!�WK�n|� � � ��;�-W*�g����!tw|� <%B�1�J��P�w��Mu^2V�����#sr$_P�Q��%�s�Ƶ-�f)��İI�YG������Pj���ţG��tkkt��fSr$A�c�8�j����
yZ��:s8�
;�b�p��_[G[�{2����['iS��f��yP�wb�xiٵ��1B�T-=Mr�=aU��ն^��7�'���r�2��0�[&��V ���v�h"Š���������81{H{������KQ�O�'oc�y��0Ơ���qj��|����%c�P�BXz 2�2���o	�:�A:(�����d�oe����yl�C��(mƋ��8u&�oaȬ+y�&�B����ٔ��|��G^�����ݟںw�#S������[.t>��ueŊ��:�!���(�y+�������d?Ѿ��Z�}�����Qv]Ʌ�n�<��IH��XbM���gX�6 �<˶�n� u׉�+��F����G�5�^R����Q�k�´^���)0Ʌ�iS�����\�ӥNM�Ƥ�Mh��E�/�*��4X�d��K�O��+Z}�N�׺Tz��L{$�B��{���%�r$�.-�Y����Ty9�u�@�!돍����o5����O�O5o ˛F"e����9����!��>\_� &T��2:X	8B]!a�+�u�(�U�J��]��p.SWA�>e�k 6��u�/�O�FR�_�F�DQ/J�%J��D�e�Ztk�;�0b��XN���rуk]����T�����Mͭ�\�lx�X��,���"�mm��o`*y~��Rx�0p�Z�7=-���ʹό>�>���U`�\S_�R�f-��뷱�C^�$���#0������A��PSR0,�J)�[@��c�R��oj}��7Uq�oLa����X�P�]�-|:
z��)��Y��tDY�L����7��uk�L/��n{s�.�/W�w��;�_�Ϣ��^Xk�t�o�M𸭂U��e$���P�!�O���l�~C���c*R�i=2C���98G`�y���p�v�B�5�&QyJ�U������!��y�g���}�wXN�:4^%o�ܬ�+�0�.6y�9�VT0\AJ�n.���u��q>����U�H,�jT�Ů�%V��@GX���ב7��LAq!� �V���1�b����':���C/�����@��߯Qߥ>���&�W!�;���4K:^�+���+nY���'(�o,�cے��I-�.(C�@�}u��\����
����h<+��]&u3��R���ȸ�LB�.�۬��w�YX�e^?0����L�d|�M��#��um��XHTnX6�w�!a�*�57(�?֐e�5I[��Wv��i�Ht?�^V�ِ!S�>�̫��}���Y��^H*��:�e%D	����2���(��j�����W~�fʎ_��G��i���\�+my�[,�@�C|>���sB�ʀU��%��a��O�S�a`q`*g�N�Xˬ �ٗ��n��ű4����r���̸�ȯ�y�؇�P���"a�;�~ٸ̞!"��`�BY(�	��pC��L kg�=���r�)x���u�|t�*�޶�����3mH8�ط'jx.���ƷK9��+���a�J��c;1�35k��m+�}��*�:��z7�1Jl��ޯ �ƃ��"N*R�GĲ���	y!���̙	����� �*�Xp4/��y9~2��r'�̪�g�xJ �B�(ꬴT\LW�
r�g��39��Uz�j�b{q����2I�-}劆�r<���#��:N݅t�m�o�F� 6�L��'a���8��׍K^��U��g�h�`ttS��:Eq���j�A�.��7[�l�e�b��$1-�I��M�M�}��o)��d�%����2��k ��u*����*N0�aX�v].��.i����Ǟ�;ё.���_�����8���!�Ī���-Ă����oRj��ܓ��L4�ģ�=����?*��TA��ky�n�n^
�� �U���4(�c����?b3�'#	�m���Wv�����u�ݟ����"|&���p`\ck��O��D+�y?65P6ÀW��a���X�z�@��� ]��g��8��Ǻ*$H�ӋM�c�޶c�b����<��3h3�vP��[K��z�eW�{�(�K��WבYRCtJ�p�_������}H���#�{Ө@%|"f��t��M�cr�3�z]YTOt�<�O�#sX��Y�͹{�q���d��45�M<��wU�X�F�9l��~�����L���d��S�Z!'����x��|�9_���瘣 �g!�4v���$�������>��t0t�I34�'�0X��D�����+�Ys����������r"�,�-�\4.͇�����?�-h�M�^�վ���?�74�a~�}{ek(�Ƌ,��׼C�2��r]��94m�|��8��]0�^5!�P�8���ӷϹ��-��]?@Ҟ΃Jq���A��e��ƲG�=tt�u@=4��<�w�<�s¬ðG��]�X���^Z���,m�E�� �%������U�Bd@OE?>]ta�(���GcϢ�9�aG2|cӏ蠔M���y��ԁĘ�����˄��sdh����vHsy��S�x�?�\=�8j�vu���#���"����o<�V�oo4hJF,w�H+U�5c����'5
^|8HH]�(p�&?@kvv{�b9�^�|)��T8S{ewD��e�����6y�'�S����`ĸWp��\�{)0_���7$�!g�RZ����������R�|Ϧ�!.g��1r��d�~�*��fB���kv�;!j�ǿ��#XJ���$��������_�0��90�(���s�s=���J^�MO芓-�.r���h���`��A'[?��*O�Q��8ږЕ��]�~����(�����G�z=.6s�d₳��>��/r\��RΪ�wN�;���1M�I�5�x�u)7j+&���w����lM愅R��MnR���h�����W#њ;���~��6}�|I��Eʅ��;j��m��/N\���l��V�A�� )@w(�
�K�c�9�G��/3%Ƽ���g�~�^ �m��PƧ#�
���L����_��}�������}�:�sF}��t|i�G���bF��J�8T	,���+6#>��;Q�5��,V]����̶�����S�Q���([�v4����T�o�ns|:��g�4�� ���|i�}��{����B]�R9��r,9^'��F��$��PΆ94�X�����w���n�))p����7����R��r�W����T4^0�Bg�AKX肐~��P��oeĪ%V�4��~$$�I}�!���$&�M�Pf��R��>������0 %���ɵ<�`�:�a�z�Y�����%2Aſ2���<��^�d 6K<j��E��YL�l�=~\Fq����,4���Ϸh\k!��N�8����������;#��(����44�d�)Yŷ,�M�Q"�^�$�S��=��(�����4��<���'`w77u�/-��](9NER1�0C��ǔH��� �%�3mB�{&�O>�w^Z?�L�B��8�h�}|%o�}(�`Է� ͒��o�=/F0r�	M;����pr[��J�A���+9fx��tQ��*)�Ӱ��$	����$+)�Y��.�!b͉�]�}=���Y��.\���uI>wtL�L�n��mi�n'pbj�����z~���
bt&K.Nt�o�Sj��ɯPe�^�@��hS<ͥ�a��gU�
۟,&�˖Q0D�@ �=������,z��j)s��V�Bn��Ӗ-4I�8��Q9���ck�$@���D=Wt~��2�!h��cR'l"�*��q�_�� �F���P&�F�C_v��[.����i����}%C�v�%�v���
=���fm�I�x�Li��4�QR�N�Șd'���}e õI��c��j4]�D:aq�P2�2u�(2<��s�n��KYsl�`N�����s���iEBj�ɺ/"\��*�7�����0����U��u��{UP����C���:�@��/�o�¼ߡWz���*<�z��$��Xvt�]�) �5�v�*�W��B�>�����a^N�i��Y�z(/��I��d5ԅ��$�9̛D۰�7~��b�L�Zd���H=,��햫Uv�s���]��K}k �t�Drp`��\؃���I�a$��f]�䅎_�B=�#O��Ug�*'��"�y�1��E9��{[X��$�t����R�F���
ʙ!\�9�ڸ�=0#�
?Fq�A䱋f1�)�N����ZX&�Q����Vt�d�N�Oٙ��/��H �
&��%���QH�y~#�֘���ۊ�6�Z��%%�4�$�m�e��΂qb���R4�V$�[�L)�]u������kL�o�V�֪�
��_* ��
�j
�ơ8���6�Wv5Ab�������P�4��R�fXh��d�V�.�l�?>/�zq�Z_����,�A"<h�*�h-'�Y~٦�p0G�Y�._);��A.��+����~	��Z�ڤE�?y^�uޭ&�l�!94%#�&�=�h�&�������gG']V�a0�^=v}�<�����l@>]ݗ��EUoDT�Aq,��C�w�p�ֵFW�^������a@)mn=�L��L�|G��_������o�I��ã�N�������������h��5�	+�-xFx0�3���g����w�Q���E�0g0W�b�z��o���g�`[��Jt��;K��Oy#B�s���־�&��k{���|���^'�'e�.g�F����à��Vk��f���哳���ܭ� b�a����/��'3����{P��=�^먋���mk���]�}�5��ǉ��餉W�2�K:�����("�$�����b�W+���9+h{8��t������^OS�<*�����PR��<.���ӏݬ_o�#�\B����8����wH�5N�)���m=�AEa��`~CU�*UЧ�l܁!�9����ik���9��DW"��s�"�����47�T�A%��)|xo��S��@�qQh`�r�q+LQ�@e��;�;�C?8O�n"���T�S�hVD���(��Km��P�ެ�,��~�x��?���H���Z�J`��\���v�AM�p��F�?E�=4e�����~�K��p�B���� O��8��j�Ea�D��-sm�1�(Ѣ,� O��:�uT|5/�9���!�<����a�(PP�Ǭ�"�Ɗ��r��Cָ�Y3��Wgbn�k��dW<����#+g�7��ېї��~+�� Q��ʸ��7CRܞe��9��NT�K=�XSJ��~=�1ê���:zU�yR�A��`�i͞5��M`e�~�2Ϩ�F5�����vD�g�[-�n�1�f�!�-՜��.�>T�sgG�9�Tt���X�7e�J4����_3�Ƞd���c7N�B��%�ȋ��6������=�μ�0�������cWQ�������(���#<J���<e����#�[7
�;o>Fx�b�Y��w)�n���$^6�4j~g�c	�6�>�׀8����r�p�J�4	��ud�`C���
�ѥ�8}��:ݬ���X�d҈��;-e>��l�����o�CZBً���'��X⥃��!��[�|nD�V�g�;�v��)L54'Oo�;Ňd�xq}=ۅ��ٸ)@���>0>RJo�"�ƻ�Ĳ�I:ƌ��:C���P����b
;ͽ*�N/'#J�%���i��&G �;��]�����&�/�W�������M� P���^����