// megafunction wizard: %ALTPLL%VBB%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: altpll

// ============================================================
// File Name: pll_sdram.v
// Megafunction Name(s):
// 			altpll
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 13.1.1 Build 166 11/26/2013 SJ Full Version
// ************************************************************

//Copyright (C) 1991-2013 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions
//and other software and tools, and its AMPP partner logic
//functions, and any output files from any of the foregoing
//(including device programming or simulation files), and any
//associated documentation or information are expressly subject
//to the terms and conditions of the Altera Program License
//Subscription Agreement, Altera MegaCore Function License
//Agreement, or other applicable license agreement, including,
//without limitation, that your use is for the sole purpose of
//programming logic devices manufactured by Altera and sold by
//Altera or its authorized distributors.  Please refer to the
//applicable agreement for further details.

module pll_sdram (
           areset,
           inclk0,
           c0,
           c1,
           locked );

input	areset;
input	inclk0;
output	c0;
output	c1;
output	locked;
`ifndef ALTERA_RESERVED_QIS
        // synopsys translate_off
`endif
        tri0	areset;
`ifndef ALTERA_RESERVED_QIS
        // synopsys translate_on
`endif

        endmodule

        // ============================================================
        // CNX file retrieval info
        // ============================================================
        // Retrieval info: PRIVATE: ACTIVECLK_CHECK STRING "0"
        // Retrieval info: PRIVATE: BANDWIDTH STRING "1.000"
        // Retrieval info: PRIVATE: BANDWIDTH_FEATURE_ENABLED STRING "1"
        // Retrieval info: PRIVATE: BANDWIDTH_FREQ_UNIT STRING "MHz"
        // Retrieval info: PRIVATE: BANDWIDTH_PRESET STRING "Low"
        // Retrieval info: PRIVATE: BANDWIDTH_USE_AUTO STRING "1"
        // Retrieval info: PRIVATE: BANDWIDTH_USE_PRESET STRING "0"
        // Retrieval info: PRIVATE: CLKBAD_SWITCHOVER_CHECK STRING "0"
        // Retrieval info: PRIVATE: CLKLOSS_CHECK STRING "0"
        // Retrieval info: PRIVATE: CLKSWITCH_CHECK STRING "0"
        // Retrieval info: PRIVATE: CNX_NO_COMPENSATE_RADIO STRING "0"
        // Retrieval info: PRIVATE: CREATE_CLKBAD_CHECK STRING "0"
        // Retrieval info: PRIVATE: CREATE_INCLK1_CHECK STRING "0"
        // Retrieval info: PRIVATE: CUR_DEDICATED_CLK STRING "c0"
        // Retrieval info: PRIVATE: CUR_FBIN_CLK STRING "c0"
        // Retrieval info: PRIVATE: DEVICE_SPEED_GRADE STRING "6"
        // Retrieval info: PRIVATE: DIV_FACTOR0 NUMERIC "3"
        // Retrieval info: PRIVATE: DIV_FACTOR1 NUMERIC "3"
        // Retrieval info: PRIVATE: DUTY_CYCLE0 STRING "50.00000000"
        // Retrieval info: PRIVATE: DUTY_CYCLE1 STRING "50.00000000"
        // Retrieval info: PRIVATE: EFF_OUTPUT_FREQ_VALUE0 STRING "133.333328"
        // Retrieval info: PRIVATE: EFF_OUTPUT_FREQ_VALUE1 STRING "133.333328"
        // Retrieval info: PRIVATE: EXPLICIT_SWITCHOVER_COUNTER STRING "0"
        // Retrieval info: PRIVATE: EXT_FEEDBACK_RADIO STRING "0"
        // Retrieval info: PRIVATE: GLOCKED_COUNTER_EDIT_CHANGED STRING "1"
        // Retrieval info: PRIVATE: GLOCKED_FEATURE_ENABLED STRING "0"
        // Retrieval info: PRIVATE: GLOCKED_MODE_CHECK STRING "0"
        // Retrieval info: PRIVATE: GLOCK_COUNTER_EDIT NUMERIC "1048575"
        // Retrieval info: PRIVATE: HAS_MANUAL_SWITCHOVER STRING "1"
        // Retrieval info: PRIVATE: INCLK0_FREQ_EDIT STRING "50.000"
        // Retrieval info: PRIVATE: INCLK0_FREQ_UNIT_COMBO STRING "MHz"
        // Retrieval info: PRIVATE: INCLK1_FREQ_EDIT STRING "100.000"
        // Retrieval info: PRIVATE: INCLK1_FREQ_EDIT_CHANGED STRING "1"
        // Retrieval info: PRIVATE: INCLK1_FREQ_UNIT_CHANGED STRING "1"
        // Retrieval info: PRIVATE: INCLK1_FREQ_UNIT_COMBO STRING "MHz"
        // Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone III"
        // Retrieval info: PRIVATE: INT_FEEDBACK__MODE_RADIO STRING "1"
        // Retrieval info: PRIVATE: LOCKED_OUTPUT_CHECK STRING "1"
        // Retrieval info: PRIVATE: LONG_SCAN_RADIO STRING "1"
        // Retrieval info: PRIVATE: LVDS_MODE_DATA_RATE STRING "Not Available"
        // Retrieval info: PRIVATE: LVDS_MODE_DATA_RATE_DIRTY NUMERIC "0"
        // Retrieval info: PRIVATE: LVDS_PHASE_SHIFT_UNIT0 STRING "deg"
        // Retrieval info: PRIVATE: LVDS_PHASE_SHIFT_UNIT1 STRING "deg"
        // Retrieval info: PRIVATE: MIG_DEVICE_SPEED_GRADE STRING "Any"
        // Retrieval info: PRIVATE: MIRROR_CLK0 STRING "0"
        // Retrieval info: PRIVATE: MIRROR_CLK1 STRING "0"
        // Retrieval info: PRIVATE: MULT_FACTOR0 NUMERIC "8"
        // Retrieval info: PRIVATE: MULT_FACTOR1 NUMERIC "8"
        // Retrieval info: PRIVATE: NORMAL_MODE_RADIO STRING "1"
        // Retrieval info: PRIVATE: OUTPUT_FREQ0 STRING "100.00000000"
        // Retrieval info: PRIVATE: OUTPUT_FREQ1 STRING "100.00000000"
        // Retrieval info: PRIVATE: OUTPUT_FREQ_MODE0 STRING "0"
        // Retrieval info: PRIVATE: OUTPUT_FREQ_MODE1 STRING "0"
        // Retrieval info: PRIVATE: OUTPUT_FREQ_UNIT0 STRING "MHz"
        // Retrieval info: PRIVATE: OUTPUT_FREQ_UNIT1 STRING "MHz"
        // Retrieval info: PRIVATE: PHASE_RECONFIG_FEATURE_ENABLED STRING "1"
        // Retrieval info: PRIVATE: PHASE_RECONFIG_INPUTS_CHECK STRING "0"
        // Retrieval info: PRIVATE: PHASE_SHIFT0 STRING "0.00000000"
        // Retrieval info: PRIVATE: PHASE_SHIFT1 STRING "-3.00000000"
        // Retrieval info: PRIVATE: PHASE_SHIFT_STEP_ENABLED_CHECK STRING "0"
        // Retrieval info: PRIVATE: PHASE_SHIFT_UNIT0 STRING "deg"
        // Retrieval info: PRIVATE: PHASE_SHIFT_UNIT1 STRING "ns"
        // Retrieval info: PRIVATE: PLL_ADVANCED_PARAM_CHECK STRING "0"
        // Retrieval info: PRIVATE: PLL_ARESET_CHECK STRING "1"
        // Retrieval info: PRIVATE: PLL_AUTOPLL_CHECK NUMERIC "1"
        // Retrieval info: PRIVATE: PLL_ENHPLL_CHECK NUMERIC "0"
        // Retrieval info: PRIVATE: PLL_FASTPLL_CHECK NUMERIC "0"
        // Retrieval info: PRIVATE: PLL_FBMIMIC_CHECK STRING "0"
        // Retrieval info: PRIVATE: PLL_LVDS_PLL_CHECK NUMERIC "0"
        // Retrieval info: PRIVATE: PLL_PFDENA_CHECK STRING "0"
        // Retrieval info: PRIVATE: PLL_TARGET_HARCOPY_CHECK NUMERIC "0"
        // Retrieval info: PRIVATE: PRIMARY_CLK_COMBO STRING "inclk0"
        // Retrieval info: PRIVATE: RECONFIG_FILE STRING "pll_sdram.mif"
        // Retrieval info: PRIVATE: SACN_INPUTS_CHECK STRING "0"
        // Retrieval info: PRIVATE: SCAN_FEATURE_ENABLED STRING "1"
        // Retrieval info: PRIVATE: SELF_RESET_LOCK_LOSS STRING "0"
        // Retrieval info: PRIVATE: SHORT_SCAN_RADIO STRING "0"
        // Retrieval info: PRIVATE: SPREAD_FEATURE_ENABLED STRING "0"
        // Retrieval info: PRIVATE: SPREAD_FREQ STRING "50.000"
        // Retrieval info: PRIVATE: SPREAD_FREQ_UNIT STRING "KHz"
        // Retrieval info: PRIVATE: SPREAD_PERCENT STRING "0.500"
        // Retrieval info: PRIVATE: SPREAD_USE STRING "0"
        // Retrieval info: PRIVATE: SRC_SYNCH_COMP_RADIO STRING "0"
        // Retrieval info: PRIVATE: STICKY_CLK0 STRING "1"
        // Retrieval info: PRIVATE: STICKY_CLK1 STRING "1"
        // Retrieval info: PRIVATE: SWITCHOVER_COUNT_EDIT NUMERIC "1"
        // Retrieval info: PRIVATE: SWITCHOVER_FEATURE_ENABLED STRING "1"
        // Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "1"
        // Retrieval info: PRIVATE: USE_CLK0 STRING "1"
        // Retrieval info: PRIVATE: USE_CLK1 STRING "1"
        // Retrieval info: PRIVATE: USE_CLKENA0 STRING "0"
        // Retrieval info: PRIVATE: USE_CLKENA1 STRING "0"
        // Retrieval info: PRIVATE: USE_MIL_SPEED_GRADE NUMERIC "0"
        // Retrieval info: PRIVATE: ZERO_DELAY_RADIO STRING "0"
        // Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
        // Retrieval info: CONSTANT: BANDWIDTH_TYPE STRING "AUTO"
        // Retrieval info: CONSTANT: CLK0_DIVIDE_BY NUMERIC "3"
        // Retrieval info: CONSTANT: CLK0_DUTY_CYCLE NUMERIC "50"
        // Retrieval info: CONSTANT: CLK0_MULTIPLY_BY NUMERIC "8"
        // Retrieval info: CONSTANT: CLK0_PHASE_SHIFT STRING "0"
        // Retrieval info: CONSTANT: CLK1_DIVIDE_BY NUMERIC "3"
        // Retrieval info: CONSTANT: CLK1_DUTY_CYCLE NUMERIC "50"
        // Retrieval info: CONSTANT: CLK1_MULTIPLY_BY NUMERIC "8"
        // Retrieval info: CONSTANT: CLK1_PHASE_SHIFT STRING "-3000"
        // Retrieval info: CONSTANT: COMPENSATE_CLOCK STRING "CLK0"
        // Retrieval info: CONSTANT: INCLK0_INPUT_FREQUENCY NUMERIC "20000"
        // Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone III"
        // Retrieval info: CONSTANT: LPM_TYPE STRING "altpll"
        // Retrieval info: CONSTANT: OPERATION_MODE STRING "NORMAL"
        // Retrieval info: CONSTANT: PLL_TYPE STRING "AUTO"
        // Retrieval info: CONSTANT: PORT_ACTIVECLOCK STRING "PORT_UNUSED"
        // Retrieval info: CONSTANT: PORT_ARESET STRING "PORT_USED"
        // Retrieval info: CONSTANT: PORT_CLKBAD0 STRING "PORT_UNUSED"
        // Retrieval info: CONSTANT: PORT_CLKBAD1 STRING "PORT_UNUSED"
        // Retrieval info: CONSTANT: PORT_CLKLOSS STRING "PORT_UNUSED"
        // Retrieval info: CONSTANT: PORT_CLKSWITCH STRING "PORT_UNUSED"
        // Retrieval info: CONSTANT: PORT_CONFIGUPDATE STRING "PORT_UNUSED"
        // Retrieval info: CONSTANT: PORT_FBIN STRING "PORT_UNUSED"
        // Retrieval info: CONSTANT: PORT_INCLK0 STRING "PORT_USED"
        // Retrieval info: CONSTANT: PORT_INCLK1 STRING "PORT_UNUSED"
        // Retrieval info: CONSTANT: PORT_LOCKED STRING "PORT_USED"
        // Retrieval info: CONSTANT: PORT_PFDENA STRING "PORT_UNUSED"
        // Retrieval info: CONSTANT: PORT_PHASECOUNTERSELECT STRING "PORT_UNUSED"
        // Retrieval info: CONSTANT: PORT_PHASEDONE STRING "PORT_UNUSED"
        // Retrieval info: CONSTANT: PORT_PHASESTEP STRING "PORT_UNUSED"
        // Retrieval info: CONSTANT: PORT_PHASEUPDOWN STRING "PORT_UNUSED"
        // Retrieval info: CONSTANT: PORT_PLLENA STRING "PORT_UNUSED"
        // Retrieval info: CONSTANT: PORT_SCANACLR STRING "PORT_UNUSED"
        // Retrieval info: CONSTANT: PORT_SCANCLK STRING "PORT_UNUSED"
        // Retrieval info: CONSTANT: PORT_SCANCLKENA STRING "PORT_UNUSED"
        // Retrieval info: CONSTANT: PORT_SCANDATA STRING "PORT_UNUSED"
        // Retrieval info: CONSTANT: PORT_SCANDATAOUT STRING "PORT_UNUSED"
        // Retrieval info: CONSTANT: PORT_SCANDONE STRING "PORT_UNUSED"
        // Retrieval info: CONSTANT: PORT_SCANREAD STRING "PORT_UNUSED"
        // Retrieval info: CONSTANT: PORT_SCANWRITE STRING "PORT_UNUSED"
        // Retrieval info: CONSTANT: PORT_clk0 STRING "PORT_USED"
        // Retrieval info: CONSTANT: PORT_clk1 STRING "PORT_USED"
        // Retrieval info: CONSTANT: PORT_clk2 STRING "PORT_UNUSED"
        // Retrieval info: CONSTANT: PORT_clk3 STRING "PORT_UNUSED"
        // Retrieval info: CONSTANT: PORT_clk4 STRING "PORT_UNUSED"
        // Retrieval info: CONSTANT: PORT_clk5 STRING "PORT_UNUSED"
        // Retrieval info: CONSTANT: PORT_clkena0 STRING "PORT_UNUSED"
        // Retrieval info: CONSTANT: PORT_clkena1 STRING "PORT_UNUSED"
        // Retrieval info: CONSTANT: PORT_clkena2 STRING "PORT_UNUSED"
        // Retrieval info: CONSTANT: PORT_clkena3 STRING "PORT_UNUSED"
        // Retrieval info: CONSTANT: PORT_clkena4 STRING "PORT_UNUSED"
        // Retrieval info: CONSTANT: PORT_clkena5 STRING "PORT_UNUSED"
        // Retrieval info: CONSTANT: PORT_extclk0 STRING "PORT_UNUSED"
        // Retrieval info: CONSTANT: PORT_extclk1 STRING "PORT_UNUSED"
        // Retrieval info: CONSTANT: PORT_extclk2 STRING "PORT_UNUSED"
        // Retrieval info: CONSTANT: PORT_extclk3 STRING "PORT_UNUSED"
        // Retrieval info: CONSTANT: SELF_RESET_ON_LOSS_LOCK STRING "OFF"
        // Retrieval info: CONSTANT: WIDTH_CLOCK NUMERIC "5"
        // Retrieval info: USED_PORT: @clk 0 0 5 0 OUTPUT_CLK_EXT VCC "@clk[4..0]"
        // Retrieval info: USED_PORT: areset 0 0 0 0 INPUT GND "areset"
        // Retrieval info: USED_PORT: c0 0 0 0 0 OUTPUT_CLK_EXT VCC "c0"
        // Retrieval info: USED_PORT: c1 0 0 0 0 OUTPUT_CLK_EXT VCC "c1"
        // Retrieval info: USED_PORT: inclk0 0 0 0 0 INPUT_CLK_EXT GND "inclk0"
        // Retrieval info: USED_PORT: locked 0 0 0 0 OUTPUT GND "locked"
        // Retrieval info: CONNECT: @areset 0 0 0 0 areset 0 0 0 0
        // Retrieval info: CONNECT: @inclk 0 0 1 1 GND 0 0 0 0
        // Retrieval info: CONNECT: @inclk 0 0 1 0 inclk0 0 0 0 0
        // Retrieval info: CONNECT: c0 0 0 0 0 @clk 0 0 1 0
        // Retrieval info: CONNECT: c1 0 0 0 0 @clk 0 0 1 1
        // Retrieval info: CONNECT: locked 0 0 0 0 @locked 0 0 0 0
        // Retrieval info: GEN_FILE: TYPE_NORMAL pll_sdram.v TRUE
        // Retrieval info: GEN_FILE: TYPE_NORMAL pll_sdram.ppf TRUE
        // Retrieval info: GEN_FILE: TYPE_NORMAL pll_sdram.inc FALSE
        // Retrieval info: GEN_FILE: TYPE_NORMAL pll_sdram.cmp FALSE
        // Retrieval info: GEN_FILE: TYPE_NORMAL pll_sdram.bsf FALSE
        // Retrieval info: GEN_FILE: TYPE_NORMAL pll_sdram_inst.v FALSE
        // Retrieval info: GEN_FILE: TYPE_NORMAL pll_sdram_bb.v TRUE
        // Retrieval info: GEN_FILE: TYPE_NORMAL pll_sdram_syn.v TRUE
        // Retrieval info: LIB_FILE: altera_mf
        // Retrieval info: CBX_MODULE_PREFIX: ON
