��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\���V�fnvx��ÍG_;�ȅe�~�>���9�>��Y;�0GN����Sl�N���ϙeh��ji򇢋�>����8=VGK7h����H�k5���|�o��6W�]6����]�<T /�����b�(�7��Ɯ4��>	Љ�����5�Qᶓ��V�}#uo�CF_��Dba�b�/xB��r�H�����t���hlݑ���K�Ͱ�X!]�/��#l1�����h����sQ�J�PL�2$�{���*�������M �������Og�� :���&y��H������{p�PI�E;q �p��Z�(Q��*xƃwbP�ɕ1F+"w�3t��t�FF�Z��jh� ���f�f�N�j�.R&�և7��ضٔ{O��\d�)���ֻ�*�hL�Nfr��pf�p{�������anj>�!�����|��_}R����Z�3�"��,ުE;�b��`�x�O�dƪ�+׌��5�`ٟԋ~B�R����3u`^̻Eϸ��b���d����<�	������xF6������ml���o3�>�ūڑ��X�Ӵ���5�d��]�O�v�ǯ4�'ԆW��>���C�R@#H ��7��,<T~��W��>#�k+m`�;�/m���+�l�d(�g� g��^J%�6�-�X�_�W�%�Q��Ϊ������f|M��fE;c��@����B�s0H���S!g�)b�_-^t|σl�^�Ӕ�	$
y#�uꭽt�ް�YKOT	��47K(�pu4��?k�eS3���u3NQ�5�	2��@G�oI�fF�eO�~��]\��^P|�t��I���:�Ej醬)~Uj]���#,	і1���nnL�V��:s�y�Xkl-(�3�������~������׭40Bw��?/�UX��3�9�fm�Y V�Pښ�`��!��`�]v�u�1L��|*�������{�T��s������kċ�n�c=im�]R���ڄ�<�)�&�(������u�Dm�Wr�=rT��7|$�р�C��o$�0���,�P�F���@'y0��-Cr�6lsk�gMo�.��YO��gx�������<F�g���֯�u����y��]���S�GyZL�ݶfҶ#�^���G�V��6j��ymg�m 4w{g��މ����X�5�X��4���r����;����-�U�H'�T�Iu�p�<`hyX�t��v��c�oZ�n��ݜ��y�*���� ��J]��|'1,��r���iC�$̚��!����؞yǡ#l��f��T��}=�5\F)\�W)���p��&�jO
1��?��N���&RLbP(�?����RvR���7-���]`�Kd <<L�a)���A�}'�tiG��2p����]`����AU�z<� mު��6��S�0���[�Z�U�Y@�F�5�O�V�x�W�,>�T2>V�(�k&!h��n��(����E�<%�I�'���o����d_W״�GX����	(�:�
	������'� [��0�E�4"s.|w{O�\�ˬ���,J���]_۝0H�L�;�T��@��_��]B$(C*�M�+iX޳�Netx�켕��i9�"%��;d_��;g0N(��Y�7.�[���yc�N�e8ʿy;�γ%L���7��94߃w~ C������{K:��Y�����n�9
�</��Rg����j�H6�<,���������4�x҃���o�F矋���2M��%A�>��t��(Z�����7��1���m�%�����L �|ݪT��&�Re,te�a\T���&��x�y��U�����ʐ���05��w��e}B9����1�9��Jv��6�p)�r��_+G2Nch+Qy��ǖ��+*��A8~T��%c2�R����/�!�nO���Ƣ����y���5!���}<�����\Fr(˰��0�Q�e�P�@�F8l�i��H=Pv��ਪ�9|K*"��-��tvT���g:T�L�p-,x����Aa.�0�����)A��u|�d����d6.B+�<Y�����~�"�9��6�?�P�j��T�/��󾂧B RZ34����F�]�I�4�઻ҫ�e��������<o�#���)h������\�����;���� W(D�&#����͛�.
���?�����G�%�ߩ2�A����W�����ܦ�{�cK��S=�xŢ��?ǘ�N$軙ϲ��^9$S�w�	9������\�e�J���^H�}d�C4�F��D�;�󸎃IH��� y�M�����ж�	w*,�[ �t��{E��G��<�~VN�6sa�7��S��;C���ݱm"/�)��]OR�+=߀k��){b�̷L����ڷe�x�FX���V����8*����VA{pBu�:�_�v]�M����sC!���3X�b㱦�r�f\]L�O�Ӯ�U����r��H��cVM�i
��n�U@�3c�g�]��EX{č�Ӵ��L:�3��Gg&���8�_��/�������dT�̀�xo�!�]IN䍯�Z>�]�|U��k��o�ׇfA.���7Ȃ���Nb���TLWF�r/����ɻ	�M�fc{���o�LV$�o�I�3?tc�x;�_R#'���ʻ�Bi?v�F ��{q��u������^�qw�S��`2���9���@�$"S���,�\� ��v���fs����u9�P_%�#���P�����;�L��J/[�v�㟗|&5tS�E���J�*�l~�e|{T�'Q-�1��Նm������'N/",|�d��0����jd��я``�m���7�KН`�ժ`U9t��J]o/�Z�L]��U6:oG+������Nn���&���~���W|CL���әS>�aS�	��g��^	��!�H4O~��(Z��:f�T�o����O.�-��~ M<����@��'���6b�r*��4��[�8	����b\�P�g��J�b�}2j��D�cW�$g��"%��-�5����d/��i�V�`�����c��21�͠Į	P�����I��y5�~TF��ڨVw���w��/��1����g3�.xy��=��CGRď��:Z/��D���C"����-V��2O8�R�Zl��?W�\Kt�}�M�m�!��}Q���G��m�����i���kP�3�{@����XN�w_%�y��̽�b�Ʃh�s����Eօf�3�4Z�&P�&�W�y�aQ̷j4fW��:�{��3��I���0`�f�����Yv���j�)0�"4���A4�`�^�����b@
 �};�W����$A��X��Ƿ���;}L�po�G甡9(>V�
��#F�uc��5�,���S(��������^�[���N��B�ɛ/�2�M��Վ�6�c�Wӂ�����`�!URDU>���z.mm^pl~G���-��N��~QL
 �^Rj�Mӑ[Z�1����~���qt�s���%��8(p٥,x�(���ӬC�v:E���t�A�|�J�µƻ�^�su�N��IPyD��>�Z�B@�"i��(�JNSa���R2�-u��������<���nYW=#��c�
�O5���j<�)3���/������m�-7����]XOj΋s�y�:�����_C~7Xu�/�����cp�v�v�d�\�g�;���e�0+�Y��8�`{��q#"r~R#8zo3�T(��d�/3>^_ZB,�1����XdDɉOHN�M�7z���0Cb}Z�����*��{ ]_s�C�i܁ ���E���j�MxׯE��J�<mg�ԀŁ�L1|m�(�>(	�Y�#�"w�	�Q)9�8����h�z�1�{��餪~%�&`cp��y�"�s��M�T��n����+�B��	J��\؏���T/sڂ��0�Y-���r'���I��]�������ڑ#J���T@tՐ�kAM��[��Q��@�����3�T�s�sr�v���d?�W|���1Ik2�M��rl.���/]8Do(�2��8���\Gt#�j]|�#!{ ~�z�=fIy�;�!�50&O��:���-�u�'ĺpj���"��(F���N��+�&(ݨ��C
� pF��x5��}���j��L�N��3��ߥ�Jw��R�
*��VI�����6�2C�B9I���>\���3w���ȕ�.�J�3�d�Z"p:��~W{Lw2�:]n ,�����A!}Q���|�����Yc������ѩa��M튿��·��ΏM�̘�ũ�;�)������I ��K�;��&v�%ATЯ���Zfy��z����'�C혰I�\��қ��AXq���S�U�z��a�9������CR�F�?�6�G��þ��kM!����&���@�e
=�=��^PÕKꜳ�x ��4��4{ug���o	~jN��D��{���	�n��F���ә�I��\\&yF��i�9�j;�>����Ǜ��$'y��k����r���ԗ�6�~�h�hZ ű�����Ee��	�$Z� �i���D�����UJ((�)��3�O�,H����F}?�4�~YH٬��q؍�"��l'1�VZ,�eP 5pg�pM�%�Y���Q�3r+�!}Ӡ+9�u��o,Ď�I&T�";J9�q�c\^(�m'��'�+d���ǔ@�-��f�;Q��M#�5�
�qS|m�g_��"�G��?��G|QPRPT!}/���ͨ�bmH�F*|���|<h��|��>S�>��r����xޜ	��.�nه�C�����*ϪV����w���w�r%n��2��θ|��D��Zu�4pj���I�e��t �0���S�o�dAߗ\<�P	r7�� )3�������]�j�u���2�«� H����o�vX4t=su\�MjU='�TN�����L�I{)	=y�����ZS2���#Z��;Xyn�� �NH5�Kg:5߿�vԧ�}u��I��f��QD�<�R<M��1�n���ܒ%e�V�����v#�b	Џ������H�n-B�֑[�r��jZ���sk�J�Mmٙ�
���BTƙ���Ȃ5�lҎ�����[���u>��S̆��-��N]0���?����0�i�Z��i�7�s���4A��>���p�!M�X@��`�%�| �l��Vu^fP�.��	�ˊ�7������כ��D�ު��Vթ�3�P #y��������G藣�j"Э�[Gk�'�Pӈ�(k�W��I'�f�{7��X�����/*ߣ78��~5Ğl��éY�8���c��8`��x!�]�R+�ԤVo��k��G�6"�ˑ���+9�R�x�AS�@���X*�E�pL=�/��M�)eB�j�~�0MԠ��0o/I.j�?�GR���+Q�k�O�g'š����Qz���M�*��M�.6x���Y��iyn��Q��}�*%��� ? 'arؗw��^��q{��C2ͫ��3{U�����ŭd��T����l���[�]p��!�`VK�\�>�6��,ĉ�&�iy��Ͻ�F��~��ګ�����%��KhX�4�@�1%͆���s����5�t@5��q�Pt3˛	�K�4����D����T������?J�S43�RP��qvJyl6����dO���@C5�� ��ȣ�i\t��2tZw��~����fd**Jf���s�S�Ꭸ���mr�R���8���k4V|�v+"`2�܎&y,�9���|Y���X`z�Bm��GH����,��˧c�z-��hY���mN�Cª�T���X�N���B��B!������5������un��C��~ФH�3�~D�I_��\2'��B{5�j�Xh�l6}4OUFwxE��+n|�{��>	��&�Pi�����t��⛒K����[��l��FKElw/1�C	%�Φ��0��^��(���s#J�6�ۘ�7�D˕�a�	��v��<�C��q6)庼���hP�ic��~$/���'V���͔ڇ���{ә]�]���b*3���u$�R��skIr��r��[�w��V�@���]m�u�In��;2nW\Y����E���l��,�yV�Z�s*�����+��=���;�1Q�5�eL��"�35)�.��=���8�ݠy7o��G���6���mԷ'u��K:a<�-��"��0�uM�q\MO�jN%��F�*��.��\���H�R�e�+Wz���h����H����X�$d��w}�nk���<�x�lK ��K�_Α�u��Tz�q_R ��.X$�Rk��Lm��Gk�]p$�ݬ��=�Ro��Y����w�74.�_9������K9���BQS�2�F�b^�(�nH3�y��wڴ�N5:>�� �}X�Ts�]])F6����%�I�0Bh=�uǫ0]�5��J��O~��l$��V%.��+�En�ȴ�4�TXC>xW��ɇZg[q��z&`�6$W���'�V�n ���f#�]N�j��n�y3�i�m(ԩx� �P��l��/��N�U�2O9�/Z/%r%<Y�4r�$��O=Iُ��ƻ����o3�� �B=�� to�hH
O�>d-�iW�
��=8�"�|��vQ���ж:YW# '�$۠�>�"Ȧ&�4a܌��eob�Q�^|�.�?�BJm�ӫ�ְ��, �B&�/��j'h�d�q���S�塇�"0S���|1��'Cx��p�͢��͓��Z�o�	�s��4���!�j��,�;��U�]��8��y��Rލ�6�Μ���Y��(rr�� v�}�)v\m'����*g�^��è j�ET��GK�=n�5䞜��鈋o��oq7#xH�o��+J�:&D����6[*��f��l�>R5��?z�6\&B)�"	��)�~�P#C_h�'p���W�[�s��﵇"����а�,�[��bC;��̀O�d���v=�3�(�K�2�����
m�?�u0(��+�!��qy+���t{/�|o>^������5�!���&��SX}C	F+���p�H�$��D��ڹr�la����}I�El�iЅ�%���]������Y�B�#�b(�Ϳ�Tn]���	SW����;�*�K�[��=��&bqj�����/�&��}�&zM*������䐧>�j/��ӫ�zF,�}P�����^$�J�@��A#5]:d3v�"�"i�,�\\�Quv�"�٘xRfa<�VX�ɖ[��{�x�զ�ʢ������Ɵ��EF�3�tΈ��_h�eҧ��!�(�%�������?N�&��G�rD�<����&)�
�vW��Fs�`��So����[\8*N��������x�Q�eW[E����J��0L_���񴪏�/��М�
�,�4���~*p�1�AF�o$��lu%.�_�_/R�dM���ޔ%}C����1���(���y�5���ׯ}"a��/��:(Vعːf�����RP@:G NcXN��t��+@�wڳ�����}�������Rg�5ueU�%��	i؈#V�(9�HlB�[#��kACcDI`�g�4D��/Xm)�Q'�P�%�Ǟi����Ԃ�1Dr�G���ҙ��D�[7��545l�Jհ~[��m�q�/u9ʧ�*��`yٛ4YƋ������̵J��ג�'`	G�U֓,�U��=��_�Oe�8y[����MԔH�״qD�8z�1���9C�0��!`H�Zl�nùg���%�s��6����Jn\:������^�n�픠ŀ`�>����<a��ͤ(�ݩ7([ҡ���4䦐�:[��<���먦+��VM�HzT?��8��jUk�w����ql8x�A��h
���e/\W�k7:�`/�E	��1BNL�-�/K��#o���,4,9�/I8����G��{}���U�� 4]*�VLU���,4��x����?[�����R��9o$R��<\�_��U�W�V��J:��%��}�Q�|�y�+�"���"�;����+;�I�(�u<U�By�b!��Ԥ|I�:ǴXM�EOK�O��{F�T�o�"�20)K��`��;M���`�U>�A������N�x+7�G9���M<�>.�b�uUIa�P�'$[
�t�h��>���@�P� ����X����)?4�3����9ܼ�f����#��Ng�a��p���Q9
f5!�+|<� j>�� OW�"���t����9]���E��灓t$�"i�T���MH�Z���W,4�^&E	�6�"^�	�f;�R��i.y�{*���M�3�O��-^�0+�Z�}�#[<Y���Yކ�=訡9<V΁_��@[n��/�Va�0\�P��jW��>�ͻ����O�TE���{�sʹ	2� uB�v}���E�0/J?��O�$����J����=r��~IӲ���w�;]� 
��I�.�M�u<ļ���%�dl�OJ���ir���"l�r�3d�0�u��:��J�g0�6�JM�4�0*\v�g��1��v[���eM����$.K@?�wF�2Ϳ���?�.�+�4�E�8�����p�w�{|V6�X�lE���2�TNɒ���j(�h	p�0͞gH��r������@��^W��=U�/%��G4�X�	QK�o_�����/p��Uj�gw����h5�<�Rݞ�n�j���{}2�Q��挰ɸI�&N�g�1ߒ����[ܢ�62��S�(Yd4-�vL�z�;�W/io���l*^M����n���~������x�1av�ΰ�-����o����J�J�:/A����("�9��V���D��N�/5)���p��ƒr�E|Xz�&�$L��[.~.��s�'lP�"OK|FϢ��8�-� �W����h1��a5����������N����خ_��0�iH��Yr�ک�,(&�]ɩ��g�#���䇓�W���(
��c�Mcޣ*�<���bnY	�:���#M�����:��:t�yw�K�aYPg��soΣ��Iu|t��%Ģ�r��r%�e�Έ���Tj��L׳x��E�����Pe��l��Y`���zf�����A�Ds�L��q��GT��r�=؜�妽t�����S��8v�S@����F)^Yp>3�&�"��8��	�L[��/&���IL��f`f��`e�#����o�NI�x6�q���HT��uDr��b�nG&����Rg�~X�o���"��%�I��E�&�%���F��=�L�<HJ?F�93��Gt� �`����2�6�b�H�/U?m?�8\�>a'/C`���B��HD����_�OS��BlT�`<�c�sz����=��)�"�)V�?�7�u�:w������U/|R��QS2����^��}���*���ꙥ���O�[b��[[�e�R%�����K�ex��8��2oӦ&a��V�<��0�:8��cӈN���$����=�h*
�� g�L���s�����x��{rYS���Q�0��TM����%�ZK�������R�o�uM?aѳE�t_���9!���-�T��5}� $���EJX��F9��U0w�@�8�E�{�U�j�XI��/ق=!6���B�%�����>̯֝�|`�R��MY�P���WԔb�;��-LM�C�P`	GX�!$���N���x�b��K�k̘����'�#|!��\v��V�	�$�����w���d�6%6�R���4٥�$����C%��ɢ�u�����I�tk��{���IW� `��v����߽�:�ZN�>h�[xT�	���:�#_q9\��RW[��39��K
U!4�N�%�OkJ�\,�w���;B�#�:_.}������u�
8g�i�t F�`��&u.I�rJ��|��?�����!�e�o�v~8��BD� �%�VK���Kz��!�������z ��L�d����2Nb|YD���by
��Xdj�i��B,^����-�9�C	@P;^¡ R~ո�.���kbf��c0�S�G��%#��s�����CH��Ov������H���)��D�@�^�Q�v���%��ȣ��d}ܘ������L��]C�y�ps3W�E�Kj�m�'.�`5k.|����Pw܅���Q����(�`k�˱�Up|���q{�)|I%ܢ/4���	�F-�܍�ߡ��L�Ñ�Vq�_;�k��C��El�Lbe�S8a�P� |ؓ��I�u���8�ݖW4�6�V
��_.jw&�R��0��W<C�h��^�m�֧$�l��z"�.x8ƪJQ Ӓxs<�a?�l�E4i�N��][�q�;Ў
[����K!'׳�j���<�7����Z�F���l�:Ȏ�gef5�w�ԃC4w��Ȱ����9��iGa$t�b�U����o $8�����]Z������]��*j���<�Mf�7�d�il?p�D;�R.���r(�����?�
���&?~Rw�;�� �ۓ���a��`�k��gBi{n��
5%%��Rd�N��2�2�|1@�KS�dʥ��@��jh��RE ������ �O; (��Vq寔]��x�cM+����
$K\����;�j�z�ߐxU�Q��"�\	>ΦGg�����f�:�6Er��!���g$�K2��	n�!�����6�.n
!$sSl��r���,�(9R{1oF�N�M/l߁ս�NgP��7�� Ҙpt����Q?����Q���UeB��xa���s/�m@W�����W�tf_O�a�`wm^�v�T��h@T�^h�T�g���P���ͮZ<1+4����9>��\�|������ :�d̥�o���@�;�W��P��v�#W�8���eS����5���z� �1��w94itTR��C��`c	!_@|��n��6�7i����}zBY�� n��1K0l���hv��\�%�_~a�k*��<7�
���1h�p��0{��lH�D�%�ߣ��9{����KӏS����L�Y1qBW�ӳ�R�>�h���Rś�,[�����-u�����U���X%??N�m�vnl�ܰآ4(�܏����Zޅ���+O��4����C>9	O�K%��]��m酰-�YSP`L����y�������kk��<�Q�����R�6K嶲^zE�m���a����yH_Y�W����ۀ!Zռ?'
�;t=��?�����i�D-X��j���@�JF�֋
��GK��:1K��j�7=K^��~{3� �5إ.����+C��jd�s����	��1��o�۫-|�Eπ3��U�r�Q�X��)&�@#˫MaG��Th�Ok�na����c�q���kj��8kO��I��ڂ���U��l0�S׊$�����^�{��N��X�C{-�G�+�.*݃�X���|�rs�5������|?��Ȅ~�[[9���Neu�σ5['}j�Y�E�p�[ƃP�]a�e�o�	;?����I��q0�0��l~AT�v�7��a��Dsk�>&�D1���E�r3���b���|.�$�%͐�IR$B՞��-��V����E׎uE��RoL��h��p`t���>��i��\��c���-9�FH�JR���dj�v��^�Yt�px��;Uh��s�����8� ���!Y~��˥ք���'7<��6���<��窬�\J�gǿczb�q��	y �ƚ�D�*�?;kq U��=�^�u��2�N��N0>��c)#��[��Er����lFCNAȾN[=�#���������� ֝ɝw�Z{�)4}�(FfX�ہ����
�G=d���������c�ؾ���Nn��h|�^<��DV��D���i[[_�{4Xmۨa�Mp��*{w�yٹ�8/+��fY��
.o���І�ycF�v��N@5V�b��5�����+}vn�ԨjѦ��*�DCⵍ�������In�L��rs_�� bc�3?�T�ďD�h�i���-WW�[}�1K�aL%�2���3�)c���<Q�F)1UI1̽�y��{��b����`Y`?���S'�d@�o��@�>�v��G/�PDQ���/Ӡ�k#	OB\��d:��,��"�,y7��?c��t���iѱ��&���ky+�y�p�'NA��n�u�m�/�I������vM�]��Ә��@�^�����c-���İ
1t�(�CA�ot���e�	X�ՋIpN*e�J���(��_�G�/�W��!�7����E�X��V���v�s���lP� ���|��D��%��	Q:��H	���#��M���� �@���U���/)��d��Uz1AVԮoN�XW���{B�O�w��b�@��C�׹�n V.�q2F/��j�L�1Vt6�͖�o]��P��y�09	�U�Cn�S�8�;�|��Zr�2Of(�
֌w;�O �`8H�}��h̑��8�/s�[�3'��pq�-�\��n� m���ӈ�T�����6$�1oT�Z�H��a����U T#����"�_�s��[��*�%W������
k��쪖|rY�_)M��u����[{��ݩ�B�vk�l<^�r�3 ��R$�ΰR�b`�È��w����	�ҧ��反���?a�#�u���4MsUD�4a����~-R`��r-c5���w�{ֵ��"E�[۪�~h�
{\uhRXvd�Z���Q1۞�8��qMZHS^M�����N�2���A���\�#�*����Ng�@��*LV�ʏ�U>BMޠ�iQ�ڋ�R�2�5�� <Y�B����ު+��u���4�"����Ťd�-qn4[��[S�3 J�̕�(mA�!?�\�6!�깂�9�9�A[O]Š��C5�9�ܱ�^L�hƉ�81e�sBOL��d%�5N�������«�e��2��T���@�8R,��M�鹃�P�e�o1�`y�?&E�EG����y6��)�FR筱q����д1齗�K(�D��]q�����t��tgg*"�o�
z
���[\]s�`��M��F(���iʝ}P��%.D��@���Ԯ�C9�(��48cՔX�-�Gz�eʕS-�����8�0�6�%�Aދ�����RA�?�QƖ^?z����u���J�;ɶV�8H���(\W�eu]�=������˽;I_�Cm���e;&XͿ*�����u�d%�ʆHސ�y�X�qB�bF@��j�����x�3�3=�XR!���Q"�1Α�L��h%el�Y%u�X��$F w����ST/6!�"��!��y���.,���g�&L_�6$����}�/�c��g����BTY�_�<� ?+W�d_E\`y�V�V0.;���gZ��
z�@*%uM����a[�;�\�����J<l ��J��>J���{��K''��BA�<݋������EV��؋�ަ��d��q6���8����0_Ȃ����T~�n;L��8?�2g;5��_����pM�����g��?�_�D|/��؂�f;-��������JV%��@~A����A{�lam؍���L�<�����kwt}[OK����PX��U�;����u�؎�ݾ�iJ�zx��[�tףL��p+�S
�͌�������%�1���Ռ�N)�)�$Ϲ��p��\ P֊g��;���]}6�,+�V����\�5L�'z��s?s��?<7{����JW4S
�j�}d���a���#^��Pt��MQ���x�E�-��6���p��ʐk�p�S��1�vw��	��[m�B8S��xq�`�eߓ���kh�M`�e
2��a���&�
"��b����T�^[�`�G,��J�zj�;"�'#��1c[f��cǧ����Ae�A��r��5��$���+R��N�(y�����o�=�r��mX"�t�D�P�hS���w۸����Z�o	ۇj�͖R6�Ps��˻�Es�d��y�c�w0�E�3�a<	��Z$�|�P �02ÚS&|��.�ל�9�;�����{�k�տ��� ��1~GJ|�=���3J;��������.-Ua�e�М��S/B_)����e�L�N+�Y�%;<�ɍ��c)wzFt{A=3vm��$��ʔ$8�i&��*
H�ݢ�S�
�`�	��Z�������,m�5DGJKB�[�O:��;��R�CNv.���X5!u�H��A��,=�ma�.�uN�>�0Gqe�A�A�b�S���:\�W^���|���͕���>Ӏ"��/~xK��Dy)��w����RPL0Zy��'z�w>>�7H�T=��:�êè%��jhep���^7̿��U\@Kn8�+�;��V�߿��(���V���Uo9��qr��5�)��9����aq ?�`�DԛKU�;��Jɐ��tn��v�����]
�Y�zQ���R{:�?��=[�X�Z�X��1�IYo]�)�1s�!�	+R��-k���m'm�Xx�A@��e�@O�Pn_��h'�Z�\7�D25�B�4/���8����o�)$�|"����&��8$�/E*��G��j2鏢�@��.���q{�ꈻH��ׂWL��Z���J'�yu�I�	����#�N7�@�k�����o��:����%I�(�������چ����Q<�;���aÔ�Z��Sς.9��7�~ِ[�<3{:_����mV���)��4입t7"�s͓���*��ȏ6�)�mdL��R�X%�W�L:9��F� Z��ao�*eRN���ǋ�˕��9�k��A�
� |n��x�n[Ѧ��~0��73Mjhn����U7[a���[�cԊ���n��M���f5]\5@@:bʩ��&���u�����XurZ d��A#n�\��i��C�pud<�*P�+��U?�(G=~���'<Fc`��/�Uq
�/l�;��+�������y�P�~������fĻ��_�^�+:I"�*�£�P��z����;����tm�/��������_[���&ް��[��[p��̯W�-�Ӄ�-�0z��`�KlT^�1��`l-�ޡ嬁RO�1���o�����e���PW]Wl�@��(����͆;��{���M�4�.�L��0���E�ɔ����D�a��!�¢Q�Y���ꏬ
S�N_F�m��	֣ᣈ�f�7�zf=�Ŵ�����'@�~x�QT��e�Nム�"$�1,�Ifs�!�"�F�u�*w���E�f��T��@߮�r�;_�TתQp#q4�w g���'�1֋����ar�QK�a}��1�D4��&/��!v6=����m����ڞk�4�{���NJD_N�#M����+I�\�:?bO$���K�S5bk�%�X��&��)�!N:gV
��<�@�~���~Hn��"%�J�"uK�׃1�����u�Ԭn$1�B���ǽ7�;�����x��/,z��|H<wA'��f�6��]�Z� ?4^!u���e�8	���`�����Q�ڴPL�O���^=7�G��k�kLsY��i��l��B������ߢdQ�&#�ś���	%=za�g���ۉ��b
@�%����K�FxR@qR�wc����`��寽��IA}ЫO��������6��O�F�o�k!��xY֕�;"��Y��6���M`^���0kXL�Ċ�¯��b��Dn�2Z�F�|e��?���ޖ���h�i�g���4��f�SNJ���ձo5%õv��ⶵ�mM�	v����&IGi����Xe��(��kmX�`��+�MW����j%"aL������ca��#���2����i ~�����e��ex����?��9��d/	_B5���^	�=;�(��ږ{�����y��.�B�js������*sX�����&XӮْ�*�ohv`BH=�<��������N�;K�J;K|b�1���6˚켣�������z��+��d��q[�#'�~�v۠g�8x��,1%��I_��BMi�!�ȇ�[�$�Zu~E��`���X�,|>��0���Jd�����D�m�sN�B���8�е������j�@Z���S؈�j����c���uq���5���H�?���_B��.����6���ӽ��4i�jf�NZ2��.	L�}H/�,8�<�QͤM wɎp��v�s&��R�#RS��)�&��}ny�=]�p��!M�0�� p�'\qL&�W�uh	N��gJ�}F��1�t��O�ۺ����*3���"�f �c����ңh�����?~{�2�H�ɫ/|Ⱦ����zA /G8�k�O<�k��7-8�*\I�Z�vF��TW_�1*סBj�1�e�r�u�y��������h��wl��wȀ��v��}Lw����ʍ�@�\o!��d�sG3H���������wڷ�z���v}
�����4�K�8&z��4�WZ������N�Rh68_(a�%b��&�T򞓻����'�b鞭����_��Q%yw����M��ݮ�y^А�Q��y��`����KTC +�d����c�B�F㻭� ��s�PX1L��_����u(��ՙH���^�Z���j'�m�w���-��ژH-p���'�pk���:I7?[h�� 8'�q���b�7���O��W�N֎�Ѹ� ܚ���I�p�_��Q%��L���f9]+35��ñZw�6vY݋��M���~�F�h�Q��*0ޏs��sQ�j��j�qG�����ݛt,<��4�j��B�G�];+~��
���WNX�	j�M�����O��%�@���#R�Ě��V��-l��i,�g����1�o@�s�(`Hy���v��2q;] x"��_崙*l�����U��{Jܓ��]@�n	�L�Sb�x3�>����h!��b�gy;/q^/9��d�'�
�Dh���=Š1 m�t%)���a�K&��˲�~��F�}M	+�D�#n�����
3�I�"��� SCY����/v;�[9Ch-���r�i�F��u�U��Ŗ�������b�C܄�^�% ��وf4�ӎ������jày`��8N�8�lLӚ��y�J8�"�Kt��M���bWΓ?DS	�t�	0XC�ܱ���X?�7�"eϲ�)U�v���
�~���C2�U�S��a0ܥ7�X�Mc��e��tpmD.jӉ�x�iB(cM'
PDM�¦7��я�������,PA�:���j�(�ԏ(��	�J0����k � ��V�X��N<_����e2�]��Q�>ɖ�q��l%��Ņ�-�
�����p̛��g�5{�%>�ܹW�x���ﱄ�PLZN8*���
f��1QȀ��rZM�xD���= �6K�*: �Ur�B�Ff�5��kJ���[�i��4�k5���(�e���0���U<^�5� Yߓ�]V�+���nȞș�U���+�`�*���ګ��	�1yL껕�m�Sl,�M��X>��O��.���<)6����Tب6�R�K%�;2��NX�}�K)��u�����r�fJ����d&g�gy�)���o���Xa8U�1�2�}�����VH�j��!��B/���D}ve@G�7w����)S�g<��o}Lu����+h�E�ΕŸ۳DX���`Ρpm=A��f^���lO���������7`{ժТ���8�s�^�"S��P�]r0�P���5:���<������}�h��y���~?g;�!:�du�^�hC�J-%�fY�*̆�ק����AuB'���&�B���Q ,� �eY��Z�.�^gVto��[͜�i���m����7������fJZ[:J��/#�F��-��>wOz�C[���u����#`J<΄﷼�Gుu��:q���9���� �D��+$��Y��4���`��r�m
�c�w<�S�����|�kA{��b���<�i��_�/8-1q��*�'�e3�U,��X&��Sg��I�0fZ���/��/��k)�7�,"D��q�	E)�#a�Ƈ�׌�3��p�O�m�5�x��3��e��N���"����jܞL
�^�1���A�:z�UN���kHc@ܞ ��+�N/��\��B0�N5�B��X�'m�io�L�ҏ����i1�̭��m�t��vQ*�l�R�L�d��G8i�?�-�ڋ��E�;�����]r��U��pv���q���W!�p��o�z��^��K^&%�����>u�%K�8���� ��8�{��k�Źmkw��8xj�'���8�՘�b1�y��x�꭛}�U���$8Mm0������C���	Dɏ(�ҡ���!7.���E(�������HG:Ad�#5�گ́ϕ��4�$�!��"b��܌N���'X��� �`�KEA�]|p �D3:�/���(�fbbGw=�.̚��[�+Is��G�/��,�)�g�I��9z�^����փZ`�u���($(��f3$���s���r��Zg���A���N�	x�_ܚ�Se�:):���(ؚOc��n�Og �ϡ�2k�1��g�����vT��ey؉�t������,kw- ����4���R�#�! �̄�Ų�ї݅�΢�_��+�*���il.x��ŗ�]A:���+��a�Z��L��.5x��~�3�[�*�&=��'�eI�.��@L%1v��>���X��eo��<��fC��K7�o�e��|+l�	]��ק��sG�[���ה�nH逮��@cp)��u��TN��kn�s� ��Ѕ���ne}��V.=��Mi;�q��lJ��> ���hWjb�d}i*��^Q5��s
��t���l����0l�uJwIp�H]�y�<UO�G�7��)X2�E��2����8@����m��G��Ȅ�Ug�;��AH0R�R~V���a;�6ma`nk��o�g���|�o⥒��e�'#�}Т8Y[�&�)���O`F��(�W��$����(RFOS�{џՊ��l�B{p�����a4�x��'T�XRx�u5���։B3��BBȷ�wm�2�ȏ�U��2 $q�s?� ��9�r�y��2��9Dl�K��n��0�g��i��G����$8�ɮH0�>���'qǟ8�Cb�܋5�;C�5�䬚�s1��R]�vO�h|+C2�GPI���c�>O������2�u��J.s�^�*��
oah�;V�W�!��VIxp�{G�_�*���b�����Y}wI�8 kD
�lx��t��Z��O	�v�z'�����^��DWZ�`����o������BDf��#��Jj&���®�W��<(Cn�]2�E���Nz�o��I#�a$a�S�U5��-����oMJ~�p�g��Å���v���I
��NzC���]aϛ��=sm��,�u�Y�M����G/d��U�q��Pط�b�R���nܤ���i�EP�� h~���>�ZCp�@�������Lh>j-ع7K��_=iTT3��%��7'�4�eV*wwN����u�e�v����\�b�o�	�p��cz��r�*�{�VD(��gw36��.���	8ek"�ļ�ML�j7I���H��c)&��z�����Mޥ��/�ۘ:m�[���8ذ�5���k�\��lr��xH1��:��D�F+\�Sβ�{�{���u#������` �p\żEr����� "*�i<ר��#��pђ۠R"�T3r�꘠�mؓ�I��o�$�����<���'ւ���GC)��!7�r���A�?TK��1�6g��S8��	�?IH������NЁ�;6"�
b)���N�H�?ՠ��i���a����<��8�jc�����������_N*6��a;��4�1���7��Xq"��W���#�+��e*."J�n�*\�[?B)1�:{����R	���Z�q������(��weV�&l�����f��b�!�Gܺ5�D��%FÚ��n���4��S�`XC�JEr�~� >�֜f�"�!�B��D�d�:�"�`��Q��6�b��N��-ќs���Y%c7P��aq^C��@�nsP�P����ފ���o��o�%o�iB�	_�+)C�*ɹzq���jz¸II0���z�?���h��(�V�r4����wբ(�Z�}l>+�ĕ���|l7������0�\ܙܠI^�a'��ݱX=@0w�0�!g�a۵6~����їmG����<�ncJ��S��ͭ���僲��z���7:;Џ�a��L�@9|���#�=!���������ܓT?���6�V����t�H=�E��1F=�^��PV1�������P�����R�f�e9N�v��ы<f�G��b
,�ڎǏ�m/�!H @r��?Y�� ����ɔ�MЉU�-9�� 
�~5;Q��"_a/s���o�܇�J-W:j|$�0~�.�{<�W�*�� �)K.�v`��&� o7��+��/������27��u�޸F��=h(ق����o����x]4��٭����^�E���'�o���l[	�"#�q8A>u����5����1"Ϗ3����@)��ѳ�b%v�鎱T�8�9�?z�KV�h�<\������y��P,84c�k�wb%�������U�ZF��"��hn���W��'��p�.J/H![#�Ɂ��t�k��Í#��O�β.�R���	��0�S���0@
A>�[��.!�(��تϪ��pZ���U�gOT; ��E�C5ֈ,��67�D}�S=�nh������v�;[�:})݉�fiͼ�OU�Y%��+\5:lh�OYf�sCZ������Ʃ��Væ!M	��gYZ�8]Ŝ�o)/����UgYn���U�3\��)Kj�
(uQ�z	7�DY�F˘���8�.;0T0bi���qizd������}/d�)	}/�:k�z+�`D\����@2�I��Q5�]�y,)��[�<#���ʍDC`��c��6���c�j���ϧR��A)�{��f�4
`qb�jŭ*`�*��_Ho�2����c�'��ۭ��{T�����wp!�gw(�C��P� ��66�� *b�WnY�Mu~X�]¿���]����x�e�{ܨ�f�4��j���V�#�cԼ�TT�.��ޤ�ދ�07�A e��V��9�> 1�a�_�u�m<Fc7�����%y��BF"�n�����W�1�3VY�M�(Z3���/
:aN���;��yb�6�㙨�m�)������=�N���Y��-ж��\(��O��
\|� �/�N�����:h����X�Yg���H=$�����p�/Rz�c5�}��1�� �������~0��/�Sj�.�����\�Ҟ�C7n~��=�z�'g��g�e�D�"��(��>p�?�]Z�pCW�$�y@�	��a��!��������ɷi�s���)cNY�Z�hH�e`�T�$1x�����"ղ��H�#��P>1�談�Hx�� �O��	x�H#�E��K�c"������Y�̋��:5�K����q�Q����h�c����=�AC�=�B�þ�KX�˃'t�ayf�g4�� �e�մ���/��ﷲ��,>g����QMK[Y�-�����
 �����pqޞ�x��9F,�C�DZ�ϴ���5��1�Aq�`��G8L/��x��|a�~o>Թ�V�u�����`�ccP__=]�m?Qۛ�&��b��ф$;F�d�=A����A����T��*��',���YC�5h%�2\���3��n�(����F"g�~���SN�?[1[bO1�w���n_O�]�09�Hs9m��F�jg��UR�� qs�;n5PoG}��jq��T7��8l���R6dy������r�;za��c����y�B�?�>���]ư����r:���/+Kh(�V��v��\���3�j��;�|�˘��*lQf������:9?z�� ��	��63P�]h&(�&���V��鍔�ڡH攙�n����U:���3C���t�@c�d1j7�����~���`��s+~�6x3�NN�5ýM�Z�����C��I���B��O����U8�c���
5o�~R�B��1���'v���U*&O�²�{��2�z����l�5Y�Z����-#��J�M���3�q�*t{04y�A� Ōf���.z.y�)�)���dE,o�7�)*۽YM<++�EP�i'y��$^0#s;���c�����^Ҟ��W�x��abJ��k�%����lc��`�Z��ğ�t�
�P��J^���t�W��CK��A�K��8W%��Am�7˰8��~��=��Z�2͗�Un��b�`���(Qe�l!�UP��	�CU���U��(~}`��ݯ+��f���  �*R�e�������xq�#���A��M�6r�.p�����k�>>�����Ur,#z�� k���[E��p��_��/��9�҇�����\.�$�X���A�۷J��}�i�:�k�Oh��c����i���Wŵ��R@O��9N��$��I�D.�t" �Q_MKN�ٝ��Ĝ���H^)l�Bxz|	\�ґ�;!��{���.`���<
��+r��ɽt��r5��a��a�2߷�F�[�yJ�(�D����%Bȭ�6�R)SG~��� �v�n��T�%��'PY���eB	\N���=�Qs�|�RI@0K�����^���:n�v��C+��?�v��i�`�MN-`^̾1�ճ�?����hF;�+Tg�Ӄ���(���ӧs����r��i��B�H\�QY.���V� i���N�S]y�P�=:W:ࡔǖm"H��!J5�r��Tx�qخ�M�qIx�Ȩc��.����0�~~�KmW!�j��~	@�l��aV]RC;��2��7h]�Oiw�u�����v���1����C I�d/cWt��e���ݫꂋl}4yPs|V�x��@u�h���f���ֻ3/|�����3��c*��� \8�R��{OIU�<�:Ҁc,�~�i�G��&E�2�T�!��e�5��AM��'`p�c��G�!��C`m�@�2��k�d���Z��`�(�_=���|je���R°N�]�S��H���`��;�Q_kQ�-�}���v�����7މ6c�����r��`7��sW��V��f������^���ՠ<<#�]�Qq?���}��W+R��v8A�kb��O�x��:E�F��2��y3M+�����KM�{�ĳrF!��`��]�O(�(Z��0
�	#!I�o��E<q��.��I[�?8�7b(�GM�~$�uv��?���d�Ɔf��<r��p��d�Ŧ,x|�p�$�Y8(+xW��HPڅ�e��%c͆ސ�9U�U��I���dӐq�	�g�� �(�S�Z�e����L��ɐ�P�I��|�3���~�I�r�J��&�ZC��n<��0���F�ܔ|e�ј��ꓝg�BN���gL���D4�1G���c�Uř����	ko���ZJ����)� �/Ce�n[�k�w��ȧ�a���P��A/yWE2�r�'�y��������RU��L�ȧ���6��G�O��e����x�)r�`�ru�I��U�E����B���S�aX��11D�oY���Y@n/����V���9廥9�'� �噯�v	����i�ԁ��6�:0)������Y�o�~J�m��RW�܀�����u���s� '�%�jGI��:�":G��tj�?�Q�\�u��{���hVͣ�+uݿ���� �%��i�M}kt�&Y� v~b�g�[
�R���b<`ԚC�kũoH��&����I^)���c+�6�E2}x|p�-��׽�XH����d�N�����v}5}s}f�~�wܒ�zBk՜E���QV�Ĵ�./��OWQ�T(5����BP�P��Ac���V�1mPo�U�n0����t��O��S
��y2����	X�K��_1�4�!��Q���k	G����}�-\�÷м��1cU'lN�6���<3Z�m������MM��^�g%lF���7�'�<!d��r�b�~&�K�)?�X���)O�[%`������?3S�Uh_9q4r�g��p������2��|�/P߼Q'ie��d����&O�9��`P�	o����]�����hY�,��W���9%��1'e�`s�;�q ) S�@�]g�Z��ݫȀ����J��8�����BS�ǰ���~�&���lD��=�1��Y:�>���-ݾB����;����
'Y(�*�z����+�_44��ii��_ڃw�\������������B�Ϳ����]�H@�"8� `�'�=��+g�ޫc6�Z�,xC�r��ؼ��G����'���@�r��t�Q�������eEvx?�w8fubmow/��N��S������H�8�>�O�}ʨ���C� �W��U�eǣ�F�c}h�:ifW�n������ �@q��|�||����p�`pO/�yy,)}
����y?�^�CAn7��4=�?����������$D���&Ӵ
U�a�M�Sb��x��1�4�����8�������3�(w��Ua��)8���Zjs���3
�F�'�Rj}j���fFbڨ�j9�"�
W�䧆���$wX�,r?���� xV��4s����8S�S���|�-G�s�M�ֱyLw�JC�
���H��q�<�@�\P�u�mfKwׁ�b�O� /�ƒ�|! �T1�GӕH���J�}����$��~(h�JY��:���
0=Ǣ�����I2÷��E �h�.� �Ə���X;��R|	7�a�+����,�P���Nt��x��IG�Hi�P�	��5tP���j���\�[v�t�7h��D�8��cE�Y�:��A�:P�l��;�$�K�d�1��-�(gd�482G�
ː��2R�B��p����M6����S�/N�B�-a�J�'�(͆��TI�y� �\��?k܃&H���6*|7E.6��O�8���$�V%��YS(P a�?G^�y�l��A1s�DG''T}��k��)J@�$Ǡ�}k�/!���Am�?��u�Ϥ��݀G���Ҏ���p532J�wh��Vt-'�����D$˄M�3,�Q�Ř��i_�_�ͩ`��o�mD�I�c��]N�N�h~�W�^>^��  ��<<.��������0Z�� �3}ޥxQ-�.ݫ��1��u�%'�gf��v�/+�H��E��:�5�I�K�Az��0ɞ�D�k	F��_�+"��Q��:�_$�d��kA����,4�;qLjsz����+6�l�F?Һ)�-��!�uM|�0x����Y��'Kp�J��#�q^��:s;Gz7v���u�����z�|sN �~�R_H��c�
���
%������>2��Ĩ������O�`��A(4"{�b�N�<+�u���VE�ߓ$�����Z����|�Z��\9]E�����b�ŧ�1�tMZ�\̕}��E����k�4�?{����M���i;���i�a�x�XD���\�!��!*�X�]�񣘥���j%B>���fݜr�̥���iQ2�h��ձJ���<F22�=��Q�ǛGV�\C�����'���m�x�j��/�C*�ӑ��w:�(?���� �jz��G�4`�؃k��$K<�m�X4x,q���+�SJ���-�'�O5�(��(	A�I��o��M�w(���b�>?���C^��2�I"X�AW��bSC�X�D������n���	��ez���	�TdY3�xa��pE���dp��q�6]�兿F Mq�e}C�9�$��	�o77��ؒ�����S�~���.kNS )�l�˄0����g#Ǳ�c[��Wi˹ɶ�y:�HE`kE�#��%r>o��R�D�����Z�6�,_���޶�	�i
��{Hm��?e<��ꡣ��9�!���~�����~[uP|��Yhí ͫqE!Tӽ��Je ���2E�LH(�[�DK2?2�9C����u��R1�b,ZaR6��p>�x�\�R��IU�'Y��o�#(�񍽣��"����iG�d��l��W�6S2�!4��� ���?�wNv��Ѻ�U��uSZ����P;�G��d��uH y����ٗ0�m����kx�������GTڞ}��rRw���{��Z��h��,hf�w���Z�g�G�qU�֗�)'�?IV� �zy����/h!M!�p���$�]���x5J��H7 �*�w/q,���q3t�o^^���'����8��GFq�y˔~R��9�J��Lj���d��ĖD$^a���*�I���X@L-��?k�gpFo�ah6�f�T�� �5'7���W���j��Tn� ���bUX2�N��@V����\3���A+�BN;<�wb_��?�	�U�3a~5�X"���W�q)�׺B�����C�����=	w:E�n;���W���n��}Qa��
��I{����4��9?�2�|$6�a����x���7hx�,S�&���z��#�dO�ſ�32�����=�\8/��â_��A����>� ETN�>*�Pב��Vh$��/(9�o5!#�4�9C˱��@�<2B�J�4�Pc���֒�(��N 6�������]�+�i���K�8�3�$8�D�$R�U��s�?�D||X�|OD��R���E@�A�tW�q�������S�ͅ���A=&kp\����/E�Y�1ȹ~��j�VO�xz��6�'Ep��2%3�P�+��4���?8=wK�����j5&����߭��Ξ�u�=R$i��!j-��id�{�ɭ�����Cw�w��@�@yz��V_(�6� ��������1=Dv���>#)(�4PӜ�(FʓJ�34'7�9�h'���x�m�.L���{VzV�'%Q�%,6��F'�yA�(j�+�&���b�fli֤���m$��ypD&�����jc� �1�2��@-�e0�,�'��좒e�J1�L��l�.=��wV���%���=�S �j����K�K��y�T]S���9;��|K��� � ��G����D���n̒���1J�o�Ķ�\O>��H�z�oܕG<`v�z!x�h0<_�C�H	��ᘞ���sv�8�ϋd�㍢���n�Yj������%�k�9�^e����:��F9|�L����N��NN�h,=���	���~�Irq�v�6~�nWYKh�jZD6!yϲj���<.�-!�qbl��0*�<�
��.���-��=P�T0��Q�ب���D2�4M�2m��2����F�ݡ��[�F��W6c�g�λXljY�u�|�z�6��Y�UW�㑫��u�B�@?��ֿy H@�CZ��{U޻���e>��ؒ���Y�ۨY::ّ�:5�ѱ�~�m�D�ܯ�/����w�ǋB���X���z�{s[-�՟����禒vr$q~���30����'�pj�>i0�
��j-�uS�X�N����*�iG�wtx��d��J�������#1G��B���G�����.촇��qE�$N;�L*�RQ��D�b��K�6h*<S�?�-�OH��tm��!)8,M2�M�}3����5�����PX�>ݩrq�`ԅ����F�$��?���x�b��8N�s�ҧۗ�l]����j8��GO�H�j<��0n��g�8�LY(p� �����s-7��o]�!MM�S:���f.89�e���n2,0ma�+�bkg
s4�22�Rǈ�Ӝ�߶%���5r t�N "_&��Q/�����҉Lr����;�9K��v~ d�x"xKj6.쓸�u9,])���p�������g������t,���Og��L�5{'�7$�1FM[v\�8�~�n��y�Y4,���J��ce׫��F����@�2� �X���xlQ�'k)g텖����c�(u��	�vd�T�H L�W~٩'�74,C��>;���2>X���@F�8R�`;`�Mr�a4P����+��h*�mҠP[�M��"�6I��|�z;��q�Rw@�Ұ�8/&�o�Զ,�p6�;���\�X)����f�|�sH]A���x#��	nD��o6ZU�eupW/���ij��|�n��;���{TrP0��ӭI]_�am������-7]���9�ޖ!��bc�6>�~��t2x�(`��`Iطm���qP������}�՚.d�`�?��m�N]��9��Y�a��� 8he�M�50��b��Bn���I���tv��CFP�712§�b��4�/��b�h�a�7�5��ǩ�*s����D[�p�yz4�X�͟{��
�v�(?�щ�ͳ�y|U�)Ɖ�^ڭx��0�C���ϰ�5�'�ᔅT�u`�V1@8Xjwc����O���!*����ԩ��"4��"j3����|��K�)6�LQ݁�-F�P�QH'� ��B5�������*�����gǅ��-t��8W=�ЛU
�c����x[E��~��4�f
���=�����%��Dn��pt��������������l��V�+����a�Y��H�����]�+��x�CiA)c���rUc��}׊�jIu�&���"�ơ�\������ͶC�X ����7��+G�u:d��5T�� �[J�F#��'�`XGi�7�T��=:���2bb���#D�p&���e�;��!d��2[=��i���G�(���`�1N-�D)����&�l�"vNֹ��P�E�����������mo3خDq��Rg���=W*l�#���؇��Q󶈷q�����ND�(����+����]N<���h|)��:�P3��B�;<�����g ,��]�	�f.5�/hXr�\��V +9)�����ѬG��J��{(��>�w�,mD��ئoP���,A�������=Q	ďUt���:= P�nV�Dm#�w�����C6��p�H� v	�7�-�y��_-�[ׄ�?W��P̩ʧ${P��PzfFY_����P���ww46u����v�7X)7 �#�܊�v���ʚ,J`m鑷�"�T����I��SpLz!�`Ũ�t{6[)��^r9�������A�|^6�~�A!�T�ԇ�K���-�p/�-V)�'���"�D��W�4M3�9RF�\M���
�0��|fM*[C���oU��S�n����2Q��jS�kTNq�h���,�L���+n��� ȕ c�<���G��=�j�Wt�yH��Kl��"U=Y�J̡�߻�x<ձGrpW¸������k㮟D9�ݣ�]{P�� ��wPx�QM+%6�_�r�677-=4�$6��L�<t�eB��K�5�.�_���<��}͉������Ed/���Rw��Q�}n�t)�p�eK>-�$��ɛ߯�I3�[���с����t�ҫ"_r=�L(?Z�}��~NQ����1�cw����Q�ma�>�N��5'Z��q��@�"��T�����[f�}��|�+��C�kg%�r��������E;�Mߧ�.�x�(��2��"�=E��܆H,g�i��Jo.ɔ%�f���F�;��%��� �3�*>���&\isC�� ������(�'�{��qVE�d��m���X���i��YV�Œ�K�M�8Ff�"G�A��X'��`,cŸڠzpnT
+�0:�'w>]���or�9�t�,4D�-%H\1tC*j�X�X�B�발�``Xf ��@�����4*i=tnA���������?N�ƀ�� ��/��z� ^��[~Y(0,����?־�~׋��	4&�U�Xpyp�!i�����m�w�~��U�T佅4�_�k´3j����*�k�.z'�d����S� H
L}���r{gn�����T=��a�5��^�)Ɵ���#��!M�Z�uH��s� ��I?[!7L��O#�ef�LRD 7����$���(V �+@���8!@�4�X�_��]IT�l[��k�޶����xlf�s�_Um�"��*
z:�;�����oI�rcܳrk4;�D{���a#��Z�D����Y����'4�U�	��]j��o�e�4�Y�DBڸ����"F�U���P��I7�2�j�l�#J��w�m�S�`�oh�T=!��q"����
M���@9�E(�)�e�� ���w�ZU�0�-`�pJ��Gv�="5�G��W�G��NS�"������|OEG���+dZ[8�N�3�ً|�dB�5"�h���~�2���տ͈�պ�L�n`\��K4VK�tz�%�#�F�U��l7[T��@]�N�����5i���=�؟�q{wz*Ɇ8�!�8y^�>����kk�b=�w���eDՔI�?Ex���EIg�,�Q��;�Z���r��O�$]�3��_Z�г<;鞺^$5Agh���b ��ᙈ�"��?v�b{t*R�ŷw,/�i���x�����Z{�4��Qe�QhF^I���@⪀U��͖�"���`���������L��kc[�f����h�G����CI7nr޷//In��SB�ic �H9�gF�����
��5+�@)Z?���h�.��dG�Y�^)���[��u�vo2{��&T�|�.BhD0����(��"�U�O�w�PGQ;�kg��#c ����S�k]�xPf��c2�3\��3�q���6&wwG`�V��B��%[|�m��jŨV\�`�1���d��e�j�WW��d�]���_:�y&@5����Z���䪄��}�u`����l7�/s�֩^y�zID����C"��x^� ��5���z�q��,�SLg8 ������Q���e��u�RK�J)~�@�3y�ܕ&����:���d�#�,qY��ø ���s��\�ᇅh�m߂�^�+ؘ�ei�JUj��	����̔��B��j;i�a��ip������fQ���R.S��>������Y��&��"������[��Kx�9ڋ=�����e�^A��K�/
OX�Ė�S�rR�%��Z��&c�S���u<v�O�%k5�I絳���ע�"����=R.���d%�&����Q�g�S�ͼlq�X	����N��3�s�L*�O�,Y��.ː�i���;�����)��`���W@o'7Մ�j��!�{�^v���@�	�>��e��{�:��� ����u���C���Z}Qrglr�e5 2�ˁ�#l���H)j�ǆ5�`�-��>�Dh�n\C�於}��񋟤@�h������NOh�mH̟&�.���Cf��5Ch�@U@�u.�[5�K��Pn���� ���s��=��������uao���mo�5QǪd�?L�⧂�]D�G(���uO�!�'h�R�;u����1eH�×X�8}���Pk'$Sp<?���4�������␗�?_V�ĶD~�SO墳.�Ԯ�}4����1���1A�~(E�#�ݵ��<x�I,��zQq��+7�u�a���U�$ �̡	��ˍ�<󋪺k��Is��A���Rǰ5I"�ޙ3jӝ�DS<��kQzݍq�uS�C){�6y ^GEȏPdн������nz%-�N�J�.�*�z*u��Ј�i�41��h(�Ѩ$��7�j�Q>�1��[@y>���>����ّvXk��w���+�:g���5�Н�bB�d��z��j�#HOG�ְ�p20]Iܐ��"o�����t�,ܦ�wx�U��+��	���q�R��҄vѓ�O^���x����ڤ�5���Ɉ��˗��=B�6�XK��d��]�ו��$s�s��qнz_�qa$����}����w�c�)�K��+׭��Z�F����]�=Im�Ml�>�q4=�0��#{~�IQ;�Ԯ��[�Qo�:��>��θ�/L���v��C�em�}ο'F̳����Ӆ�B�iv��n_�ho��C�Ł�;�|\������V̩HPɹ=��7Iα�4��x��FB5%?k_ҡ1]�y;(�Ҹ�h�WR �PX�6���kї��Dd�����.8S����w�b_p��4Q+�u
����Nb��G�ֺ����*v�&�5����2��D|�Q�S�i~�G�6#<[��?��'�q�-0v
��?�	ģ�u��H6�.8lG�.�`S�x��s=ɝ���Ĵc(���ߌU2�����-���N�]�X�#�x=t��9�
x6ZV������u���3�&㛇U���rIaa��0�����'���&c�9�j���_���ϗV�6 ���
j��oF\[M1߶��|��1Q/3RN\I�`g��5���#k�Y,����b�Wx�/T����0ވ �
��'YK�c4�����2��9p�Q�/ �0Xfp�ap�!�pRL���x/������um��ޝ]5mg��X*��(�-dAu� {��b��,�Ŵ�@���Ps�&��ZkC�f���U�U^����p�ʵ͊8�����T$��Ү�����H�}Q�r3�qY�Jԁ�V5KP_�I�	��}�@����s"��d~t�o%��(�d��=������9��I輔��Q��`5߻^��Ȇ��7��a|~�&�~7N�>W�}���s?���s�g��+��� ��Ҿ���c��g`W[+�/��-63�[|��T���7�+ 5�y��(�{] ��H�Т��]f�)"��7V��ϝ���-&�tR�ل�[��=����烤�b��z'
� ��s�s����:����0�-��������EBf\Y���s��2���$�0[Dx"4�7�n�r5�5[���>�e@i��UR93��-(l��XP��5?�'ׅ��~������j����&q؈��*A��,��f�d�K6�-�xE����4�ϊV�f 'Ϩ���}͸�-a~v
��d��0��8ו�ѫ�8�ߔ�
����ks�X����G��Z����#�'�Ev���'�l�<dV��P'���L#;�,V;����g��vk� 3J��O����F�"z��G�8s��7[���J�1�����4z	\?����gx�a�}!��֭�9<R�.�H})Gdu��۾e�c��aK5KI
�dC ��c�n��i��e���盚�1_�`1���d�����xc�,K)�>�b�/~�ԕI�8�M�ۅH!���V�X6�����@f�b��o�̮�ix��%ϸ�a�����"�m�����F�ʻ��1�C͆)q�(����`�S��w<d.�6����`�����5>J���A��W9���@�*zt)��6�|S��i�1&Ō��\B�MF<�g���<���\x>��\/Wf=�} �� q��
`�J��#���M��c�:A�z�������_�V�k����ŢZ�ж6*�uom���B�|?�dj_o7)��D㬱!Lk�}�����.Z����{[�|M*��̗TY�j�+��}\V/�[�[сPE�
ᙃ��U�x���ӽuO6s'D�Qbg����"�G����F�E �u��j��
d��)���U�t��|�|b�����˹y8 4Ҥ��1>�*��(Q���#�/��ywX���y*iӐ�5�B݉�w�W���/�=����UOe�V��#�9�F�0�bVGzU����`��u��0�,�q=n�@��=og`�5�\��q\S�s4d�Ì��w+���#�o�6(�(x�szE�����R�Ө�;��|4R��v�}=К����p??1����1�0�I6�aŏ�Y�^��������vEZ
�ފ,��hS���]/_��fh�D���< ���B懃�p0~�g1�c�svY��Q��.�J��Op���Qָ��;(৤�.}V�}�H�M�����k���}�4M�`^�N]N_E�����������3�[m���ڳ��h�L�SxM�N���E�U��	��U~62��^����ĸĹEI<u��c򞉮M�_PR��D� 	����$#�`��<��C�c��7D�8��*/�������s��F?!t`7���A\W\9帙�;�!��{C��h���a��Ԯ}�I�ԛ�
��`�pM�9�^��&'����s-a��{YZ��Ӑ>��=P�����!�X�5�A�p`x�咮e����f�޿vnc�=5��i
�Ȣȸ"?$�փ��ɃU�z��NN��mA�:+�_��=БL��D'����ߔ����v�Dz�r,IZ-
��=��߄��z7�-�d����C�p۠>u��cm�adʆ�)V�i+����3wF%wTH���E���t]��t���o�E��]m���&�ŝ����bR�����}�4�Ji_��3��((���������p�M1�,r��K�'Q�h�b�H�k�#��N������23��cn��çD�mb�]�������5@}��䨝j	�$[��Ӿ�v��WL��eQ��*�����tfAq��fq����*��<�&$ӌ�B�N"}!�����Ľ�S����8��@o]�����7#c������)��n'W��dP1�M<B�
z���K0�^&����0+V���`��{�"7C#�gm�-՚  �����W|+�m�at��
����]�W�^3���ܺk6��c��u[M6�ɛ��������ea�v�0���:89kF��l(t�~��5�����3��K@_��L'�������b���˜���?h*���'�������M�)C]�7��Fﺺ�%�&����5���Ira�����$�֍�/=]��y��M��MO�N*�z��c#��n�.���jQ�4�\y���80|޻�H�*��k�Z_l���:��gPPQ�1����o��Y�����8�!{���v{4/hS0'��xy4*� �������&�S��XN�}s��K7���g@������<U�e�g���g�sƭ��WcA���kT[�R�߬]E6ì�������r�DC{�;�*|� � ����A�$�����4����pn���Q��).g���s��ZIg��y������XX��N��8ō4(�`�K�Xƒ���p�>�քi�PJ�^�|��%wl�����{U��ӂo���� ϧKz����B�O�[��]
4�'���W�*��@����c�~��9�c�*����6���v7zD�e/-#s���؟&ykg��T�+��8��!����l�V�Z	M$;X��)����1ԯ�N��:_y����'��k>��ia\X���9�=Lx��j,�,71�z�N�L%
N�-
n�h�C���o#d���������V��7U(�9w�:��N�n��!�a7|HoF��M���&RəR�[L!�JwTޣ���?�J�I=��>����J�_aP���`R�n%�c_��=8Sr��̎�ܰ�]~�3��a���S}��jM��G�����-B����
iNyGr&�ۆ�Z��i`5t��6���]�Ǌw<'l!�ű�W�L�e���t�	��bWD��y�&�����L��8}�Xʪ����q��x�^�:�uW��Ԉ��iϴ�`.?�M?#E�3�SD��L!g������m��P����_4o����l�ɵ��K2x��_3+ۿKm��(�-���Y�%��I��<^��8��V��;.�Ԝ>L�5y��� �SS���/�oY>�4{Y� �H=���Pe��|E��'k�+���{���|e^:kg���]�3�/J?��{@��O�Ѵ��]����n�O^%�t���p�D� ��f?ބ@��^Wr��n����e������7�j�boO��J�
���7��<�3ƥ�����.l��Y�t'՜��|7�.�D�p���E����c��}��m*�'P�̤�s	����Z+k�Np`X��7h܈Nsc�]V"�6���o�.���m߆�4_^ɭ]��!�ŵ<L:J/r*&�� �)jT�8p���O���o'��������
|HN�S��	s|l��������&m@+�$�v-ɨI���Y{��檲~�2�Y��HN\�`���9t�\BL�ף��E�������������O��� �(X��P���,�=m�v�W�b�t���J�a���Ϣ�T=��烇�Ǔ�x�6m�T�3�wb�~��D��Y����L-�Ƥ���e%��0آ$�$[ml�ی��Чa���
���#��x?��Uj���`�����OM�Z[�C����wD)4���X0����Q��_ ���ÔstvӾ{Ѹ�WL��
Z���%�+q)���g����?�Q���⠴�-ջ �L�uT�ٮ�q�X��FO���pu�e{e�6f>��+��(��榥w2�L�x�+�n;Zb��v �r��H�9��c��H�x��y�_�AUU��./@S#���<�TA�b罱��J�R� ������~F��wY��(�d��di���B���I����(�g�6�;�n��Ӌ���g��j���h�.y* LU:BR��k$�4�BP2i��=tSD��3R��H$�X"���Ƙ?�n�,6�?�	���92�D����>�#p�Z	?;����bѫ��۶�j92���C|��)�t��ӑ/c�'I#��g�.p(	j��s�E�g���p"��斴+'t���W�P
��&�cˈ�L�t	a�>Ffvc¹!���� R=iӇ^�8�n�_A�4��b]d��V�Kyd��(7�`WIL�ل4�ʍō@JfCY�Lg6[���V�[J���x��B%153ϗG�Llż�{4��_tM��,���|���aD�$�xj�� �K��޲V�Uo	�FǑ=������γVY`��p��n��J!�Ӷ<�����?���+ ��M-Y4�mqa.l��HB��g�`��F7�;s]A��~y>�A��u�R�^��ѐ�t��<�h�T� �%�v�����.��*VH�M��Lc�AaF����h���ngN���}1i]�42!�qk���������e���F�wp�e����n�5���j����ӌ4!J1�u`B���r���7���h�ѧ����N�����V��Mz@�ܗų��)l�j:�W���"_��d]/j>��#V��I��G8�(���_�|�6�$E*��Q%�-�7]��@��I�Π�D�s:ஜ�7
4�n���9E-� j��4�j��~O�:��=U�L�ՠ����LL1݇bɟȩ6���M4�УIÉ�� zp���K�)��� (B�0Q}�\��܎��.�
�����R��!�}C�W��|'�xr6��S���MZ��f3��4�q�$�{/�l�X�������i"K���3��«~]Z�b'�8g�L�ʭ�g+�G0&�F�m���ub{�{�\�MT���QZ�����J!��B��Z1��:��=v�:����5,����]���+e�����g����O������GA��(ؖ�~w�_r�+%X�+������O�$��坤/���:	���T�v���L{.���4��[[�z����!L�ؙ>!�0�hvx��S��4�K*�_V�[w���d��F���\�LU�}�����t�:��=(���R���I�D��r��-�����a��s,P���;�	��~�����ba~`\]fOV�ɔ����hDA\yMe�#�ߵw�y���5��9yav=,:�
�81�=�R�>g�5ɑ�������ѐ��^���a#/5�G�b �@�ե�֖}�1^�H�'��6:�W&�MS��A<���ML�G����;��Su(c���V���g"��R�kAq�!F�j/*d�%׳��&$7MJu�
\,Q*���5�2}Do5�Z�߰�Ty& ~��j����w�7F<�X4��C���x^q�b�5m��D�&�5p^�gj����#>В}�Xv(<��/�<�?O2Q���m5�D�����$����S�Ş��Q���)3)ɥP�OQC�����s���þ�uqK��Iǩ�������M�V���j�#���?$ٿ�9���h�d����o���r�%�J�Dt�G�,�g�HOMS}�����NDh��xp�^��J��E���U�-����e�Պ��lr���*�W��2s?)��)H�~q��W�s�T���a��+	�©9Q<���&l}Iع�z�a��W����~� �gx��W�G��t���P+��dB��es��	���N��Q�Ì�_=��}��!��3�U�?"Szc�13����	�Ih	�@M[��p�(yv[�=���'F�,1�,-d�*$%v�`�RA�z uTA����*r8!gb((x	��\a.���a&��)��n2����\�iOҠD@�a��1`7��#�i�A��Wd�9}b��M��CY	ۇ��<�- ܽ˳��6��������N/�8|�sX�K���(��UT�.�S'�S��|�#�J/%Wi"��0�R����λs��IY�y���␪�8_^P%���4��g!���)N8Iz̦������EU�O?��� ,�0�Ճa���ގUܼF��bz��(�@8	���ZO�2��+�*���FfC��_*�{��v��m�|��C9�s.���VK�8�g��of�֋c�8��VI��:���6��Fb�I��ȋ��@�/�ˁ}P����#�w�*�]8~�`e������[c��L�S %��g|��g�{h����=}-9���s�R����glU�u��*S7΍�� ��]��5�p
,�C�I���4"e��V��

�#І:�#fu#�E_&���z��mC����d`+��\���L���'M�}}��-��!��Y)�oX���pK5��YvmG4��{��<��/�x�����GXe�T��mB�8�&���M����oԿ҇>��F�p+�{DQ-!��B� �UM�f���g�BTXb�����ꑭ�<^��y�k��/�1���i���
��5�&�WuIB��u�_��
 ���;��m:��=T�]���V��&"����Jn�+�� ���:��N�awk��E����{��l�(��'$̼F8ba�i�K�P�3��u�������5�$d|m��=~l�4�-����	���&�W�T�N�-M^��hw���	&�\h�W�J�y�)S������'�W~+b��y���Mp�<{��L)�l����Ag������N�D1��k���[0^�'lt��'-���.�
���g�hgU���l&a#�UPM	p���s �r�L�?�r��;I��r��*;��ٗW�����,��CnW޻���Ȼ�ȍl�K�UӀN2J�[vn�3�������I)=��O"��	�]R����{I�I��O���/�~���.�|�� @��*� �J���;�;`V��פ�Ek^�J���ٞ������e9�f��a��GUPp�q�H���Q"��:\'s����	Lc��]��e//�ê+	s�E~��L�	.��u��p��;B%�����f�9]{���
�=���� [+Dv��y/4����h@����|Tso�V���T��{^��@�)��9W���K������1�����d���ȮQ �{�����D=ܺ�r${��d�)ጼ&:,L^Ǵo4�0�,��_d��h�{f·��q�ۚ0��S�Z�
Nf%+�>͋�fHz��[7�;�T�f׌?UykbS�lJ��������.�t��J�`J�ś�@=�x~b�13�K�sw�u�䏾��n�Lq�m�?�2��s�R�2U�(otj�"|����c��;ly�Yɬ�{=�l�A��y˾�0S�~�t��S����$ܵ�fc*���g�XNu�j�=1�78O]w��)«j��NT|R���j#b�TeG^�+����)!� ��KSh�8�4zb�,�dh|䧳kޱ��2�FK��	|��O��^�>�����%�M��2_)��[	����^5?-��L y�'�Q��^�)J3`=]`Q|�"L�!� ��0WU�*�̥-.q�h��6��$٤��A&��V��)�%��(Lע�Cx1�����WYϤ�
WmB����?���Q�pU�Xe�{"�J^�_�D���<�nOao��x7��H�����=q.ţ-_�=6���N�y���N�6��K� ���
�Ძ��2h�rgC#�%��[�<W�4�W؀z;E����ݯG��eU	�in_^���&��8y�Q���XU��t���J��	Hdg�
��*��燕���4�6�����o+gF�6_��5 ����fErae!� k"����$ serr�/�f����a��U�i���=�eM'UǔaIwJ����Ia��IΨ���L)�ñ�������#뜷h�frd������{�Zڡ�K�eD�	"6t�/6&�� Ր�<�^IDgË�/Y
D6��qy3g6@Eq�w��_��6w���sB����v]K߀]`�)���������T�JxtEi�-���-��o�=�V->.P�o����q�#�����{�e���r3�X��R��y=�޶b >Nw�,�}.�{���C(��~�:���d2�yݠ�ʩ��}Dt��/
����ܘ�	��?�ւ԰��㶵39��W�. ���L#�ב+kSҭ���~C!�#r�N�eY�����*��,���H�qQ�d��$`��fGcs9�OǂR��῭�Mvް|3F�U���!4�Ʈ�t���DH3&��#D~�94�|�&��ܳ�,���(����ms8��!C),��x(�f4T���NϦRr�vpI9��i�D)i�0P�|��z��*2-��Ҁ�^���-��:��if3a��E�F��{�!�u����<�
�n~���v�p����ZRC��a�
i����Dm��|J�u�n�n��=;�RY��h�t7v,ǰQX���e8ue�be+��8��St&MS�QGn���袙�O�y`��:�o���>7�����S���8m@�?���z�k�j"B�C�8�W�*�I5VS��C���x��Ե#T-�����pge[������5�<R���3]�Ⱦtb�
����QT�J\�9�c+�b8��W6��259e��
~A�����zJP	���oYG��V�\�'M�xs)l>F���W{��p��|��L"0�jO�m�N�e�
+�Tk���,��"����u��-Pb��S�.��^ĺ�5�ﯟ�:4���	b��Q#BO��e�O:��l�P+Ͳ�eф�OC�@���M����N�������ON���E�4�:�TN_�4����;f��
y��,z�l2��u�mJY��_��Xb[�]�!�U3h�,��z��q�Y���0����!7b��.���G���6�Aǖ!	km�%�Ξ�d����C��I�1g����e�YN���^y���dE^�\��B�J�lU8@�_X"_��b�d:µ�jh���K'f������09�tzI���WQ�Q�ȡ3��Á�}53�����4ς�2�f@Z���|6�6�6�y�"�3��p 32��@.����h�5W�[#�a��A/�:�J��2yd&�R��Lbw��USU�����{̛IE&�B�ͦ�|ʛG�w5�rǙ�������g�"��7�jp
�R
���I��5�D�<��Vz+CF?y�2w{k�zfOwJ�?V��S�����8|]���& ��Ǿ|@ӑ�'�q�����f��E0%5O��d��V�����'��5+s��'ܣp�; �M}t�ݶ%��R[d��5>�̰��O�)wz�i�t��+~����'���{���=�4���w4�LS_=��!M����B����Yny�oB���!�F)����;��xL���3ш�������*\R���*�Fo>-�3�U�B�
�0�o�M2[�%��FL�e�8�o�cBw�[2a�
k�5�o��`Sp39\��+�!�*�v��Gy]��y&�eCefC�@}�y���3�b��2�2����� �	T���j	�=q�[��GX���G�_⧿~(d�y��V0��ǩ�3��R�r�!�+*BCb�m�9�m�{)¤�1����0:c��P����'���	d����l'qf�Q!d���:�`�W�~��\��L���>���e�SJQHv˞B�e���9�t����Z 6D+��p��B6�ϡ��)4��A?�T8~�$��1�)(3h���� 3�N�����^��ƶo���Z��$����/�^�S�̅+yo���d��U�Db̽���S�`�Ǐ����;4dl��j�e[L����
�V��-�T� ���G�lJZ=b�l!z?��pF�A%X����}B�ho����Ң?�L��;��2}�}A�&�����ƌ*�{�_@�,8�qFS��r^�f��-ٲ��;n�,�>=�$��1�8g��kFYf�om������n~��"�����a>�
�#k���qD��Vħ�uv>QL�w��Q"����!4��2��.�^0��mVd>�$��ׄ|/(I����o��k�aNޗ�>?U�d�/wg�u��W"����(��b<xx\���:l}�xstr)�D���*iE_���4Q�����]Ȗw��'��
A+�c�7��|F���-�V�W�ra�5hđlT~v���^ԏ_8��=�?H�0�BK�Q*|�l��s��om�7��S� �M�ɹ��\��E&~��^�q�^$P�n��c.�eY�Z�qk�o����!��} y]2��u�CW���vZ�[FE42���hE%O5�-����?��+���߲|����5(�Y�<	�����[���OU�V jdGъ$��4T KV��n��=@M��+��B��R��j���޿H�2��sH��W>��&n�^�is%���(x�Ũ�ɚ����/�՚���7�o��{� �ӥJ�FKk+ۮ�)_(�nv�WC�y=��Զ2-U�Dţ�{�*eE���s{zD��;l�$�<����ֱ�}�&��L%C�
{����m�C��Q��M�%B�)3�-g�턬�4]�f�Ҝ\�i�s��v�ݥŋY��C�B�-ϓ�q������l i��烦���9��YP�n��b��s� �K/r��N�5���Zp	��X@r2��( ��x 0)<�(gM���f	�`-�b��`��<Alx�a�N�C��E�i��ПO��W�թ���^�r����?\)�~�=��-dW��)��V�C��#�h5�=u�;����Llț�F-#^D[�-�Ui5F�Y�b��Оby� P���S��ъ2o"�p��*2g�?"Q���ˀ;3�2sj1�Z;rz)��2�?�����'�G7H���Kb5g�\T�Pi[ߑm�$�q���R�_G��y�^ߘ��]��$H�k_i,�I�ϖ�hq�M�[MgS�[/��X���®�jn���u���8K���+n�;_�ձ��\w���:� �f���0��� 9���N�H�
�a�հ?�-�{�n���n�o��t+p��f\�h����A��Ӭ{��D������(eͻ_��a�@�v�|�rl�SL,�d����)�&�⧟��G�qB�'bu�S6b�$�`0�4�z������~�EAg�+���6��uTĜ���X�p�{�O����x3��2�:S��bs��ha4��� �����:U3�\��>���z'	�"ҊJ|�rlq4�Rn����9�x&�Zoڏ˩��By'J@����Ʒ�2���͢zY�Y^�u\�G�����3*�o��Yϫ��
�b��&��vϥ�$�7�@�0Ȳ��q���wE�56Wn�I)�������2o�<�X���Y�8��3*��i�:<�B�|��6
P`nU�崳4�>*�A��^�	nXj�eJ��}iA ��L�܄l��jʽj��,Pa�;`�>Mn*uܠ�VaN�[�����V����%<��GJ��s��a ޣo��RD6���*��G����s�B
_OF�ؗ��I���?4]oڪ}��U0��?��u$�ш�5.����u���ԩ�6�(pu�`�D������0��i	�%�D1�����ÿ��V���W����\�0f��l�7s�?�Y=�͙|�%wr���W;S0�C��a����"6��J�
�rv�%
����l�u���� ή�cFW1�dsNf�U��d����"�y%�9h�-�|�VY�����}��z���N4��1)w,��فl�=D�}�lW�Wa�M1k���O֬A�ׅ�]�]�V{�r�[��W��)��g�8�ʹ�}s���ڔ��X�E��5��,���U ��=�ZyC�Dȭ�dZvd?�G*����,���7�O��-��]���A�2$��4�3C�V��bPL���N�R}Sk��#Ռ�"º�t+9ůޗEd,�x^�
��
��X>^�C��k����(iG�	/sݽc��;�8[��{��_�Ť�/k8Am��e��Au۝�^�~�^G|��s� JsB��c��y�)ݼw� �ߞ�eN����'7�����eh|��t��� �MơR�Ge�)/O���w��)��m�L�u<��ac ��lr��i,��a��:#D�(eҥh���h3�������t�X�VCl���x59��|)+0c2�ǆ�i��"�9�POW���j迕��-�̭|���'ZF ���4��'I`z�V����ʳ=r@����l�2.��ł�� ��h����2��4u��X3��p��pV���x%��`�$~��7o�l��F<��ɚh|
xx9�ɭа&�`���O1�xF���?����2�Z�17p�PvI�)ݻ��{���k���=C���/���ǯ���׵܀.�Z����-?�(���~���_�;IH}�j}l�)2]��>���A8�Q5Dp���,�#��ٯ�m����,��Afd*�&n��X���n_�Sd��N��R]D��L���ļn�9P-�>�P��e7�=F�0�#v6��U���<�S��:s��������	a��<�'�.,~hԴ�����Ӊz�%��XY4��g����=uO(sg꠮�ub��� ���2YQ�ʞ�����ר�+��F����FHU�y��3�TuL.%L�<�?q����Hc���N���Aͤ��vn�J�7,;�u�(�y8<�����f��$*� �5���o�`��>J�5V�;(�R�v�#�<��Q�Y.m�h����(������}����S��Xz L�5��\W�x�H
竲C�H�+HN��oW��h��eLg�6��jS[5}���z��|���7.�i=�7��L��չ�R��Y]N.[�ߙIv2_�,KT���)��	��{�z��V=�wVa�aq�F����FJ ��n��Ê���2��_����}�U����䱒a���Xei�����E�~����S�:��Y�j��E�I�� �Ο���tA��Ȗ=�<4� ��m_�t�G�r�0o*d�Y�,����m՝'}��22ީ�a����w���䗱n^��W�Ug����p�؟�!sݮ���m��b�ʙ<�|�Q�P�S⹍k	E\�Y���kz�y�>P㧾��������z����m�͐��w�>L��KxS�q�mL����th|���R��L�=oM�C6�����a,��b~�K?YzQ��c��	��x�\�J�k��3E4�f����F�U4!��^�7��`�I�w�'�~�	�1�X�=	 {J2X+�>��(���S�9X�{���ݠA��"�����`pw�:�u�6!CE��$2�P��}�W��W�ؽn_�C��`WGB%8���F��/�R]��LQ�]��<����s9�k��}F��_o��2cb0�/�Q�FD�F,^��,PڨB��l�5��s/����@o(�a�s��_��U��:`<�U�k�侫irW��֢;F���Ղ������(���,h�qѷ2{� G߇�|�k���ƅor幓��tG�hp�jq:т߿9�u�2bЉ>�3g��K]b�z;C�aZ�� �KA�e�ʬ��<�C}! �<H`�*˻G.�̙���� ���nN"���*k��ޯO�*E�?O1�v��9cLk�+���y���nEi�R�F�mO 㵥�Q&��to�I��`'r:��H�_���F7��)�U?Ճ�KA�A.~��hK_K[v7���WW2dw�%-}bS��΀ �V�Qt�!�*���g��.
hx0Lp�x<Nw�"iF�%��T�7p���R��Cu���{�P6 ��48�X��|�JR�F�%\O�LJE�sG�0+��e6�:�K����.�Zu��A&�Hө�c��������?���9�hc��<�I*���>�����a�w�驧RL������	QJ�%,I0qSX�R?�}�Õ>� ��?�u{�n��fR&��eߛ
�x��[W�@��y�X.9�c�m�gw(D0��c� �j���N��������g�ر�W_"⡟N�*ܺ޻���KϹ		���V� �zQ^��Wfd�&w
�R����.�g���� 1��]s�mҗE��.v"U��HzB��,��"��"���݊&��W��iF�
������H�����;�fPpB�s�a��N!_zFb^�~KO "ƫ���V�Lw��h���82�W�*>�� �'ߖO�5<g���ՙ�RT�"�{%M�����6i�<:ڬ�BZb;�0�����`�Ci�<�
���"���R}���#��b�T���g-oPխ�*�j�w�%Љ�R�Tny\IA�xf�-�s�#�}�����S�o���,DNj;W��>�h��@�'cv.p��?J�h��8�P���Ri'��>��#"D���5���ߜ��W��n[��J����v�a��")ռ8�OQ���y3�����JegU�n�*.Dv^�G�Q\��ʤ� 
d�tΠJ?�l���zΎ������ (c/���������\9 �1���z �e�Vr2[m���%���g;����� ��T�.��!dG�1��C$P���T��KwKv#ے���Ym���u͵��(�@�K%���I�0��pt{|b$ ����rvS�{{	y�P���J��0����|���6V�\rȿ���K�"O��ʚ��b�=��.P+�O^H����^do
��?ww�/\�ӌ��	`�	דS�ƢS� W�x�) ,0�<q(�&��%eQ�1��p,ժ}͊�(�k�3E�����b�-��>�7��S_�k�@�6T����hA2����j-�C�w�d@,�#�Ύy�=v��A��j5�U4I���������
�N�m`m'FA$&�?s���e���h�J5��l���Fmn�f�z�@SY�$w7p7��1��e{�p���{�G�0�7��ag���ˬ�o�f�q��Q��g��f�n��p�iE�ؽ�?σJE��`޸�)�{�w����3���C��Ӄ���Ŝ&���e��(��eO=��M��L}�)}©�З�]��V��U{Ǜs1z\y�~ p8/���9�QH��A
 EoiWl?�*�\&�J4� 3��t��jst��/"���S�~�T��IB��Ru,|��'�����>,)��ע��q����?	Ό�5!~��;�k<Iŭ^$'� D!4I�	@q�E?�-*֒����)��I'����&,�c�����\�(���FA�R�R|��"ʀ�cs^��.���=S˃L"�iy�@���!@eY5��61k�ؾ�Pa��O�	��n���O���UC�7�`c�9t_[��������7�I�&�b{�p��Z���]�ĩ�.���d�.hr0�uN9?v\H����d�#3O���>�D����U!��:,G�.�F"��n��JM�� ��d������d����i;h�4_(`�}�)�����
�C`��ɷfm0PRI0�{E#�NL��j{<��듩+v(�T�o�%����-H�Գ�J_��1���D�Ĕ�BRh��}�����8��F	�>�	p����Q�po%�}��֖j���&�t"�?�E��UW�g��Ѝ�l%Trn������!�d���h5���]ް����p�ߕ���ml�4����ٮ�0�X�����<c҉C(ψҕە��n85��.��+�}�"�U�/K<�3�`Hg��hnY�h�,���x����h������l�܀���Ǝ�Q�%'����װނ: ���U�QH��z�����j!��:�'`�3�k���LeC���S����P{��rF�L,��q1����̗�]2@��j�tyg&����ٲ#�
��8AI�t�]�X��%[�����s}/7���
zO!�{�ܧ<��51Ne�z��%:g0��=��(�`n*S�P\Aq��`[%$X��[�Er���QT�����|�/5�x�/�}M�l*��3j��2��Q����#�������B�c's��y`/pD���ёW���gD4r�!���ͺ,���?1N���[�_��'^���k�Xx#
�=�*�	;����˝���A�,�h��� ����6N�nQ�z��Yl�܍D���_JѮ$���!���M�(�R�ë���v��lG`�H� 2�y������^$`�|_b�iQNy,;#V~����|��UC�eM!�X��3�o^�@�[u��gJ��ez���<W�)^VR��qK{���b�bW�^=׀	��x�Q:Н�f%b�+��:5�NZ��"�i���7���&��K0:��<���[WY	��,�P�_��f��h��&���޼� �8#�n�pJՇЁ-��v����R=���@27����"�`jn�e: ��g�O8i������;s�����Ln�^0,�{p�9c�B+����LJy�詎JLۄ�:�7C��
NЙL��)+DMF��q�gRS�w��q�eo"�cvה^����@x����/e�_t�Y�Sg7̱�������dFY��N�����r���[�c.oJY��C'��z�"��I��*68c�n5w��Y���:b!|!��)���ױ6��	'ܦo?/�a��O��b����9V-;���O���L �v��r)s尡j�Ҵxi�8��G���Pdї5ĝ!2����g/�b�Hi3�C�:|�/�sN$�߼KI���OiX'>%Б��������} 33�H>�S�.��#�16�r�Ux100�S�	�Qm�Ef`� .4�?�WjH2�$��	<k�]/N�/��<�RDsM�@��r;߃tj}��Wf��%`V��^OL��/R��=;9��'�̩)(ˠ��Ɛ�x0t��^O��a��R#*�Y���.nZIjpk1�?�[	UW3����\�X�!�I+H�R�wCѸ��̭��Ry�P�3,�,������'��'�7|�����L��)�o0��Z�?6�pb�l(���ۥ����XXv�c�:��Q|(��a���S�D�M-�4��u-��v�$��M\�����k�cG�QF��QN�tc��o��D��{����++&Q���$��h�!��&22z�4�(�ۡT�u�!��vw"��B�yH@q�e�2[��֐���^ng��aX��b�o�T�Sj��R6d,Ѵu ����u�2�ZDp>�)p��H�?Ne9����+�6CQ�Y�ر��3���ā�؝��X������t�1�1yU�����->k�ы.Z�>�S�'�:M�$�} s���و��v2��~y�`JW��O7r�b���O�1(	��*���w��^i0 �g���"�	�_h�_��q�#�"�A��6n�;�C���g�x͖�5����Zr�Pì�R8L��=�4�f���݈�S񲽒x�i�WAcP=+�+*E�F ��,K��"J�(\�1�T��QN���"[��!iV�k�FN�,�#3���[�u'�	#�h0VI9f�9S^�ۙ��7��/z�����h|���V�2���A���;a� �o��6 	�w�03P,&��Cq���C�,�Mq�9�Q�'~j���������}��x�/Fz���<ppj�Vh���_;�������}H���@\zL���Z��%�$�g��0���5���j&Jz=������#�/�P��C:��4�5h�����.��ou�s��*4��S�_s�M���^H��Au��Ch�������u���	�s[�n��r�o6�k8n�@�}�:������4�)��M(z�Ug�T#o���<L5d��r��>
NI,�pG��P��)7:�8�B����d��v����^�3�0_K����e*���46���2)F�4���q��T�6�J޵[�+Z��ꦸ8�8ڷd����ct]��F�IwH�Ye�q��T�D��hqpK\^��G�9�����!��KR8�'1�����5�'h��1Ҹ��dtx�`���p~~�3����6��{�lb�&\��u��˟t׍h_}v�_fSZ�S�	V$Z�_�l�y��Kz������$���3LC6��@��큋���>�4&P��� 0{cv���
�|Yq���l.[ط�,��?��~*�ۖ���}��{Ӱs�s���3z��!�yg���c����J֦k��`S� ߼-r|�m_Ҭ̡�kU���B\�m��Q�l2'�2�4}�m�PXc�j�F�q��ş�M��k����r����H�%�"X�`O_&��#zE���֤+"�Iq#�R(żG��J��p��h5���ߥ�-�/�vA ��0v�(��ַbK7t�?�/I2�xc�R�qU4o���%{�����l�Ҹ�u��r��|f��?�w��yP���{�5�/zS3�'��X��I�x��x�n<�y�K)�)7M�ZoUfe-�bZ�I�׼��e���Q���yWhl��彘���fP[_��^2no&�M�m?�oJL	��
�A�ڦ�˅�#�����u�J��� N��2D��Uߎe�{EDY	X�V��=�#@!�*�/��:���pX_�Z�@���(2�e�}�t��v�I�m�?af��yJ���a���Q�D7����4UG����ιBOX�#��a��5V��j_??"�$���;������>�"�9�b�\�+ٵ�e�`�x�;�+v�◞�S��	���1��y��Q}��x�U���e�)�����1)+�-7����"�ȺhuA�W�3�!�@�+���=@	�?�Qh�v1�H��N�iUj����ڪRK�FEJO�=���K�FQBP�|J>�k��L ����V��\��gգq�  [�o7� ~Zù�m��������0@`$G1a��S�HH��=�M7���,2��6�/<��̗}�^�G�-�\���,S�kl/�t�ߍI����g�Y50�҇ƪC�kA]�2r�:���|�
��V���n����>�@[�;��ۑ��ܻ�t�8��́�E]�N T���?�x���N ����-��0��d��=����?��;P�	���7$�N�#|���݄.@kz��2��n�`�G�ٌ��}��D;��c�h�M��(���7J-�*�H�&qk�2K�8����y�N����t�N��˪���L*����n+	Յ3l���~^l_+�.��mh9���d<8�P3UtY�.�ܘ�����M�5]�3�^�Q��^B��R�R��"�0=�#̧�ꊀ��w#N�W�_Lӵ�x�I�>���B��%��<Y�9�Mg���z� �R<��1��o��N*��l:�w��zl�H�Ƭ��<�纛rׇ�3��z;���Zs�_Q�Yp�&��͞u[4|�;�SR6�����0n���UJ�T(�
�k>=�|��' ���#)2�.��m�Ob��82�&�a���M�D��YN�-�h�lT���f�Nq7���/g�G�)�#^$4�ZS��=h����h�f�?j���*��m�x1�[�a����0Ei�ٯV�+x���q7����qW�W���%����2��ml���l¨��QO�w����f�5��}��O��]����5�(mF>k+�}5j�;�|���p�ʇ�f��.X�����;��~-�����Pq�e�fz���a� VCF�J�5>��&пiҮ�)P*��6j���y�z�w���1&�����
K�֕~p}E�ĻR����c���4X�㄂#_JmcNć�����B,���b!_��Y�*�E;�K�D�x0�S�&۳9,�yyI���w���$�?Q=$F�[Yu�ğ�݊�X
�Ӏ��2`"���.��gp�}����z�$9q�lD�b��5���_�/�X�?�<����hU�|d�0�t�i`]v<���D_TT��p��T�`t^`�C �: �E#{�[��L�a�$�}�\����2q,�`T��[-��V3��]�]̗�dȓ�nz;��j﵆f��ېvi����{}�z{U����+����_����BC&5	W.|:DK��t���ˏ��Lt�q�NT#J��{����y͹���߬"����L�*�ym�[��j,���� �x�`\�@�5����6�������4� �{�S�_O��报]5M7��#R���w����O=ܭ�XVݤo且n��<#��_X:���e�"��Q�^v�T�6erOpU���Tk.��sc��*tE�&-ʻ[���X��{��*�Ĵ�XW��*����bՏMM��Y��yX��<�t.��o6�d*���i���߂�b49?�Qgm����Y���Ќn"��^-O��Ne4agL)�Tg0�X�h����qE,� �em��������#��/�����$�˲��&�G�[8}�t��M/J�
���m�����l�r�4<�QgH%��$����&	���G��6�͍\��L/J�?1hr�7}����*�����"M��+�X��;�^v�x#?B��7d�T�� hJ�4�0Y��8z�⌓$O�G��A\�Sr��Ǝ��=�_���֖�~��By�;>�H	��Ӌ���v�1jO,�)42f�+�t4m�zIX���]fM�X�L+̽/y�03c��̩au'�P￦ԙ�!ڠ{���;�5�ғ�E��f���M�O����4�WIJ"��i!�k�}
Y�������L	v��F.>��j�?�[H�U�j�G;Z[�kf���%q�9n�����5�4e)��OF��9G� Y0�a)�|�ۄO�]J��An+|}���HߣACG�����zɯ��6��R�1�fu,�"}�싶A�K���ŊT2���͚�Y��>5JJE��Z�r�����U����P�.���������g�"E��T��a��u6�3	��%�Lq
v$\"Ĝ�b�>3%X7�����'
��@:��~X�v�H��\�lÜ1'���c�Xlr]�J��]1s����U�k3^�����Q�qe�Bse�M�;�(Օ%Aڬx("E[��Kb��]� ��J~Z�:��X�O�{� ��PM�;��"%֣?�"n�0��⾷�N1M��S^m�e��T�+ty�╮>��bѮ$a��/��a��*��F�.m���[5���5V�U��@�ţd�6���>��|����?xP�m22d&���h/� �6�<�Vx�4`�ƥ�CoH�Ժ{���~��S��h�U�`�
����&M�*jYz �>8�RZ����=AYY&�����C��P�wZ��>�jjʪ1T��I�t�p�m��^:Op�ʸ�k+EʘS%�M��&�8�L/�d������ֆ�.H�ީ�Ɩ{���<t�P��#��>��Q�cs�}ؙ#vs$Ĭԙ��o��N��эCYS�����\y�E��d[ԋ/&m���G廝ؓ��}��S��W;��q����\Gg&6���K֬	����9�]ǧ���x!VTڭL5
�&D4wǖmz�LÑѥ��8��l%�1�hYC`��6^EA�L�|%�.��_x6� 5\���M��	(��N�:�=}�g�5��h`qX��J�����-�
!�����Km�+��5T3r�,	� Ύ#^����D�b�}u�"��M�Dl,�o�K��G������@~6�:Ty���!)�=�>+�)�����&:tÈ��lu#�b�qN=��u���55fw���ƌq=����+ouNҊy7�ا��V����6q��[�u0"�!k��]�� �9s2�(Ql�7S�j��n��d��*Ҥ�_����!��K���H�,����=��)���]4"��7+E��U�JO�[�~�ne~��֎�6�d�X󭴝fW�D8B�1E�&ϟ�������
�����A���z�^4���u�����o��\�y����6��۲��%Kᨫ͍AP���}��$�����L|J�-�S����%������+z����H3 r����d�8�v�P�sfW���ǜ���i��R��j�\�c=���⫄�x�3�ng+���1 ;�1"&�����%�j�z(c�u�.�JA�O���OS%��#Ͷ�e5BK��@rm~���A�N붌Ė��3ގΕ�=�O�\oխ>9�?��/�a����J��A8�ɲ<�z3�V�5*������v�a��ݨzm��~$q��fSH�ָ��-MK��g�.���>�+A�h�w�oi�/��ސ�پ���x�$�Y�I��#�|�|�#������"�>���t�������9���cՎ�'�7�;8@�2�B���2Y�Z�_ܤ�Uo�ƄU�z�,#O\3�������)yt�Jz�T|�$��VMT
IeG�M��?G�~_'�}3��{��^Mf&�����{�}��h�܍5 Zr�Y�/���1>LS]�ZP����\�
�e������!�t�]+cV���BZ�'�)��ɑ\�:O��d&*f��{���_ʍk�}Dm�L/�QF�eJ�+ݗ�;Γ��ٴ\�G�bnR}-�I
�S�r�
c�Y�����Ns��2[���z���[�[&�8T�DQ�O$z'sS��_�2cI&�e�.����;R&oca�?�j��UL{+����ߞ��������Z<;D�GB0t$��;�4L���Eң�v^''s`����=a����VX27Rﶾ�Fƪܝ�5��7��?iT��l������ڥ3��a������Gü�B�|c>dK#��V������"tϩR+d�w �>�Ɨ���2�"X@,�`31D�\t2�ݏ^Ёx Ӭ�����u (��9���<����$�2����!��D�&�ȧ4Li��)�Z�ʥC�*�WFm����ͷ\���R�Y�CBĆ	F�G��Cz5h:��:n�lP����c��FQ�?C�p;�U#w���V<�����Fo�#vMk<�Z,�U��K��n_�d��#����3e�&�mH�B�@�k����I�$%HY�~?�����ٞG+{��[(�e����b������r���ggC
Ɩ�s�:]��G�vW|�&?��EsM[��es?��])m�I��OK-ݯ�dͩ�V.��*y�a^�br������[PZb���ݺZ0�m��`���Q�� ɐ[���>�Ӄ[��
�V���p-��y3{I#+}+�F'�lY��w0��	<�c���DÓ& �����'�p�����S+��+����3�Qm~I	��+���ɷ�7��%a]>��v$��:�Qͺ�� |�y�z{��$,�����sO���e�$�J�U�i�����m�F[�'V�D+- h`�H2e�W�5�]�m`���1e̚=������D� ݓm$@O�]�F¾���ӔY�^��-�4��:��Mn��+ȏ�U�b�J���★��2Wʌ�g��vmڮ�َ�Q������^c�r����5n Ӓ�E+�Ԩk{���nߖ�-�!�7 ��ќ���b����i��E�#a�B�U��%���Ħ\}����1�U�8�8:�����^���[y���OLJ1���K�����g�V�E�O?ȮiF���۷�׾8P���[��6ojI�a��V�眜�]���YAa��ESQ}��5��\�M����a����kw[Bc�O\�W��L�ёoj_I����6cd�G_��73�ʡEgA��x �����un����1������qP���T���9����\_P�;����<�x����N-���,��t�y�>=�~I(^�m�1�C�CcoD���`�(�V���3ppe��}Ⱦ$� ���!O��Q��2	m(�]��g�"A��ѤY)A	8��-+��#�M�=L�i��ewr,8N���LZ#��dD@�PU���H@\T���VwV�]���c��s
cK��������.t�u��t9k#�v>��gC@wN	�O��!���[���؜���b��_u쾵�?�z��-D��j$�,Y��)d��x�IYQo�O3�e�T����`�HVa$Oj�]�d�E��4*�3Kq~%_Ӽ��l�M�#�44�!j�&Ɠ��m�r2�hG��a�S��J���V<�*�@AH�ľ�7-X8e��Eݞ�aQv-?�l�gg��W1B�Qg�~� w%�A�lx"m'BM���q���,��j>s�e�~u!��f���6��<�,�魖�ɂ�<�k��3� 4�G�u��mڱ��f`(��	6���������������'譝�t�Ն"�bA`7x�&`>x�U�eG����A���,�9�����S`w)��q�Y�������o����S���M�C�>?zm�P�yY}�U_�"|K�ܚ0	w�V{	!��D6�� V���Y���ܥ�}�
Pe(��E�}"ן�u�Pj���Z����T��n[e��B3��Z��� ����P���{�o�>S~)G.�t� �=%�5�];�߳M	��h	�+�C��ۖa�i�htz4�٭��<�>'�o�D�P>TUS�����U���@�� �e�]3�AV���iQ�K,��+FpwIb{˻��-��))�Ng
!���A���d{"f~r*�mq�N�[l17��o���1»�O_fB�	��	�)y]6#A�C�jBJE��x;m&�zb�o��u����k�>s�z憒����D���j�ôa�۶�O��-��W�gRUDL���$[ �q�����j��4`�^�+<�|)wC��)h��
�#�#�:�P�dQ��/�w"�����{����K�=����x,ޒc��[��F?bt&�����>�LĢ�i�/ �>�
e	�@��0*��r<�\�7�}������.�[��ݷ���Xb�C�՚]���U��6x������hp�9G���i�߷����ج���j,Mc��5:�M��Bv��~�����"�3r�J2�_��M� ��h���Q��g
�<&�:������ޣ �;��ʼ���4$��ց��ONAH�gS����.?�@��R�"��"���t�թD�z��p.�K8�4��C¤%$3a�ڵ�97D���ԭ��{��q�G��dF�,!�e�4S=4�x�Y�n@�u�<C���|�����{�G7��d���谞��P���P �.�D�'ϊ���؄#4�H���[s��%:� ����^C�
�e��j�FC+E��>��O��V��n���*������Y=��68�g����'?Q��=�+cܫ�F���j,c��3><[ޭX9{�Q�Q�~��ց��Bli����@-����
�&�e�#�o="R �(tV�͡�%y�<�ֵnZ��l�"%-07��|4h&���|����Sq�d	���Z�� ��c�وcc���1���� �u.�>�>Z��ڌ9ٙ�|"�:��f>���j��#(v��¼��FSj�B3W�����LѓĹ�WN�W��X�@4%˛����������@��T��	��M(�v�jbl�j�	CsNj��S��A�₽~fG���g����]qk�����u�d��ݗO7�)���y��j����˔=  ۛ�+ڻP@=����⮷kЂ�g8M�\])�i��oB[��$�yL����P�WC�n�����L[^S�\f�V�`Ԣ�8֑ƚ=��ƋSV����YLrG��4���/H/%7>�G/|�p�r�1̡gK�Y0[���Q����:~�o�[֛'��.�dcS�����Ҥ�n��<��(��������ޅ������OM��G�0���èu�6�5k����Ƒejv�!9v�;\4��;o�`����|��m�#���/��D#5z^v�.��e�\���n6:5.��sr���,ܥ�L�$R�爊�V2h~������@9�����y�P�v:4I�Yv}��[���8�4aq:�,����
ή(�����mo��1����[�s�-���l�V�+q:�θ{6�	�H�h�;9�]�h�k�bt�y�� dN����Xw�� �I#�^+C$6g0�26��ǭ] �*�Jx��/x�d�"��0AK��C� ��u�~�=6�L�j�����O����'��/�x�����a�_�ί�Ҟ3��:��1�=�\`�XK�J��鋀Q5�vw�}$��ʪ��^���
q��Q�=}-;l�d�Т,���xH���9��E��/4�|��?+�B��,>�xDXw�K�����f~��i�$���r�?п��F�A�u�� �������0�N8���mm�b΀-�����_ʹ�p��E�� �7�M'̽Ly��8m	��d�tz�>���D��j�6�ea��PE�Q�i����q�ho�?/��ʹJ�o��FD�c�t�<�7Nҡ��*�����syC�]Ďf��.�mtN1�-��v˔Gb�u�5.�LM��Jܣ��E�u�1f99&nh틉����6����� �1"��q�t[��FP��b�+�'�w�/���<�f�Mm��^6#��4�M��d&�*	�~��[�hۇr}]˒eҐ����{Èξe k���f|��ń�R�;�n�����~��d���@b�ｭ�&nX0���K{�Ԃn�`Ж�!���x�
k{�W���g�/ҿxV�.m� ���Ǹ�D����!��[���j��Ke�ή�"�_���)�7(R �&3̭PJ��k���\n.f7�'(*�.�{�Ek�(���:����lb����Ise�x#���A�i��y�$D�(Ж�ύd���m>��cǞ��~���m�<yH�.���yi!�%g��O=p�q���)דЀO�p-.�eN$;�|S5V@��J��O��2�z��H�+��Ӛ�"�M+Ħz�L&�J4(�q��<~o�AI�� ܖ�B"�h�c��Q�G�+%�s�$p�&��q��͊m ^�cPe
�X{.�^��~L^ՙȬ�5��.t
�n�7�5�}e������*g׍����݁&mk�G��jt�V�^qޠ��>�z*bW�o K�(gK��4�O0�w7��uViS2��Rv�{�{��U 3�>�d�R���0��"�*����~S�}�uk	���d� 4ɒ�O9��[��I�L�Ӥ��Gmȼ��dSs��܄gmSO$Y߉���� 	���[k .w����Kr^��L�-+k\ǂ.��rkv��4�i��lh_��x~����
�&9�� ���s;0d}��J�n��HM�����n҇k]�[N\�TP��� �\�p� �G͟�bf�Ɍ��N�-���s�C< �@y�o�+@�����2qP;x�	;�aط�KHY�B��F��W
��G x���;-��Xt�Qo�Q�5L�h�z�sV�~
c�n{��+\���$.w��������L2�ԉ2`��a�+����T�K�~�S��Qk����bH������w��S����O����އ3�װ�u%�V��c�|?Y��p������ ���X,�׾����';�[u??qԼ��^4 �r�|�`�	�u?��@���Ԑ�����<WQ
�-m���P��aO �̀�x��f7�Fй�yj�.�b�Y^M���sn�#z�?H��8+e�j�1/ͮ�E�f�0�F�@9Y���u$��m�N
�����d`�ȏDzeMm��_�n�<#��qz�ހJ�z��L��T��d{������2ncG8`�l �R'3�k	��滐غ�1�k2Z�/��	��{��*�fs���������C吝�,�z9��{����c9[��1о��Ȫ�&A�A3Ն�*t������I�䙓B'�|���ԍyp��
��I�AUQ-�!�,��8@�P�]�U[��D	�ă���iƔ���&�NX�v;���c�V9)L��Ӊv���b ]�m����ڕeo�V�ک�A�����꧉:�?�<Y�����k�(�i;�������$:(���͹�8�)�=*�h�C���$2H`=��Z<~�?��DK6���nd�ɭ3#>'�H��Gnh��c> s� ��U�t������	��A5��a�:yS��a�6w�0以�õ ��3�H�$2�^��k�&v�M��['ƌ��B��8m���ѹ50L��qK�in��������x��'�}�pM����y%Jw��w��=m�r-<󣮊E�����_L���Qiz'[�������]�/����ϋ);w�d���6�o�h3n��5��E+S�p[5��#���u�� (�t�B�u��V�����/��.,	��wi�:�r�e;�Ρ�,����N���*��b|�{�j��W0+ax����Wр,G�&H��R����Zn
���&mt�h;!+¹�ɰ��-4)�i?�m��X0�h#��`fċmժp���8ЃG�x�G����m�A���0��X���П�e����[�����Ǔ[Q����>��p;�~��O���)%�h��D"�l�؝�}�����.����n�.Cg��Ґ��� �h�s���fu�����Z��~�fT�"Κ�%h�|.�M�>���8�T�:��:���a�d�E28�s~�A�s^�j��r�#��Cj���>3���>���ǻ��M���Z������;��~���p���@���}Љ�l�0tw����3�!����W>$n!����(|�fkZ�Ռ�1��#���;0��b�����*z�z�L7�F=�^r&&{L���60�֒=�.��$���v�����b�xs�S�;�M�Z!H?�~��(dlN-�'ط�v Ub֜�r	��hH�LfuE6�b�GI�"=�~�o�����7�Frcz _t��ba�B�H�<�{@c�`�����l�'ؐ���^K.�jj"�!���-j+{��:�BS��p#yX��5v
;�D�Wz_r.%��f�YT�ަ�6^�]g��v�G,mm��W��B�wX�1>Z~ B�(t�UGU��X��10��#��ڨ�wѩiYz!���k�/w
��D�N�!tUs�%А�0Mt?�^�Yy����ŵ}��&��Ea3����|.%�,��S���3ڧ5�~�٦{T��ᮥq_w��֘#��ܖ�ز��2b���R�U�RF��K�����.>|)�_d�^),~I���	75�.��Y�	��.�Y����0LW�.;�%�2C����}�`�<����>W�M�у��ب�h :�5E��j����f.<y\�ew��F�����{6X�|����L�j�-�>Pٹ�s]bS��(7ڃ�.�4�ɜ������n~�ƾ.�*��%t4y}�����6�ا�T=$�ڐ~'<���պ?��O�t��ᾌ5�b��%շKՔ*LN#Z���/4��IU�^(Dۋ������L!��3�~)�آ�L��eK��-��(�N����9���jsok���p.��(���U��I�2N�p��u�עOZ�8�d�f�j���0��b2�����z��v��I�VW��V�����sD��D�ψ���H��mT�ty�d�u¿0�Of�)7�ވ䑯�� �Yr�v�r�F0�I)�y�j���.�j�2�*���u9\G8���j��}�gl W��Z,�n/�Rd$���DT�Ӷq�U{|`{��}�ꠃ�&RR���ksq�0@�f}�r�"�/��;nc�4A<nAz0�� �~</����i���.����P�~cS��_� �'O.S$퍼\=PWR�C
��}�
�Z�0�B��.�@f$�WN���Y&�q'���K��"�剥�=8�m�^$�m���j� �N���0��V�_���q���;HI�[��,\=�d*Y� �m�J����mW3���>|~���hl ,'��UUn��o� ��J�?GkU�/�'�V��b������ZH�'��e�}�����ջ̚��z���-:
�YB��1'q��Bh�?�(m�َ�L;J��&�gh���E?oTRa$��@��g�\'�z>�T�����V������S�\�A��e��Î�9�hL�dR!�b`OSidim�4�s�v�\�T�Mp��#:�ώ��;�;YB%&m6S���q��b�?�3OM݌5��:q�6$ߔ��A��wNKEφ~c��J�1��q����,��l"��~�8��_���4-����ZUxƦ��� �d�-�������b+7���ȇ׻#R�����3;2s�\��є�^�7��X�9*���?�7��د齱�胬��5'Rr���l��E$_f�{��?���։@��._��b���^�@���lӄh��6*n[f׈��/驱�5}�gY�;����X<�2�NF2��n�������1f�P{�e�;)���#q� ]�]z��%��X��/�ǲ6z�C�ND���73��/'D���-�!M�zr�Ԥ�4b)Dy�������UX���7���*�:h�G�|�gw�~�Dh��Q��/�M���<9	��˻H:�Z���l�W��)tG�¥�,��P���%ј�]��"����Џf��]y�m	����^4��%}~�a�˟�g'�hN���Zb:!�L~��!���ã�h ��=�	�I���튄�������'�,�^�֙gX������:l6�٢�^��w)�A�10sm�����,ZqV&�h���s���X�]�
���ۂ���G|:V�!Ԯ�Pifl�A����x�)��4w�_��l�',�O����U<�E��Td9��Sn�,5S��m��/���͌�r���6������Ԋ��ZYs1��c��)�7�c���
S�\Z	��y&���T�pե)�D���lOU�'�����%�vrQ�=�"y�!�\��������y �U2$�D1���\Y��r M0�\�, u�Prf)�@�n���(����q'�M�M�
��s��v���F�N5�,��!�`:5�T(���v�4�C�v����~{�c���2�.�a��}1R���T�z��{W���nc�˃�?�}����,xGd�q��^��^�'Hv�!'�m�oN����N�����7ݵ���ugSr�pO$.N�<�cFY|��9�^�n!�j2������Cg�W��h�4��7[ΒC�gNB���[@9���S�� k˦b�KFWw��ޛO�"��j�";��`"8h?�-��nD��wy���4�$�M.�`�GN�~F�@�e/�ϊx@wÆ���[�=��Ż���1��S�b�R���7]�fc4mw�[a̸	|��rI�V(PT�?ͅ޷�ҟ��-��ӓ�$��A�>�����n��c��®��%*z��=U��[I�ή�K�6U�Md�E|��oD�Q\"D:}y-d���X�80.5̓��Mi1�\9i]���-��������Ax�O��Ĭ�Y���4p��Y�}w��4�]M�pkJa6�O�eD���q��Sw;��#Eܲ�Ls��B�8gIG�*������z�����^�(m���H">�L��G0�=�T��~�0��p�Б3��'G��3.�m�.P�����O�j�?UK-ĺOp)�ךȜr�.U��hR?�G�Z�G*ƀ9�����'�K���'?>(�L�:�;����dj;`�(l���&������w�|�h����y��ۜk��)df��3a��>��4Yy�*�~hȰP���d(�H6��Q��i�"��pv"�^�&� �B%�c�������B[ɶj�N\�랏7�����hH��K�����bYYf0Dk�N!e�X�{�rn	S/�U�_;M��'n@�R(!�V�k�S��YVW�6}��f��rjܷ������J���:
E9 �Ș�jV�����Q	���Ɓգ;1��s����Ny$�,`cI����fcˏ�%51]�yL�5��	���>���U��b�-��c�-=+�.��ְ~�����:Ǳɋ:t�~�c�b�fg�ԟwrlD���U���{�~�4o���E�7�N�kY�qPFt�Vk���\�$�t����q�|)B��t�c�Y��ټ2�?S�I�>�%Y�,3�Ab���h�˫�Ssw�����8]��m�;NG%�k�5Y�%���g��X���]m�~�:�H�(:���]����O�mV\{uZ�,�:�:Fy_CV1�>�T��u�CW\3����`GL�	�$e����������t�&��F��JJ�Ob�,f�gt�K],�lw�k �f's<�7e]\�:�����RX�Z�"��:j_c�(#�׌� �0�yS���#�<�������y|ָ�*���`�i�t��VE��b1��P�E�N�-���$�%�1�rH�{��{��(�t���g���y��~ʊ�Q��DG%�h8����E�ݒ�qq�9z���窻!�m���4�{ �rH���TҚw9�*y�����}_K4�XcI^����br��[s��1�F�xbb@�p�4kf��M�>f�,S��<	(2����e��P@ݞ�p#���m�K��~̓����#
�s�Z�^�E���n���2�3���,
���M��J
x�O��s� �[��~p��������i��bv�T;�m��de����y�7���e�/h��h~�)�_�^�\R�ɪ?ZR�� n=:߷N�KEC��X4:�YV�3S��;C
,u���X0z�AW�	,}��[����\�Q�H7��=�w�cEb�3&��r�>����c3��:�!���ثhg�� �G����� }�.�|OJ�a��z�4�#�A����[��b��"�e �@�Rշ1as�&9�u���e��6�|p�s�^DZg����g�=�H���73B*$��<���3]�錬��$�,�����A���O�ks���ؘ@i��cT�`����&��L��0��.�E��*դ|��'�z|�r�ҀR��J��4CH�'��~x�B("���Wͮ�$#�"zD];�^#�Ra�^KΠWF�v9��H>I�rX΄�Ф�|�_�N�3'��g�\5�7�1���ޓ������]F��$>�хP�U]d�W�����9�4z�}�?B�OYn!�L6gJ�G���{"hu��-"_ح1|7�u#��ui���_�U�ꢹ�e�_�݀2x"!�I�o�?=�@����W匒�_Hzu�v�����Sn�ͽ䞉��Y:PV���H��og�8-�`zX2����
��-�����M#�+=�j%h�j�C�Ľo'�xq�?1t��gho;M�d�fe��R[c��^��T��=I+1���yP��c+_�v�����֝l���~��]�����q�h����)OJ}�2:�T��p�3�U�\�F!ϟ?(J$���� �=F�_�@�<+K��4�~�(�H�O�s���z3ZN�����)�I�����`ҦxM��$[���?ƛ2�Z�s���	��\�&:o?�o}S�f=��f�vU�K��s��a�&���*"�.�1p�yPrR*劎S��#֌��.��T{n(�` �ʙ9To3Dvno��WӉ9T-�\�hv���l���:4�pM7Ӕo���"���v����2n
/���r�_b��2��ܛR�TyK)J}�P�-�E�?��9'o!ՄY�q��5�t�g�?���� w=n}�}� Ĺ$z�W��C��i2�C)O����7�!=���U�Ö!o�~���ϻ�љ?�a�)j>N�{ҳc��B�����|3��������`���栛�9����;�h,��2��Z�h[-\>�H>�l�+��@���^���!��ygс�Z��4
���������3�X��(�q?�����?���)���=���5���4 ~W2� ww�#Ț��3<�An�5�1���S���������T��������%���e@|p	]�	���}0�J��\l \@/'ד(R7ٕ_6��G�FC$��}ˁ7)�0���?�ԣ�X�-2]^�ޞ�+-�V��x!r���x]@Av�����%B�|a��a��5���lz��߱��4Z+Os�m�T�ꩿI�za��=�c������:}6�BQ۶�|hi���:A�����}X��^.e_���% Sۤ�3�d0uy3���Z�n��l��Ex3R�}�|P���ټz��1N�f�uf���l ��ج��g�P3�$g���b�^�U؎Y���Ai�]OZ~��8���(��f�D�;"���ۚ:<�w��A�=�?�%�Z6R`������:5��\�p[�&�=޳i"�P�N����ʭ�RO���h&:��R��/�b��WPS��	���xj5���|_�L%���^�3v�V��z�Bi���<!�J=O�命�YB@�G�Q�S��K�Ց�ܽ�㦥%δ���=Չ� ���Y	57�#GZ�穏�g�|�W �r��V�'[䘎(�p�
��� @j|���K�-�N
J)_�]H�c>�o%�MVg43P!��8K9y��g�4��ŋ���ӳu�Q�2韰����)+ ��PY�O�{���(if�pI Z��F��3�W+sx���Gl�ف��e��o��6p��%��k^rm@�+����9�:P�9�A��q󙋂AGd ��fZ��p�vO�/����F�L$D��7sNg|���Q����\��Ok��'l�X3�Y��(΅��N�Z��=)�����`��@:�M�0B��4Z/���|Mٷоw
Py}�9��rMB��{%��poz󒒵֡ �M�
�// g�����o4O��z@�W��0h�!v-FP~� ��=E9:_y)\�*��ScM��Gs��-�-	=��E^���u>TRl��:��A~?��J�������9�k��c��u�]��e�ʬ��F����/PW�dLςP�y���H�6q��\3JVa��M5�x����}�LW�ӱQVo$����H����M�.�c��?���7�E78^^�Ԓ=H��	��9��W���$F���0%u�=���fd�����S-�:������g[,�Xi��WB�u�s"&�����lN�Q�j�q'^?�����ܬOlr���B�� �0�W�E7Z�M��E�pT�ȃRɪ����b4�%���^����~Eߡ���K�w�~F�O���3��Z�Ȇ�=6��/�l;���p�QY`�~.f
��4�(��~Ϊψ�4p�7`,����d�{]s�r��ѫif\�>DE� 6L����)�S�Ƈlk����Y�Or�W���T�J��3�^�����Z��Pkn߫A��>jgLHa/�7
j�#��hǝ3�
�����sS�$aQ�Z�̒�mM���8j!K��J����q>	�Ruc� ئw@v��V��E��7^B�2˜�'e��j�?Um/cpl����<�S������ ��)����f���ND=p�S_٣Ÿ�kJ]|ߠ�u�n�a.�lxy�wG��v��z3�*&������}����6�c�	��Q�x���?�i���r�?:�M���*Ed9W�g����p�(o�4�^x�&�&ǰ��ꌷa�h>.�%ɯ�E��?���_���e0a�[�⡘^����Z�����OFso�0���t��?�#�p��#�+T�����t���*��Ɛ,��t�a4��r����	�>�cS�("X�Xl�o�T��T��g�P^�HBx���3��&WF"���yV<1I�	p\��5���,,B���I�I`;�a�gƠ=_��t�n���X$x�<��WF��!* |]�]��u��a?�p���⹜���&��D���)�<#<G��Ό�L/:B�����1Kl�.s6��Ī���Ɵ���Խ�v���K~_���O�պ ߣ$��^y(U��o#�3�����:�,���h�4s�����F���mwm0�U]@���
}�g�A�خ��5� �V�?��jqb�&`SM��L(,.շ�i�&R�]aV}ƨ�>�	5�A�fҺ��Ͻؕ�0������Kp���n�&���e�+c�e��� ���8�7�r�.��Y�X���Ӵ��5"�v���ȪqNl���:��#��*a\���������0�нcs)�s�in��k5=�k�9�1zF�Y�_��1I�6��m�Qb������40?��A#�萮mf�&���4�����Ӄ�LuY��3�P�m>>�M]w��6P���2b������"&���h�tY�F�_��*��O\|��?î�H��[|�7�{���皂xŦ��h���%�}�N�h��=Yk��$�
��I� ˼jGk;�5u{�a<k|8ް,ٸ��W���L{��-.�V�(E��Kuޘ?�O�߳H��Xܱ8����j�j"XnS�725�xʑ	�7>O�ʹ*r>'�(�1����>���Z���e_�'�?��mw]�¤A�V~�K�m�,�7 ��h������".��l$  5C����N)V�#A�Q�5�VQ�n�C��8[Rkd%>�Ils��!�&ۊ�N���Ag��'�I�Z����J/ۡL�^C�h�� 35��0;#2��NR�� ��4����iiZ��,�:z��X��y���_>D#_=Vr�1�&�?�\+q8zy~f�6�7��*�.U�`�'> ���C�������PP�>h9ݩ�V]!��J@����d���D@�&2^��|X��#>����fVg��z}lC�Y��i{�-C�D��%U#2L�/�>%
�2�ӤC��T���Qw��>6�D �P�R�p���3bQa��4i��*/E��_�;�"1|�o�^B�����-,Sdo��f���L�m���:	�?�v�GD�LXI
��gEִ��aK=� _P����c�G�6�]M6��聞1���O1,@k�
*���v�MWf7�E�`NTw`�N�H����-V���y��G�g�S?�
����#{���95s{���Z���5_/6eh�:s�l�1��p�ԑ�	���0�Q\�@���ig;���DX�:��ln�tq\�e=,�4�<_Z�f��n���2�3���L���-�d�FD���ăx�P��H�z���K��i�4$䴴���U�_��ُ�sI.UK%*D)�Q�]�$_�z2ςf��͚z *���$|�F����͊-�!9p]=�ߣ7�U�c�"3����a B�-ݶ��5�sp�H�|�j`�.��GU%��JK�݀���#J��E��ө+L�f�zr�Zg����\�	pr2��Q'�A�d�?��ut��=ey�G��j�@�b�?P%k����JS#�Z��#*�q���W�z����X�\WC�!�7�"���Yjp1P~�vh�qc-x�G��Q�v��x'�Y;�r��W{�fh#���ύO��(�;�w-�.�׺�m���2�?x���5��kǗ �&��nm����'�j���x%�����PU�t(��;ڮo�\Z��M[�/!1O5ˡ ��{�d�X 9�M�ւP����Q7���+Q�1ǌ��Y&�q@��-ˌ��d��mg��ﻑ���,d�&Gʴ�H� ��.7��E4�� ��[w��W��#|^~����_��[����1�8��@��r:����a���3�����d汤��.#���<���h����U��V�MgJW3S��pU�ANm�ն����D3)��-�e����G�^���e���QOOu��4����Ƙj�Bv��N��w��=̉@:7B�p��4�;�!�����_����v�>�N���m����O�Թ�	��+�v�o�k��:-���g�����OGzϗ��*�9y�����T���>�8K��`��[8˸�s�C~n{�{�rӥ��v�6��M�㟇zĹ�6�0=�yJ8d��s��������[���е'" o��(�� '�nd���2�7�d~��U��8$�D�<��˴�����w��HZ6������z����"|�P$:���aA��Oa�X��SQ����~�!@�2�x��;G������3ָ����ߜ�����\p2��P�����bC���&M�'�|i��##�y2v'&3�����{��]�`�Y~��?�+V����x�CH�e(�pF��VnZ���v�(��4�g#<\�J�-��&u�R�\<�ǲ����S��{�f�)cʵ�=1��k�T<��*�#�Wf�V2 
��ү���}���o�[3������*�H5(�ْ"��$񽢼� �%��*�:G�������V���2/(˖y�r*�:,�U����$M[x�a�g�c�4mM&��[��4��M���p��u��n-3.��	��˷�q,�:�H�vئIu0���e[l��r����|���v/����@H���@ѩ���c������N���
��Y�i)��ˁ"H-+�@y	��W�o>C)���nٛ�oS�4e�s_�uR�%F�kj��(�j73WEc���?������Иo��.�0�������ȸ��+���	����g�e�lg�Mn�����r����l[��/Q��/��i�P�������)�+O����=��9<ƌ_\��Ë�D��q���ۊ����I��e?�>�^�dA���n@Y�)����Xc����rV��u:���\��9��R���Sx������~��;!?��cgmc��÷���E� gt�����kb�?�v+ڴ���s��m��[
+��"�LO��𜽋 e�<\ ���6���qK�γ���u��.��o�Qy[�;I
��~��Kג�a1ji�u0�MW��WAb?�]�;d�1�C��u�:��1��(�G������W	?,�O�\���7;c�,CJCF�}e�stխRT�O�Ks�t��t�_�s�hN�x�Q����=Z��Nf0�lH�j��j�fnQ����^V\��!�(<��u��K�U�e-�{m]��H)Y̳�ڴH��n��xpQ�%��*X��e���r���&NX����JS6$K��L�u��������bA���Xr7�.�c��M�1gĿC�0��6�W2U�:h�ō	�ޑ���a�PZv�iq4�y"@5��L��ѳ Kӯ��2F���[�����(t6�dD�OY��g�r��O������>���Sv��z�� �_��ᶠ�Z��*����\��.Dɱ"�
щ��k����@���i8GF��-��xT=��x#���1@�9c�ك�	B O��(�b���B�i\����"��к�3������}4���4,��Yj�̿<<�#H��54�Ո�* Iv��Qi^#{��%%٩b,�9dSx7�0�aD�������M�M�)����j���?�O���{xp����kD�>U�Τ���FXx5��"w�h��2�C��ɦY�c���e��S��/W*4-C���]u�V��3�Lp�F?�!�������+r����$�(Y �����[aWܘi�ǡ:��/r�΅{��^�C(́x�p"07�`��w����CN�2	�U�mt3gh[NhU�u�a�|�+���5�Jͥ�-B*-,���K�7M��[Bʽ��hġ#���|3�=����.٘[s��Z��f��N��ъt�%/�eͳ��a���XP��:lg���͈S&@�9KW)eAHͭ����,�g��7�*� Cs�Ca���L���X��⋲��UL�]�ܲŊh��<8<y���9��Vi�SB
�62&n<��8L4���j�=��Ǣu���=Ϋ�8In�3�.;I�`Ҹ�0L��tYW�%D����}��I��"kH6�j��-6�ҡ��J`ȹ	��zNz�Y�[w!��;�V��`BD����§��	2����τS��fG���!�1S�s>����x�Zd���h��#�K^b�oFΝ�� J��+��\����xO7'����O�L!���;ā��,�p���vw2���Cx
eMF?�V�q����9cOv���Ujt�p�sS�1�) �P�����^�IfC���❳���yf�Cc9<ϔ��[��d(��\�(���]�������5$�h^~��:hO�]I����cm5C�[��Y�ץ=}r��w6)U��B�[?��f�VI�̩����)�_S)��;�<E���L͓ߴ���J^���6則�h�y��p�����u������1.A��C6�Y��}��JHI�n��/���cw�%�ɽ�I�K^�����z��K���e/�PV"$�}RޘG+��=Q�<��l~'��71�E��_W>
4_x��<���@ΡP �  �U�h%��W�kf_A���&��3��Y5S���	[�3N攄-2k >a1ɮt��8���	t�� �+w��A�_gZ�}��6l�(��Iq]��1�<��~n�<kL�8�Q��2H�Kԩ����{�����R6|?4���-Ed7*��ޜ\��sN��p�3�d}�ZzAz�?��i��ZކaP��Kj����;�z?��6(ħ��R�����p>n!�I&8:B͎[³U�^��`_��Κ�� �h���`i�aF�-L��\��������?���Ks#��74�]�6���
�ʱI�@�i��%����+�n֓>�����]C��j+c���U1��GK)GN%B	�lu�+��5�~�|�4j�������kW{eW��B�_�E��z���Q��"�n�M,�M��pӄ�l�<F��7��`QQ���1*F��
�L����!|kDN�}�ݓ�q��JM�̫��m~xR9���!�!�_i���j��`?�h��5�����'n[Ê"��H"��o�<J�:s�vPg�EB�H�\bn��{Tv���.�.�H�e���n����}�<�J�e�O3!U�|#��}���{3�0C��LT��RXG�'ft%] ~?�9�^O���Ɲ(ƹ�O i�OP��V#k,�H*D��x|�;�Q� J���ڽWDp�&�u�Dv_s��9DM���#jT,�ݏ-��s�i�Y��g���YT�q'�h^(�q �~ʔ��`]��RKN/6�qxI.����%�&�ut#�����ti�йL�b�S��,�8�o� ���n{ M���E�w��y;�>�C-��]�`�"�s���2�$9H��;iV
�$�rp�������P��8+�=[����8��`��b�<G��?�=X��	��Fn��Vf&�T���Z/)�Z�Bؼ�|$�<K�9�H�=�xk��7�L���[�D(~MZ���>"�ւ��~}�nM��YY$9�?آk���z<5�\���R/k0�N��8"wHr�0v*�kf0�69��b�u^[���#��Z��K���i τ}�3q�n$�/!�+2�r�ք'ӏ����UH���l`Jxq/��C ������è8��`�iK�%d�7�,M������:(B���xJ�@&F�5����X`�-�z��5�U7�}��h'*=�8up���t*v�+i���{��x�m#_�[���Ryt �e�Wrw�^��U8���f���S):SR��\�7���A	r��lH���"�&��e~\m��d�"�1B���de�|���v�S�`�?�앏S�s �B/H��` ��*��x<l*oCqOkoX���2&��'Xa����>��՟����|��S�&U���[�*�����j7��8PM��G�$��mXXeq��`e�y˫�5)��6q7�IM]�p����ۈ;c!G��/cW�eL��=����j�>�y��Z�2��Ic_!W�k!�J�"����_��w>8�����БiM��*5.r��rɛs�$��B�+&5��~������#�.�0�����S�s��jֺ��6�u?��*���*�si+��0s�5�V���#<ء�P"����Z�J�d~�)�t8����Ȉ[���2%:�;r~��6�^��S7N��&�㲁}I5@����[�'�B�j�	M<	V�&�c�r���b2mg,��xQ�W%��/sHZ��� �򳶨�[�}Q伄�f��¢�mS�a����I}̽�&uڅ�ꠚ��[�D!���#S�(�����������J3����O�!����g��ӷਓ�
0:�^��� ���]R�J$�8.��Ҋ^(�c��)��$��߸�y�{+��iOqR��5��D���!C�1��%F���@�ވ6T��Cn?�ht;Y�k1pτ7x����x�t�C�$��`����M��&��!���6
<���b6|�%X�#�gk��|"9����'���FUq�����P��ЀDeY���8"�M��!���_ŏݜ%��Ե�<�w�j0��\٩�}��xW����(CEO5�c��0t�#��z�Ok|�*��K?,���]�7�g�ѝ�_��Z"��`қy_;�@���U��淵�e�mx��i�
*(W�$��
����~Y��9��Oۿ/<Q��E��S��R�0�N�W���?_
t�pcjuOWS+Xx��\�f�]��m�}��2�Fe����;��kN&tJ΍��u����n�Xٖ{��o�lo�1��d�]���'dG����
ӦVN�>Ń��QpGIS�
����@�ut\�3�Hxs��ߓ
��By{�s-��)�	��)�7NAD �?��EA�f��O��㦆�Z��{A?��ܜ~�N4m�q�Q95��<�*f�Z�x��{z#�J��@/��`IV-��#F%L�a(��Rqٳ�C�R5�~^6MM#�[��I[�1i��:żr����%xc��֣7x�a����]�_���E*�qgV7�#x�����!��a5��m��r�r�Vp�ˆ2�ːBD� -Z}R���ZV��4��9���Ā�qm�V��J�o���GR�A����}��NLèAۨ�4x<��QaG�B���)U�'-��)�_P�8�q�M0��/�;F�5E����>��HgU�����ɺ/c���LO�1�֋d�=��b��Gy�5c���.B���րCsW�k�2+��Fp�3<wj�_�w��KX��~��J4�&ղ�ś^��n:%9��_�|��`��/�iѮK�-TaZ���Z�F�IP6X��5�k��2�(�0����ҭ,����ǺT+n��{���ڣ^��
.�V���Y
�.3b�m&�ct(ϛVϘ��]n���H��Z�FfS[µ����L'���Vs�МC7�kنĤ/5�
��X-�cҮ| �Du�FM�=��|���$G�A�kS.E;��H@i��b�����W�ZĭxA�8'�F�+TVq��lϬF�RVǘ��?��;f�h/_�|J,�F)5jK���;����+(�a��nkS3lgR�p8�V.��I�,�:븼�}���n�C*+_i�f0����ڊC�L�Jeb�����1��	���%bYTmj��%��Q�����5�mW^���_�ET&L�u��>���
?+U.�%3WSGH���1��Y쵣3��QӺ5_SS�%ٴ�o���S��!�5��z����7��&6��]�=9�CK�f�G���w�&9J0~�����y�&��ȭvXL^�\�,w���zJ�;�u��s�Vw�&�U���aJS���>9����S͖g��^��uC4	y�0�����v�y�z�9GR�baY�������1�H����֢F�U ��$��r _�^ ���:1��]Z�^:'�?c�����xHG��U�WGW��M��Ѕ�7P��1��UP9�'�����x.�֨�Q��V$�m[1���z�Dׁ��lٯ+Ϋyj��fz>�Tr�/AJ-�b�:�]w�1�lEZM^�F��s��Boc�# �q ��74@=��.t����p!��S��SA��_�� m�A~>�E�+���U�p�Ɏvc-( �G�B�]��=nB��U���X9�%,��E��5��,#���u��|�g���h=OR�9�UN@���QC��ϋ{�ۇ�$G.,�4eg{�
WḒ�(+*��`� �ˍ�uK�(�+�	�ʔ�� ,�!�8SɅ�<��RT��Y%�ZAU�$��UN'LAS��R�P9WMZ��ϰ˂m����0؅��b� lr�$�H |���-�-/��g}�5K��/�{C��*�q\���u�de��sNޱI��heu��Q;�������ʹ��F�C��O�M2�`�S'i�ڨ���J�qS�24+��,-��_Y��q�"f�=�y퍀�����U�X���Ͱ̢y�6����_��m��B�x~�6��:�] � �Qa �H`�*Ҟ·�4Ӥ \C1��\R��������2�������˱�c�JРޛ��.��^u*�˱n,d@��q$��sXbǈm�������g��
!LD��x��s�S�F1��b4*�P=P��R�W��50��ꠟN,�����8� ��=r�D�z�ґ�>����O�R���ZBT��t/����l�}��5�*,�����L�TZ�6f'��KÐ?���}T��]�������C����Fjx��Q*|AOM����mt�`�1��A����N�o����S��3�VZv�����F�{�:��k^J�̖�g��(�[�EZWT��N>+�C���V#?�9`J�Y�M�o�H�>�BiMR�`��k���������,�bv�'
��3���5Q����sp��D�����PF[g(d��k��(�8R��a�qaݫն:��ݶXT�����@�	��a�+\1u�;�=5R_g����4�o�I�|(��^� �!�;ù���ux��y_z��#Å��g`�������-��/�W\P[)1lؤ�)`l@2�D�
_h�T
���v�wWh�~��a�B����i��h �Ơ��]� �G�~�ʙ�A,��%iz���#��_���I��=ٳ��'I-��Q������'z�����1as��Ъ��&�����e�̔H2R�XQ���8��Jf�~���-��7���J��Q�{�dy~�c ݦg�% ���5KH��T�֔�MUN'��ǜ~� O̐ޟ��{%--��u ��<엒y��,y�����ޔ����V�䎽⬉|�f,GC��_���R�4�«x�&�Xk�����4V����b*��j��Wvv4���\�do ��2|��?�z�g��	��^l�)&�qfj,�
��m)�q.mw�Vis��������MQ���g�fu.F�9�R�o*O��b�z$srwD�2�ܙ�h��Kޗ��xY��VN� ���M�=���3�"*���PYdg�����whF������i����hZY�3�&b������wk���Y��+"�EME�:���v �
S�x ���D5씅 �-q�{)��$�:�E��:���@�����Ҍr� ��q����2�3 h�s��|`�cl��mm|;{� USUl�K�������f�������OdsĽ���0�[���zEۯT2n+��N�%E�ZU�둻֊쮞���Ǖ�5�����N�h���C��B;:�p��!���u��$5�[�͜6�F�N���%�& �<	!���CSV�����,D��m�J��K2���6�Vf�G�3��l�x�fz���Z�F�4۔u�7#mx���:]j�<�R߶,�țwc�e�.�Qqҳ�v6�z��O�x���Ʈ�P6o���Y���?"d=Ȗ�r6��"��F6�Y=SJ)���ZT���1�*ܤn���N[:�LYI���Fܪ���l�y̪EM�����lya��v����!4ܳ}­���2A��+E��t�{���8�e����H�����?+;Lq@��ڱ^ߜ��A�K����#t��ITe�`k����{jB�>`��P,��5`���@{8�L&Z�V/w�.$�� ��wm-���ݥ��>0�2&V���&�t�uz?�V���[/LO��Q~[n���W�.��C�Xs+��oj{�ݰE��F��G���u���Z�P^����o�cͧ��Ԃ�.Ɣ_=r�t�Y�"�V8u@�/���M�T����F�BFX)"��D4U����m��*�8�<]��%H<;�`ސW9'�4���9Y�P�?��;Y7̇�@��k�I��ߐ�����?�#�o(MټS���5*j����� ��9��i�0u�ω�t 4��r����s=�r��+͗�����i		�y����H��
Feni���$@ ����Hw��!�"~f�cL����R�N	�
W�i�� R��^$� ������<�vu߄���B)����u�����[ϯ��Q�I�ɯ���D#z���tm��MY���A���2������?����5Gb�4����5Z���q�7�ǟR�w��Bޤ}(+��O�N*pT#Xr.3����ھmt�C8���l��*~�n)������o#՛�V�7���y����/�����-,Q�4��9�@�TҳAY��Z6$�������I�^���soo�#��0c2g݌T=��5��{n�d)�������ĶI�Hs�@� ����0꦳ts>E���$@A��{�@ڧB��D�{���ay�/Ό�t4�5�zԝ3N������*�׈l3L+�58�k� �k3�}<�H���xp�-~Z����*Ե����Sc�*�$��e�@u�n`�s�}� ���-4�3d6����ރ[��0Y�By�T��>�:V#?.�
�O��	�RK
냼!u{�� _����5��ݓ�n�%X�x����!�K�u�z.Ua.̀,��
����!�b�.�V��Wc/�z���N��	��o�B�O�h]�q�
�$�N������#��^k�D�lw��4vw_�JH������Vʔ��}�`�WϚ��9�E^�~�G�-�!�K��ߘ1�6:�t��s��2X�&��>BSؐU]m��cp����@@�SZ֌.�B�
�����^��C�3��r�J���Hn�T G�KϷ�
y�VV"��~H�0��H�?/�Ӆ7:�3* 2~�ע�����М{пL�
��ŢBɰ?�(�G���#��q����^���/D�K
i�>4�A ��N��Q)��n�b�o��򯎞HL^�X��z;�&q��qL�L_Nf�.���!����'|���LhP��!��/�;	���R�A�DU
,]hnm���	<v��]�/�^U��\�<:B:��L�-�Q��H��E}�B��F�;�#�;�?E��	�X��Y�a9&y���׆��fd�zqR�ك�+^���ף�hY���w�;��x�����-�R��ӫ��3��99[g�oM��S�t�	�tH�&���B��BiNrvm(�)���-�A�;h��k2�`|�{�U����B+h�+�'�sE
�w�w� %�&��#o���Y���6�1��d�����ʹ1���n �x>��Z����b�>�VL��!�z��]��~��G[�����Q��;3�%~�0���}��1/�ݏM�����v�E�i�L����K@gA��Y`���<5-ʸDCT�&���Ad�@�$-����[y�B����>#@Ƿ�!^E�b���}V��CE�A��+�)AT����p��@b['�ߤ��SxS�8�����X7�_1����/�M>ˏ%��P��_�V�x�`�z�CD|����3�,���0��:��P�;N����1.sг�j?T���5�����u/i~G�O��	Ԑa�عI.�!��v�J?ei0Q=���i�]f�၈H��*/3-�f���Rh�}V�o�Y��AEw4Y9Q��YvXl��;�t���ݢX��◳�ն�o�L<���j�/	����q㕆�.ǥ���%K��r�J��~�����t�f3�wMPh��n�>�z��SAq�C��Z{�`�L��p�����m�F��t�w���
�^����|7���Jf����Z��D�ϓe��͡��ޟC��!��~����������R�XO ��fXD7~�����$���
o��@J�u�Da��Y�P��  ֬t�E�n,�F�W��h���GD����?"lNB����=�w�����o��"�wkoh�����5��|0G�2��-���ܕO���ec4&>}�s��w�| �N12�<�D�؞�NI:���;P�ѥ���~��г��V��Ũa0�I�x�֑Ñ��O0�Q�`��
Rզ�O|�#��v,T����Cyg����'JmT�*��o	�3���P�m4F
�$�)	�]�B��A}0�T+!6�I�'?�)���e�Niv��az�$\��L���l �xJ�m�K��k^)4�zL��g��Pvqy3O��n#�[2*�&|��k�R!���{��u8:�r<;���,��Y}:���YZ"�U7잕���D�\��p� �<s��#��eS����m��پ�,����dM�Ӟ�RW7;!��X��Q�������I��]O#H:������=�L�[gE�(���T���1�f���:x���f*��&��V��V��D�q����O'/�!��,2�*ތ�}
ǯ�P��0��=��n�l3%�P��C<��#i봣G��R�h�+�9%&�M.���}��֧���Q��7D����E}pI��`��#o�Cy��LP�գU[H`>�i@k#�~]�{��HY��?u�%�DٶU��#�Y��峴�ľ�unC�\W�娺�u�Qh�nT�k��Y��r<`D@������k��B���I�(��X$Fl����U� .?�Sx�o>W秂���y��{I*3�*f��]�봍s���k�(�gxSCQ}�< \=��|�s�2����V����4ۜ#z�+_㻬�"#����d/B���)�݃���l��a�L_<�d�#_�j�;�	na`pXU�Cb��#�y���b�8���[�����Y-�.��4�Ū!���8xH�-GW'�4��wbA�Q�j���'����ߖ��[�u���g�^L�#_������yg&��H��3�*�Jog�o���u?�P�YW
�Rs�:@�)�&��0sSƞ-SSw$$��GP��CÜ�TLA����	�HC�{F���ZKB��^y
I�����6�T���U/'$ ��^~����dߨ�~�c��8k�A����P���o�۱
d5��!�����ƭ`tw�3�L.�$�t���z�"u�K)ɼ��nl�k̢����aj��uϨ�[Dc��{P�h�D�l��FX�LL�[{�C2w���ͦ���nt��qρe��S��b�I����lI>JGs,i��=�^�gz��F�����d
���l���~�A�u�{U2
���GZ��?�d�{Ȱ��i����2H�2��H��s��м$N��HAN���"#�����`_<!K@]�Ǣ��
p���0�\s>�(�2�{
��(=��~&��p��t,�%�OD�9-?#�����<լ�pm� h��f ��Y��9�M�c���Jl��zN��5d��x(�? �Q޵�UO�Mş��>�k2�(Bk:��-��#�C*^�l8�
�ʅe��0H��5��@��޸�]�Ξ���<ċ$��|'�niy;�z-c�1��p���\�]p`�M�u[i�IR�a��<j��	�QO���A���P�G���v��Ya_v?1΍M3�ݯk�IH�7-��E��(�^'��%���m���R����v2�f�h��kpK{�coU1��j�k8��@w[S
iUrg�)K׾),��<_Q��͙M5�:h߽4;ե/�C�@�Ԟ�����Ȭ��5�J?n����S��a�}���,�%I���>�ͦTRw �(�Z�A�)H7w���I��}HN�s#�s��_2!��h����ҿ]���h$.��_Dꊗ'D��4�3�c{�*Ck�RKL�R�\�7C)a�W��N`~�4����Q�?Х˿�̀�#!2��r�����ٌD[����_��VT��	~F�g��7�n=�(�hX-U@����,DWz�#G'�q��G���0O@���\�ćT�1�hP��C���,+���~}�~cI}���FT�;	3�M��K<N��ǄnQ��C�-n;���˞N��� �r���7.�Q~M��5%(��֦.+[<�}o(&L�������y�W`?�ׇ�q~�(�%g~N�Xڌ�.��ټ(��	"���@�@���kg�T�_�,'S�F���Xc��	$�+IN��) L�k�o��cP{@�=��@!<wΡ����w��<����a<�M��0����C>�����7��g�׍�4?�� �02�c�L��NH�e�����W��j~/W��<C�r�/X;G-</!����^�[�����������ͣJc{��w��ٹj�N��N���S5�1�7���P
����@��GM�J���m�2h(���V�鋏�4F��ab<+%L�����=��6H�7
7�wo !�����H����;�e�7Spb�?��)|L�يp;���i>"&sR`�~P��A�ؔA3�l��8�i.���Ŀ�M��Gz:�	�'s��;C��h���A�X�MƓ/J⥓�����	����+?}�Z�F�����P��s�D{j�չdR��C����������묁j����Zc�$m�g�B�o�%V�6�nl�r�gXZ��!��I=�Y������8mܘ|Q��\�IY��DH��>�B4d��Lt���-53�DlE
��Y����*jl��:s�T7C?-��<jn6dYHu��p�^9r�m'ϗ�_�0�D_�]^����8�&�8�Ţ���4�*� mPW�4�?��H�p���o��(�
vE�A�Ϥq8�pKXބܜ`+������Gp�9�D.vh��$��^�OT�g67���n咆V�|�{C�����׹e]2$�O]�����N��0i�Y����]�kueSř���P�:.�S��Gb�o����i[%^!�f����4bIyo�R�j�)�����{�߆3��\h��^�$P�Bc��T�A�Ꝣ<���ʈ#���&yc�m��-lvxE�K�	��Bo��l[����T�U�/��,��h�e�w�T)�5��~[Ӽ��"拓�����Q���ڼ�|�"B���bB���L�K������i%���;h�6]p��c��9P� �?~����:�!=�{َ �X��-��>0/`���&��W�R�ҮphH���b
`�:ڬ��rq)gL|a>_Jڳ3�o	���k��$���<<K�u�?GT��'Q�
z��X�J�T/ ���@�d�<$x{l>���/�\�k��,��5�$�>������T����"/�<6hv�9�!Z�=�V��5Ȕ���I>A�^�~������f��I�������k^�-��c�[3�;�h�"o's*p��`4?(��"�������P���?��5S�=*��wPk�0gt�}�{�F���v!���s���-D	�"������v���)�h��h`-��Nu�����W2����<�kP_^X����{9��������������5�uf+�TcWiV�70K8c<�~5~�/�Ꚍ������M�+}�A�<��m��q��«��- /m�ݲjoj*���V��y^9aJ��:�fv�i1O��o(����n;��pv��i(:�`A�����C$\��4<L3�S%&J�A����LY?�4sIs���8�s��b�X��{V��A#���ҙ�i'�xl�j���W�c'66�se���.�G����Nڞ�uL*� ��|EJhz�5�]Q��EF\�	_���o����a�.�ob�����ik�x�r:.ܶ}H���-,{��S��A5;(�b�PD��3������"X��5��D�}����*��'7�����(�H�(�k���Y�*�>�mB^�A��������u������ƍ���*?ј�[*�&f�IdBzZ@���ϒҬ��7-��=� ��^'e�::F�vA@֮�Q���"��dH»�䆕�(�2�|�����3�\��{h���ٳ~5�-2ʗ�;ݎחm��H�R|R��B�QS~סúKT�i=��� �+<���&�MLCћ0�ye�ۜ?(Wp��#�.�0L��#@
��ؔv��p�<�}�1�������x���������GɒO���ǾP%�ś1�[[;���4����X�E")+���i}��
A�C)J�n������T��y�7��[������>������r�W�i�Q�\����|�Oe�w�r���͞��1�8�;A��=x����08� )�/���0G�ڲ��������j�c��8]x��z|��yt�?d;&q7��x��{XowPuZج�0� � &%�'���N���j�R����43�?�&����x�QO,Fw����k&�󄤇�V�=�2No�����9t[1x�z|��z4Sd�Pp�w7�B���0v����H��;�{�id�ɑ�/1����;�e,��,��T&��7�I�XvTt#��j�����~$����=f#��w
W;r������4r���(\ν�*|� #�-�]M�Jg���5�U�)��׉_�Jm�	BZ��I�q1s����w�La�0��+>Nz�� xf�c�B�#�&��=�u�t��������)onլ�ۣi�P��7�rd%��&��/!k�5S��7�%A�T[:���~A�\�܊�ի��@2�z����E�k��Ú�7t�}���ᰚ�Ƣ��y�!���r����΄��^����C�	Ị@f$���F�3޵+�)���g�^�d=�x����|�֬�#�O\�� "^�`(�;�o~�<��C��r2�qZ�Z�3¡�����N�p���;!��"�m��Q"�Ts�0�����o{3_��H;�e��p�T)%��LBc�g�}��
x���G��l0ǲ����F����d�ہN���	M���&L�?I�*��;�m3Nt-�.�UF���j�F�y��"+T ��{a\�������ɲ̷�ٯ���l��j�����@n��m�	����Y�P�y��ZI�Pf��Զ���x�+�5:�Ϝ(a�Z5�j�|��n��$2�3����b�@�bj�L��1����}�J"*!4��u7�E=B�+�,�|u��ƶ��g�0&��G���P:�Շׄ~�ݠE��9��o߶)Ⱥ��&$�Z�����_�Y��_<��x�r��QW}Ǧ.5�70��$��@���mM��ed�u�؋�,���nu��>�D�hTM
a-��Y���u$�s�$�ڦ�ّ'd��:�?ܲA5F?��8�	=wI� QZ�?�f?���RZ4tc
|	����j���(��}MNS+��n��ρ
U[�瓱�����S�Tu���%�'�e�tT�����m�󸽴����Rl�w�$��xm�.*�،�Xf�J�*5W�d�v���� �i�\���� 7��B�m�|՟c| � ���l�={�f�6��BD^Ô�c>u�Ok��, g�d��r��OR��4���(��75��ІԺ�i�~o!y��J�5��{*+�Uo�_�7���|k�������k�H�������"c'���l �Q�q	U_t�#Y��i�n*��XǖI����n��_��֎T�F�J�2� ���h���?e��)zD�Xn��3����W�2�n�Ea��?�_����1���ܱ��V4A��-E��0R�dpz]�~(�Q��ᦞ�C�-
�u��؝��Դ��w#�{�ţ��������2dFl�6�DIG��Lkz�U�>y�����N����
t��a��Rt�L��N�g<�3��fJ�5ᅚYc�@׺nHHM������WT9�b�¸�)�hV���0.�e��#TG����oW�`8{���V	���4D�_P�*D>��捻`��r�)�(�a%5�e���!x����J�A~P4��X�߾��ϑmh�  �'*_�B>(S�R��-�C���b�/[8�"����z<��������lݱ=����z�d�wQD��A���$�R�X��X}xkWb����8���U��P	��G¦�rd��Ru�j��T-�?��FM��Ǳ;\E��l���ͬ=�3�����?�g�{�Wh��`~m��ق!K���y�/,&���U�Wc�on0��w�]ސҟmN�,��vf�zCV��v���Q��RD�(��$ĺ�Ҷ^x	�&ytw����/`Մ�yK�Q�H�Шx���Ph�M��T|�|եG�M^*��Cs���3_��M������Щ�{�#*9)E��S=)؜����ە������.�M3���#�lɛ{�NLo]��2O���OJ�S5O��ce�mZ1���z\	O����a��m�m���oY?0L9u�f3~���U�TZn=үy/�tZ�_�{�j��V�+�G�>��[�|�Rٹ�{�$�[���qf�b�y���â�	GH�O*4hqbrk��f�3�ޱ��u�:!G߈]��CFB6O��^��D�E�KW?ih4���Sңls�t��AU;=^,�og�}�=������S�YL2z�1H9>ɺ�D#����D��0#�%�(`�N���1w�����g&�'�x+Q�fH�D���A5�R���n�(�N�x�-��Gv���l�9Xo����ب�n�i�ka���߳3���l�~3�3O�	�:�0v�g*�6.�VeVO�x�T�]3E���]�O��%$kرQ�֢�ԙ�"������� ��y�0���I���O��GT����%w�Z�t�ь��,cg���a����C�Q{�e6��=�U>�FMRw(�Ԑ�����s����b���VM��#�SP"��sso��$�!6�7�<���SO���Ef��,��� �}��8�J
��A��'�ҙ�Ԥ��M��L�r�A��Vʘ7{��zeEqE��;�5��k�ô��.9J�JA g�����TPO�2��2�&́�^� ��^7G�EZo��k�r����{�4�#-��v)=���񸼻�"؃m�3��̷;�<@֑�q���ɨ��2Y U��U���01�zKÓ��+�_�~��羁5���'� ���7�� ��4�,]o]�{;�?s|�����n���h8+!�����Ʉ�SP����r�WPX�w��q�+�d�P�D��+��f8ߟ�����ϡ�*3�FWӊ��2�F- �7� �&��b�A��D��e��:&g����+�u�+7/O
�'�3ܥ���Y�ƔR����^Ϸ�K9�R4\f����N�F����v�#^p����D*�
mF��l�"�aځ�T�\���nM@�;��{����rf�Ut���Bi�}$��8����dp��N�_���)��\IՁ�C0)���Ȱ=�5�c'��/����<��}�+o��+�eH�<��oQ���@\��.�Nݧ�����8�w~�{��ķ�#�Lʨ�h>F�K�[(�F�H͡��(����_W`X-Zf*�||u;L �!�F�i4ԡ��K�nb��=b,	���!~gJ�x>f�����z�3-�(Ftʫ�~���ݽ2�T��,��E�ż@�f�'������PgX�G@���4p�%��W�~e��c�\r�c�.�_@�;�a�����H��
����t(�JY?�h�B����x>��+�o�g������^���XL��)}s(�a�����|!R
M�b�w�,�)�i�gΦC�7'J�i��^=E��U��yhnD&e�	�>�ȝ��
*�p������|a��@*n���
֬$|8��fx�~Kz[���3G;N$[�N`�ޗ.���a[�n�dE��AL>DV(oK�V��)9�~{(|w�t�j�+��<͔j���{��lºp��2��@-��/��(]҉Ȣ��6�_��3��G�x8�w,$��r߉BvؽU�i	\�T?���l5
PM>ɛ�솑�X�,�JP��ch��q5�g-���L����+Oc��Əv���u����Ol�ng��t�zC�C����*���tJ�!ޝ:��sF���m���W}(�Xo�T���6��|����k1G�{�099~�6c^L��#GԽo��@V�Ȓʛ]��(�e7h�:��~�`��{��IـE�5>�c�.�E2=o��L	q��:I?�8q��G;���E˳�m��Z0����C�χ.P�>� �0&g?���!M5]�@W�M3Ei9m�$3��V�r�*��B���VE�y�^b�YLr.؜ �rC7ǒ�n��8�?ʋ���� R�S�!>3#ͦ/N�b$�3��*���8��T�n�Ic�����$sw��2�9�=7���H�H��UX�[�KA�"{A�=d_��]�����5�q��n.YݧDT����˦��}�f�-��Z�«��a��1gS�D@d��h��;i��u�J�<njB<PK�9a� �D=K��TɃ�g��4<._T�xr��n�"����œ��ye�X���^�\�w �_��C���{1 ����aNN6@V��#:]���i��M���`�M@ְ�'��_�C�Ls<Y�����n��5��	� �:�
J��M�S�l ���I�hD�%���S�=��!�a��]���g����{���O	]a|�,;�_2���DYR�J���i���0�썵-�E6�ۗ�]��$Q�f�����vC)~���i���٧Q�*_�n�q߸��h��#��"#��)&z���b���ܧ5���y[��	�JU���j cY.��u���@���=�(�%U��9�$��j���aT�M��v|�Rq�.F�9�}B�x$Bڕ^�K��٧�yס�	�>���.�۲�m����`R��ä�{J�Z:rJ>Nw����)�!����7a��L����j�k�S� }n�^�us��gM�$��}aL�]YI�Il�Ћ6t�������*2��׹����j(�b��<�'����f9�9�Q�����y�߭Z!��ff�� j1���&cO� �5����'�=Z:*9��:2nc��G �/����4͖"�88#m^����ᙈZ�Pg
H��).�L���
CP'�;k���F��kݟ���^���Զ�y4�&Ҳ%���U2�tj�1�ݿ����Sے~?yC�����T�V���_)5��4�y��1
���\h���KPp�i )�<�ug�
>o{?�L)�1�~�9�*� .�J�w�*��bک�T�6�TҰ�j�S��US.>�Y	Fq�@={����-70I�0���D��u��<����H�7e�+X§����x<�����/��Ѻ�\�AS"[z��0���c�eWq�cgU�W��2�L��׀�&�F?������V��qg�
�B�q���[�*c��u���S!h[���
M�O��]P:I�.q4�v�x�u}s��r���_�LX��)g>y�܁O�'l��D�Ϸ����9B����YZ
��s!y4t�G#Vƽ�$UjGt�7�.�-�QƘH� `jUaA�;���ˆ: �÷����t��{�j��Ό�7=�t�}�&&wP<n�c㷚1hq�]�g�X��$��s�2�S� ��O@�Q�����@�v��굜���{�+��vМ�
 ��uN�7�sH�����R6��S%C8�hE�z�1x�6�dr%�"���M��d����f/r�,(���Zk/ֺ�^f�b蟎���X�Z�bW"���	�i $m��73$�m#��{��v�}:�w#i��cV#iG�n]����a�e<��ן���x���@��QH�_}���_$�$����㤏^e��n�|к��(_��"3ob���9'��_����!�~K]5�y.ߦÙ�u17��!����	��6�z��<E��'�[�2d����׿dَ}�ڝ)#��Gg�ޓ��8X�ٓK:�~��;�����$�rv�y.I.�T�S�<���u�r� 6hn�	)�U��p�_Z;�4�=�]P/�O4k퉗��|��e���c;�ؠ��;#�Yeʯ^���dߚWHp_$�nYzE�2I\�ĭI4n���+�s`��Gʬ;�5��9����%9��_�EK�F�fCV�v�8�^��6�R�����������:��ahc�,�LZ�SѦ
6^+z��r�K�����.z��/�Z٥�C�Hx��ɠ#M��H/R�O+(E��'�4P/��������f��ɨnc�&�g���X��R"���I �S7�ٺ4�.����h�7��]�yJ6��+�9{䄭7�J�7S��� >	��͆FY"8�O'_l�"'k�j&�9��lr�l�fx����+ܭgTY�/���|��8��a*����v�rAL��c�� ̮&���i堰�..��֛ ����\���d��Н	�����VY�5;+S+���pU��|���)j�I�!�_-ͬ���AR;'(�J�#h?���}�E�h0 R7�W�(�#�������=:�5�^��T4��mo�n;��茺m8�^\.���(��;򍒬L����tW	�y��"3m^xx���%��zq��#��	B]ksγ�;� ��ut�S�:�l����H�N�$u���g�R�T�m�i����=�=x#��m�[����"]�g��4����@�'�
��K��m#'��Ǻ��;���((�A��~��Ì�S�)���k	�G��Θ}{���( ��;&ճ֒ir���Iڂ�f�M��K�oa=7w^!��v^*�!S)A,3i�H+�(�ŝgz���^���<�OG+���?�:�T����r�$iq&�vY��!��$?��A�@,M��������}89vȋ.��6��iҪ��MV�Íjzԁz^av$lv1�ۢc���A��\�ȍ��z�Td�w��b��:�f�E��!�(Z+���R����
Q��_��Vy�F�О�*��+Jɽ�Gt׬@��X��g�]1 j��R"~d1���n�O�m*����z`��U�5�as��-n4_�Wy����.ZN��n��_�8Z8$�6��6��/}�0�����z�cߐL�{)	�&��`�**E�䕰�u��E��"+��2	^�����,��<�m���mLw�z\J=�'V��=?"4B]�ncި����E��_'��`�v���𗷫+���wZ���݆����B3�IzN))�)���P��\=@h�w���G�N�?<C�q���GO��U�3�a+o0~+��?{f~�bS�=�H�$~E���D�NF:����S��-��(��W�U �>�����_S)�\�vnݣ��=�k�w�|�H!�KY.��i�풠�g����<x89�p�� 1��qK���s=��o׭w���=z��f�϶Aٗ�^g��X�N��X�c������_ZFs����>����`��/Cd�?��Y��CVj���@,b^��+�z;���0rI���$��4_Fy<Y���=��TO�X�2���7��p��qST�;2g��7���Ϻ^a��T�*��Ǣ���l̬S���ظ�I�(yK
_�P3���ƚWߜ(Iݑ���*w�Uo�f
�R������u����O~mHj:�?��~���ؿ@"{��Vl(�K�<���@^�?;�E��b�Z"�{���� �(i%�`�����&^~C�}(����| �N7���9s�	*�϶��a�@�Y� �^U�ԗ�I�H�Q�ˌ��r!�q%�	*���!��@��W�)*:���G��v���&6��6ωf��7O�H;	�n�SS�,�t�4Bd=>B�s��E�`zק��e3�<g�:����'T7;Ԛ6�h����S��I�5���	��Zt�_O�h���%��|�V�ңQV��P���ov��נ�n�M1�E�2\L���d;3�3]5��q�V_��޺Y��W��r�v��a��ns~ʕ��}���N�dF�e�1w�-_Sn�T�"$��_S��g���R&�`�m��U5N�A����2�)T��X-�؜*��ђl��l��L/���;?L�+%LP�I�_�n<��N�H���xш�%<j�zY�[�ܘ:�w޼�?:�]Nw5��K�Y����QG�X��B�Q}L��H�j�Q�0<�]�U�n�1�MD�R�/Ko���X��7k(�櫓��S�/?c/jş�D,(��˖TzG�=����a�������c����|	7VW-�l[�̓�T+O�DR�����j?��^-�qO��x�b��� "ӹO��$�rG���t^ֵqc�P��2�M��lT����j(���0ޭ*WFf��{��3��.7~�G�vA^�94P���]���9��HԊ�ub|����Ƣ��[f�E�2��@w���ragd5��~��n�?!V���A�$(jl�Д9��g�_<�d�"�L��.�A�hL#���iSP�&��a3��ܓB��A�^��0��ͯ��?�;|��$�������v��$�эQ
�\�2��_��{�v6�B�T!XWL��� -y�a7pS5'S�_go���>޲��ʱ��*��FA<HP���Y�x��O8ѓ#����p�g����^߫�Ux�}ե�\Q����:K�W[�x������~v ��(텏�^�e~�^E��B���<�)��xsmlC��J���M�L��*�f�sx�޸\����]�"���+��A(�եm��K^����"y�$��B�/�z��4�\��<�a\Ywl�֫܃J,�E��quk�M�H��6s��m;ff��H(�X�����ҕ���n"Fw�ʉ1}�uYew��6�����Q�&.��8�?�>��1�^���Sg�Ս����>���9� X6}u��$s��;Y���$nso�|���03�Q'Mc69^�7��u\����
���7$r���-�Ϟ�
��(�id@i�P#tC�9���)V����0/��a�c��MC[p�� �O�̯b�L��,�d���?r��x��`/�T``�����Vr�VF�����eitE��f�`/�I��)�y�D
C��Hz�av8r�S����$IOF�V֕�3��O���^���4)���ϙ"�ݎ���uǊ�S�AF �/�Z���b���Rm���o��&�Aڗ|��s�~F0�oc��S��:��P3F~�����C̚�k,L�$�噊���g�2���w Z[Q����r�����g�-��Epx��������Q�,���qVSS*�B&��*IbQ�Z������fA�yL2�$�X
���Z����z���ޚ@x�7Z� ־QU��y��r*�jL��,)	�L�?cUwIIE�PR�U��#���vvx!��&"&:Y%!>�F��S�OΜ� "@�S����d�~û툎n�0��!�-�)Y�?P�]d>�/;��d��5g��,8��y�ʆ�C|���I��?a��Ƥ(
J���2A�OI��A�_�*QiHOo/�-��ڊZ����(�1����<�'e{�DII0R�7��ȏg-zm�P�ǝ�=%�inb���}�*z<�lL4w&4SBj�RR"��*}��K��bQp�/�b⸵������}����3�1^񫑇}Gs3���f­�vW���Ǟ�?��ܮ���*�բ�$9~��<w��1�
��O�n��T���)�cC�9Y����ZV��=AA��^H�OJ����lv
	&y�r�����c4�TB�m��sDc/"�̐s���a��A�Y؁54�@b�x6�E[�̑�l�(��q|�K�.�{;�2�	�Y�V�Z�UR�j�Z1[��W��\�R�ʟv�~߆Q�u����<b���$9�P�u�g14+��r�9D��4�ʊ�Q:�!jE[u�2�U���
����Zt�;�ֿu���0�.�W7�԰2���`W�em�d�CKϸԟ��A�� ].߀R=� �=�׼����S<��'���;N]�(�1�Wr(�ٌ����p�[j���wW���N���>�`��s|=1�S�R��u�g�#1yht}��zB�x.f�g�PVocBr��x|�/�)�gT"�u���9H��d�ڰ[x2#�E5�+k�k��k�8����$c��OK�S���F���W_C��{��Z `�?g�5 ����r��v1��jdI��|5�d�c� Y�!�~�O#���1P�0L��JI[���$m���m-��G'|:�r獱)WTK�子]E��t�xz���b*�=�kt�����!�IH
8@J3�z:��TU�x�Rx�@J�	o}��۟�jn�U䖊��	h�t��(�G%��P��C��ڂl{�l�`i��x�P�|ܐ���a���x6i�@�rGI�y�9
x�"����4!bi9��؋��P���B+��6���R��p���/��ꉨ�p�)�0N�m(�f�y#�7����a�`�������D�ʿy��ʉ:?�&xv��P(�{�XS>��#�"�r�Md��Iq,h}�Pf�D2�;WK� Y�$8E��l�7vq��c=���/��L��	+�Py�r�phF���|lH�&�qf�W1��7�I�:��_� �!Cd�=GS�W����*�u���%�]x��ѯ(�"BZ�tY뺿`�h�$c5۶9�d�&�U1��S$	yd�FD���[?u}�S���?��tt���)����R�95���@��:�)�#9f�ko�	�7F%��j��`V��щ�����u��q4x��]Tw�2�D�gU�m���r���e�hs�'�Z�-d�>�M���ڡ@�ȍ3�Ͽ�U���, �榡�i�����^�\߶Z�	f�첩iY�`����w���(J7�����$w��U�ן���b!:a.�C��<�x�1m�úz*��ual�_��:�`�hD,6Ό�a*�I�9"(>A�B��+��9mױ��:����O�TiF����3?~N����d�@��[����v,��7���9����2�+3��.�����s�8�;:�>��OC2:�a=[��(�R��C�NƊ5�.��
�F8�����M����.���QJԧ�)!?��C3Fw�DͶ\�iTn�����:	K���c����m��h,�Op'eFB�'��c,VN�~!
T�A��A���o�"��9�Yז���-�i�X��#r#u���lc각ʬ[u���5������'�J��?$Rt�O�b��<�dD���-au �&�?H��1�}��b�f�J��9==_����o���B��[tX��V�v,��=;�c���Q�CC�P3k1��"�}�6Z�[�����kP�o�ۑG�f����)g��kպ,������O}f�����Zw����Jb��2��7���l'*%�B�����_5�Ϛ�����޼�'����/T �.�k�A���:Y�i�ӿV�*�˼o�{h9&��y�Z~�w���{�o�{�K(���Ck�Un9I������?��l�}oP^Ѻբ��]�O�ƈ+���-[�ۃ������	�I���k��= �4)~~?C�hR�k ���'x����;z��-�Wg�l�M�C.0ٿ�z+��r�҄K��oG��&�x�x��-X��D��>7�'���5{�]<�0���)���n�/4�Vz�QЈC7��Mмf��HI���_�;����Z9����@}�?��8� �����8]ymQ�¾�~�ƙ�Ԓ
�㐹� ���U�����>����'&-��CvR�����*?XV���>�U�"��Y�Ȋ&ج���d�\�z��z���i�T0EE��6�$E[��o��	�v�M3��{>{0�5�,�,X|+;��ӵ��^4�'Q������)Er�M	��ҖA�8���W3H�:-���x$W r���s �'�I��g�g[�;�v���F�Lۉ��6H�����^�N��[��5I {p1}��aT�/4���+�co ��f^��Ĺ_=e���Lb츳��5�/g�y[z++���U�^��5E"��l�lC?���<�y�JF(ؽm��b��A����ҙ���r�]�~���Q᎟�'}��D��77�FQI�Yĸ����e��I1���ȷ�8BJ�T'�['��J�U���Ƃ���.<�`�zy�ڿ6<����������"l�I�w��9ZsZGYFVމ�4��Z�3Ps�+u��N����R�/�]/g3v�f��H�� X���v��e �n�nƇ�Z�2<)�Z�����/��?��I��C��?�4�T��)���vIUoi�bFa�a$�`�I�k���+���s����jE�2�����T7�s�t��H� ���Mӏa�6�vD���7
���Vr-�Յ.p�����D��t�o��e��=�&�: �o�
�k?�@�[m��TGV��yv>$�h^��v�{�P����!\��ɈO�%���ߛ�=�?�A���rZ�V���	�1k��m�b"h�jE�0����LH5#|w�y|�eߠ�Do�|�1�b�4�?���%��^�P��1dK��Qϊ}S����E�o�:6-�d0+�+�	A�}��PqQ9����{�����`�>:�h��m�h|�POZ;�rJt���q~0�Ɗ ڊ��k<�@�������˜�եFT��	xo����B�U��w�����8Ҩ05�/�xqh�����G�12��/,Rv�u��]C\��yUf��.L�?�\1{O�q��3IǗr��l��G	9	�ޫ�=�g���S��:�1�I�@
�v����?#g�̉&�7(�G.'�7mC6{��P�׊��f[	��Ǽ%*�oD_S��r_ih)թ�1�O6�hZ��Kg�?�:2��c�<��a��#fcd��o�(�k��א�B�̽E���b�XM�f�6���竣�P~�w	��W ��)E���UMG�!/�rGپ��e}Q��I�H�]2�Q(V��A��Z��0�E#��P�A*i�����@�i0^6�3c#���=A���m��잲���w�nV��:̰"j:r��9��������9�p_`�^a��+ID� �� ��]���`���0�?8�j`�UYR�n�v_<H��R;M�X�T3�f�_���U�������[�H��݂���P3��c�Ѫ;F��G�c�d�A��uA˿\���� �ܓQ��˯��9�5@eB<�>Ntw��XV���"H�!�d? P*�ԿG��ң~"�"��z4�B��%/n�.�JL˦0'���I��ǅd�V~6�U�v9&���׀�A����Vg/�U(*I�\�;�U�#qA��*�`"C�TH;6K�������G��3�9� ��LՖ1�d:�7$�lo�x�����n�q��$~4L ��VZY#�m.a�Ic�����`�0�t��Am+դ�#]���i?w�SQ������񙪇�bn�i�xU����t�n$��PE��6��4J��V����-��8M�VY_gښ�G�k$�t��$���ؾVH�Y�!��p�񸢨Gl��>�ki .M;���;ї�N�5e������4[<X\VU����;�Ө	��sݏ�._:�dUD��%">V9�M6�+3D�x�.hv>DM굕�W��&>�񬩰��:���>[�<w`av��x��d:��7��р��<[f�<��owLԲ�u.;�ŪYw.�,�5���͇����`�>B����f^���������=p��V��s,iW��C�������l�.�y���2"�ݐbZ��+�L�+�#)Å>��W:$�Xb-�2Q�+bi� �t]C{�������.LxF���4[�XE�bˑ�(��w���䣲L�Ư�����ܱ����݇��a9̑����(��\�>}4�(|2(�Z�%�>\��{$x]@���ל����g`�N/�����fs@��o���	@���� e��_�<2)�+0�������ו�o�N� ��
؜���Ɵ�2��h�k�t�[�y�"׻���nLϊ�������C"FA�j��|�6���F
���,K��Vu4���>�R�\z�۩^�^i�`-���iל�Z8f89�1D�P�񦌳��ȟ���z����MGs�������\���t���,8�B��B�&���f ��$&Q��>���#�*��m��D
�}�.֬��w������y�bb�ԡ�d��C��B����i�Q#�H�h�'H�س��5q���,�l���Yb�0{�m� vsMm
4Q��u�:%b�Rh�y�"�99���YcW!�J�Q�c�`�2���B�q2��7Z�l�����>m��3����s�Ԣ��͂��0�����T-����	�N�B�& ��5ޱ��u(��R����E=��F���l�.�I���Ѻ-KgE�Z5 n��#,A�K�-����j�_����Տ8.%?>4�'�_q��l���Bj���2r����IRCly��j7&�L;jd����#������+>*$��@ӻ����s4��~�n.s� �P͒�v8"Z���02�mj��F����Mޤfr^���/*=]g�UšoG���������u��Pg0+��`��c�b���vw-��b�_�ɑ'nv�i�5w�OK�k�yeZ4|�k�/��|ڠ�Ы��°&(�uM�`�ܳ�>��C����W'2~��,�!�����R��M���<#���>�~�`���I�k��3V:�3���Vnbq�,YX�P{%�~b��s��|��`"ʀ���9ґ	�Z�l�]*g������Z�Tyr�6��z���k���dX��QO���q��x8v
V�ZN��VSܖ��s��Y%f����h�֎T��2�V�T�cy��E�R�ڧ��fS�.�z�M�I��q����?W�Q���`��%��58[Mό\�(������ާp����ݭ˜D�m��	ȓς��e��DPnCV��@�v�n,v�yF]�U2*��/k�i�\C'�?���Ĝ�拢9H:�N���f[���Q�d9K۹�?����{e�l�C:��À܏�;����.�kF���+�#�i$*ˆ��#��X(0���W�/Y�J��3%=�J���r�v���%����� �<�^����I�����L��ڀ�.�#�Rn\��2"z�)��/ ?�|��r��e;�{&�o�K�Θ�J cw��%�>��e򜟯��}�5W[��(ٍ�h=�V��͵�Nc�V6U���\	gg5�>_T��5��r��6��vR��V�]�tE+O2���U��*mdv�]��!zP�@O���& ~9�J��,_M&1����KF�j����O⁈y0�����Q.;���(��'����T?����qs:�	�۾Ld��x����{�J?��\�?�сW��HcKZCgw@	��o(�e�bS-fko$�g���yZ)��K0�gbv��ߧc߃V���
#e���3�n�,	R�z��K���p�q�vT�ƕ�3�����c@�'��m�$�-?��t������H;9Ρ�����㟖�L3uQ�G��s�_�N;�f���f8j&��)�7�Z�!t~mY�X��tKf�E���I��1�� ��dL+��Fl���K[�~���eo	��P�,Ҭ�Lf����:e�%H�=��)��E W𒥝D��
����N��V�BIƅ������
Ǵ]w�����7w>?Ɲ�y.�j �X�|l5q㓍��tK�l�gkrc7�WQC��a� �X,��G�~M�]S
	��;���Bt�F�h���GiF�qZ+����K�����Z;�kf@���~MUw����(U|L���W])�@`Ɠ�?"���9���i�+�VL,|���d�Q[�p�I��w� Lڅ�� �Y�c;�㓿z1zpK+��=�' �QV2(�3�	+��аa�)* )>�m"g���)�S/��:���@��`.ubg���VȅԽ���{x�K]�%~V&M�y-��D�J�\�d]��DSK���"Z�#�.�o����dP�;��X~r�Q5	�[z�uz��c�~�����jU4GP����b�*��H�i��rCɟ��OL����f��ťLt)L5�!�b{���D�V�i���U�}��L���e��\��nk��_��7ī:7N���<�ۤ�B�W6p,#{up�{o��Йt;�4�n�S[��u�9�����O_����x"�����>E7 0&��RP���Ύ����ϲÝ��#l#�Q�_���j%��O�+w&ž�x�Ā�+b��L��qY��a~Y9ʦ3,�&��
���2��!�T�sr��N��^Ӟ$�꼄�1ds�H�<�U���� �p��9�VJݍIZ>�~�ō����pu�����?"�Ozܭy�"��T .:��E�h���Q߲��۷Ot��m�D��8Mw�.;8����쩌T3&���������mضe'�N�x�QZ�#i�"�����'�ok{w <Wd�U>G���iYMĢ`n�I:l.x�p�Ū��u��7�_s�����x3����:Csҁb#c�>6H�2���(�݉���U:��|�>��;a�d������̂�yE���ĳ�is�m�(�	<jݛ�k�e[u?̝��C��u�֐��ϙ$δ�L���x4=@2�`݁��԰��Cs^ ��i��\ǛlϹO']�I���`f`q�la6kRvw��U�!�W5e����$@>E@|4{�/W۱,M��k�3 ��Åh/E�%��s��R�Pp	O|z���t�P�Q�M��L�a+(�(ж}�9����s��RV�u`@�X`q��[i��m����X�G��N����9wyФbӋ�;�;4t���}�5�N9_VWIf����(}���zC�Xy�O���ǜ�X[��ۆ�a|��͎y��K�\њr?*���j?��k���3�D���jưr���%v�o�D�ʇ��'���09e�{nI�Xğ��e�G����lC�@yF`=b�o1r.~z�&���K�����*��S�1���[�Wv�%��{[I�������%\z�T/k���$����b��W,��`��T� MV`7 ���6�0�O�2�ζQ*�������������CB@����he��ǹ0�����<O�7 ���uԟcZ�A��j�)4GZ�7�l��'Ԯ����h�rV��|b�_4��̢,�F���i4����r�m+���vng����F�	��%�6�~Q���=�T��_5`ϧ熙�R��2B �!���H��fv84�kB"p��	oy���k�=��>J}l� �l�>�!��/h` o}/��t�'���'tAw�,��ua�p~5��@�M�-XS��]��Q�j��)J�j��W�� [7����_&(����`�2?{��F�Dpk+XS�LE�9;�ɭC���=;ރ��D��l�;��aI�Qu�Q�6���7�1Ӟ�57> OD��Q�X�U�v����v���M�薏��a���͎d������?�[�6�cA{Ї��'�T����=K����y�"?��
΋F�ړご�X#�NN��;�3G�n	�hu�{z2���r6~[
3��pG(o����
\qʪ�Ե�_ɮ����/�>����p�^{�٭
{��a*�hz*Z�X˝I������g;�������v��e��Ǻ�ZY)���ܻ��f��C��갣*�k��Z�ԩ�K��)�.e�b�Xx��n��O5�&k$�Y<2����~w}W��_X����zz�*��v�t�{�����f"��b�a�>_�s����z�f�!h�S�E����]!��W�f���k�:���|!�|���MC�;��_O�<h'X�H��|yV�d�A�!h���-�N��#�٫y�T^�2FF�Ҡ9�|���7�P�t{h�ۏ+� ��ʨ�0��>:D*��T�0jV�J��(�;�zx�3n&�z!������n��sfl:#�'W�H�ũZ�j�|Y�ހ[z豎��7h>[�2�8�S�y�	���N&&a�9�WF��[!��ז">�Uf\��N&� QO��'��f>�{�4Y�1��M$�F�	�B�H�%����?�����}��fqfS��b�MO�$������.6�r�0�+.��]��5�M�O��c�%�`a��M(VVj6^������LI���,�&��Y���d��L��+�*���]$Q#���������?F]�m+?�t���!��@�ܵt�7B�X<�@��HI�?W�d�2^
,�t`�ؔ��O �&��`���ն��q��g�c�I���˛�(4��>g=�n�3���kn��4ǥ��!M؍��6x;��Y���5���]Un��ҭ�#)����*�*���� ��L
��JPi۳�N�zS���@]��/�"V���EJ/d��ۼu�����_�$ju�j� �M�2��)�}�ſB[n#�pޞ#%� G�����nǈpl��ؙ?������oK��T�)b$|�����9�^v�����)[����o�8�b�(N|��NWs*և�H�Wa�+�?ݼL�G�Z�7���Qjw�C��U�Oe���9�4�(H�hPuk��R9�t$���:�/�+ޕh���8a�'k�/��雅��k��v�Y %`���|�r��vYx�yǌ�"�!�p'�4\\�?>��j�Lm�A��8Q��M}6�ïT%v��"���~G���~�x=ړ��j6����ّ3��X�"6TIפ��밨��@�a�����gI����<3 ��5I�JK�.��i[[���_]sE�<�ȟ��?Ǎ��w@=EXvX���/��t���R1qAƾ֐��5�Դ��S���-�qڐQ���82:�oT�����֯c� �8�`e#C�����	g#k�M���/h�n#�i�L�q�U%��?��T�\Ewz�{�d3	�%�����D}�%nD�5�������QhA5�ԣ/�U]�㊒�ߒ�3�{K�6����O;g����8
#��k,(>"�c���VbǶ�����٘@��:�.� ������b��� �������J.��� �,譟G���s~�����v������SW\>�t���yv�3��0�N��aʡM����ڙ� %�GǃG�%�7w	3h.d��%�w�@�� �O�͂W�jd�)x#G��RWCtY�����6p�Ysl�'��|H����V�>��ӨYRgAAx�c���#�E68-pś]&�Z#ѥB���G�H'�	s���g���yPk���v3��%}�������ʏ,�X��>`��U�m9�Z�A4�S���0�]�V�m���V~V<�?����K���4��M��T(X�omM�>��.b���{C"�K,i`n�ź$��e%��v�1��sOl:K�g��Z溝�m����}�񳤥I�����A�x��*���n�;�H�����ܘo7��n���!��rd@��x�xuc�%��h�_�%@����k�j"����,O)̸�)�^�Mc�I!\�,ZM�ݖ�FA�SZ9/����p�}�4_E���@q�E"�����E#�-�M�Ӧ\4��WY~�p&"����riQl�걙Ֆ���5L�g�> Y�$_&��m�I��Y�I���̹��f��K��6������<e	���T�shv��OL"0�FzL���J� o�˅Z}���|�f6;Y2�[�f�����.Y�������69���a]q���ߨ�����L�����CI�2��u��@��`���B��M��_5��5�n2Ni �
��'����O� �H\8�!4�9��~��=/"�8�
n��@� �k3�dTfF�a�4�˃V*��&9��k�PSV	���y����Z���W?��6x�F��ު�
	�'[ S��.d��5�\!66jOW�u�jrA��{���4�bO%��e�ځ�EZ>g"��me0g1������z�\�8�� �x���Oz*��9a�'�c��8o[�oqU�� d������=3Kձ8�%�#���z�pǱy�#d��Rb1�����H�
�!|��34Yl���8<͚���At=�1�ز��Y͞�Y�L�	0Sp@�n[��RQR��O��F�s��]X��7AG�&i_��_d�&>��~��B�J�ũo0�� x]I�AugU�pl)�s��y3
�'���C��,`}����&Wm��&�M�Yx6��AK _�}�v�%(dML{	��d&j��av���2������,_=M��:��Ҝ�Љu�ٝLf��D�J^�L��~FG�����R��̲~�kQ];�9h�/����*KB��݅E@z>�2��X=&�q�X^�` m|��p�'Z_b��<Q�6cE�� �Z����e�$� �� G�|�M������M���J]���f���dz��p,�#��M*3��B��П�O[$h�fp�GTn�9U���I݋��e�*�a3�rX ���{�Z;�U �~�\cj9*z6P�B`�x�"�O2����T����\��f�G[	�ܪ;��mLl�?.Տ���s'�	� ǊLm���� 绖+ݵ��#�|�c��a�5�2�#�)/`����[2G��(��&�v��JS����0�/6N�b�t��fPP��U��-�r�!{�R@�f*N)�*�ٹ
����7����JRI��M{�,�F��+��A�2�v����ś����GQ|����P��;_◊�r���L���x�����֙�4���,����}lu�=,<� GQ��:�ͬvB΂G����p:���ô��)�/,}�:bl�tq�Gf��Q��F ,͆p�����W�xt�L̠�dN��꣩�wˏ����b�I[!�a�?����IL�T!$Lb�ޏ�`����W�9�N���d�2Z�<.��T���&�B����f�����ieY�9j�1i@��n��(�Ǐ���(�5�/l�d0Mg�<�=�cF���D[ڂ��= �@�n-�ɺ�� �]��8T�$��j���K$(')"D��(����<K<}~��%PN�]
�����7�r�BLiP�dM���=]��(��X��_��}P�38��V�]t��t�r\�ց��ќ��f�1����8�L�h������B`�Vm��s�漍�)zj[�y�2���+U��gu�_���<k�E�>�jwl9#���� ���<�K!� �����&��kp�O�ʐ��qJL	� <���A�3�+ �C#L񿐯p_�A����5���'�E�t�9�84������X�ʠ�ȉ�~<"��Y7�Tz4-��n�f�fx�1��jA2x�>�E�u�����2�)D��Vq+ѡ�1O�j�XO�x�`O}� m�q���`�ǹ��Q?KT�t�,N�������J�~��k�k�D�v�dQ�w�vg��cfIڣ��-;�=�!�-�\.�W���qfT.u��"�/3uNh�k�0�'�ZxH(םBn�֍�Z�^�b=V�?Kg74
SR�鸳�cM1�#�)銚�Fl4��)��LF�&�FJ@;#Ы�MM�8�F)t3wS�S%���� !�k����(���u�v�3XJNY�r�j>t�	���%�}����$yp�n:0����h���1�VT����+�0~|��4�Я��
�E�k����w<ޙ!�+tő��n|ae���ǖj����#l6�<W��B�Nu�H�Li
ʍRBЪF8��
[��U.!�D�/ v ��e��i- ��,Q��@FS�723�|�)��K���q���a�y~�������7��6�塳� �9�w$%�iV�Tt�xo�q��(]j�^w_�Q����z�+>4Ǯ��X��-qC��Q2>�!I�m�Ը���,*��'Ó�I�3?��i8O��p�����I@us����������Y0/6���|�}\;�iG�����!�V�G`�]��T0��&[�84Q
�G��#9�Jݚ=���KH-�6�Qa�+��Ƈ��?��Z�d���k$�얰[���fH}*Bb:�$JtM\��8�+n��-#}J�G�WA��&����C�M#\*��n�aǫ�ł���G���ޡ���P��m��/nH}����M��qǉ"2� �
7�K�����,`R�znS>���T,i����
G���H��,�i��$�TUފLp�	@��zf���Y��N��ļ��-�O�1�¢֙�dHSx�v�v��pE����V��=��xPU��Q����%w�����2Zy4�m�}EdK�TT�o�3��cXpN�[�t<��lYjX��8R�CmC����=D͡��b��:���ѡa�+:�����$p�e��u:y�ɺK��,Y?�N�N�=dc#e�ǧ��2��|��
��_�Ҹx|����W�����Aʂ[��=r�|��)�hp��} l���OB-tx��\<f��	���*͒R�,��=��V3(\#�ip��3w��u�vʑdJ��䴤���1#l�Ga��K$̟�S(�����t.9PgNg��?����LF�xq[�]o�"nB8��ݙ�ԜQ���S��_��p�t��f�S4����f(��;B!��xw0U�3���n���i.���iH���Əq�s9��h�	8���#�,ⴼ8$��>�hҊ�c�M�Q]5E3�"�J���T��`y�|/rV��֝c���ثU��xhM�}�b��:�"�u�I��!��e���&�+�w�s�ޫ�J��ku�&zx�l�Z��O���}����E`%��L���f=y�Θ�+�Z֝�(&�!hth|����'�d��X��{�=pB�Yx��	�9)�TW$z��M�ȳRѯ�i�LL ��}p���%�Ɩg��}4-����f:���4;�c���ܖ�'{Y����)�M&���?Va� �<�WO�à��|{�ᔃ��oe�����H6M� \i0�W��{B���v���H��@\.I�Wu�j�2�G��IQ[��aK�����EG�:>�����~���k�2�ȓ]�v�k ?�q�;���c�Xa�Ʉc-�VSv+�