��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\���V�fnvx��ÍG_;�ȅe�~�>���9�>��Y;�0GN����Sl�Dg��r���Ik��
/J|Y������5gkK�W��.�mR�gzO�O`I$V�{�>^�#����<h_�nSު t:Ԅ31��e���������;�����#r$���\)
M�8�f�@�����{}�qX�S�k��(���}asWҀ�Ǝc0�Wp�X�.���bTS��r;Ϯ#} `���'�A�cl��f�<�O�mҼ�gI6�&����.\�z�ːg�Ll�*B3$-\����F��V6��\���\QL&v��k�0d�����z���v��:�8,��%F���}E��N�
.%ݹCQ*I2����"]:1.j��R�"����5D�.9/����Ə{
�r�ɣw�[��ڃ�AFF.z�,U��}��s�%no�y5��v�<���Q
��D�����/,�
������ � 5;��P7P��,�!��)4w��P&��~��9m��	t҃�7�Z������L �zŻ�6D�������Q�5/� �D��`�$!�t�-��B"��~6ЉB��f�F�|]`1X*.U��d"ӌuIZ���a�?P��CZ�t979�(Tۃ���]��2�����r&y�͌P�3��N!��g�Lٱ�W}f��)^�O�0�w�m�I=	�G��m�#'�:�G���f��[�κw4ADfrQ	�0UW(փԧ�Gt�!�5bq��O[0��)W�������8�u�d����̐���7m&��̙l��X2����2r�	�����;o�q�x��o������|��Dp	�d{�+���\W�B�!X��+�P�D{��=j��t��t��;�ًn����;-X]W�u��Ց��ի���1�:�y˒�@k`������a�8��ۮ��q���dg�zv����������X�c~�tE���ñ��B�C����	�g�P�n�V9�O۾��y����̓~���J��D�,����m��8Hl�OB(w��z\D�/�����D�m�c���d�P������ٶK�w���ai9�T���`dL|^TN>�$�j�MO/Q$}"ͩJ4뼗�}��~�(Nv�ڷ7�.�d�H�������a�yC�f˕�>�}>C�e����F2
�6=-���Z5����<Z�����]�I�G�m�)��4������.���/���r�%�A?���VpF4.aIf�L""ej- �#��e�B����&�K�"��M�S �Xx�a�8hEaÇ=����I�&�6��h*���ʤ��ޏxLՔ�鳞�$w@�� �`��W�B>��� �7^Ԛ��s�v6'���+�jσ���!��֓���X�ѤvU�XJ�N9��t�%�:r�;�ef�RE-]���mض,�Ы������ð�lD�W��*���8j�AC'F1Y��<	2h��t�喬�١��	7�]oY2W����q@� ��6^)�I֥4*0���H���ң��lձ��Bx!E��N�;zm =��/R�&�iZ�m��E����� ����#��Q�	UK@�{f
������>%+��dG��E���#X/Q�_3��䲟�o�ἴЊ
e*�C �zn��|e΄������}���������/q����FX�5?�ahL�U��$�K�닙n4��s �#�o�=���8n�'q'81���fH�^�86.���L�E�"��tf,�&���sި�8��(r��]�^J�E��Cc���x��8_`[D�Y�Gؗ\�����z�~=V����t�����^�KO���#tͱ����[����B�%���(X��V�l��Yo�7P�NWf
���v��w�'`Pkt��{�9ҭ����%�}�+L�҄oU��Ilf�V��>�aI�u��ĺ�v� V��- �;�fC�����}ƞ�&e�e��� !��Y�Yꉒir��8�)W�1JVS��ʶ�	�~�O�5�z��6�Z'C��X�A�י<$�W�[Aw�bX��W�v�}�!� ���MW�`<DR��R[��B����u������<ꅹ6f���4����š"!�(�W��]�����LV���b��_2��cx��aTcT��\����&Q	y��L�N�T(ߤR_kIk~h�t~�/E�#a�%���>�kQ	�}�Z?-덻`�t2"$�ǯ��>Z���C�=χ�P�Έso��Bx]2r���^�,����&T\�,ܢb��ǯ��:��`�ia��Մ�{��Q5����S��m��� u"D����>�L���%���O�'�|����K�����r��Gt�C���I�#f�*`�G�E�slb�W��pV�%bV�G�6h�5��eR�]��4嗢�1+	�ϚlH<�����*�6�N3�}�<��B�xjT�o��5��Y ���L��
��,��:�;L�����?�����rQ��0������� ��zv��ǃ�hf/6B��q�^$�9������!"��`r��y0&-�-��)M�!���y�/�H�� �:7���g�C�'[s͒(�A�S~h*��|�Pp��VHh��W��,�"��ԆɊ	 ��ߘO��o��;L�bW�;8�	������j��@�ޟ�2?(-f��y)����r���Y��[X�bP�N;���N�Ҋs��)V���?-j��a1������_<�~'�J1��tv?��Ob5Q��#��s�;���D��3�8�DJ�RJ �[�������Z�E�;��Z�`[g�^�Q�+�I�]���oe�g�T�#�b���fjKy2�"lN���`���� Xa���v�_���t3DTaЛ9�����c_��c��52�Yj�j�Xke��9�a�'��K�[� z����C�a�n|}D.�_�>�
�I"��� ���_��,�Z�$�*�>�&�*=��P]�#�|Q���2*J���޳�v�ߨ
b�ȼ�7'G6(��IU��o�,tL����$rtU���v����0�^�!ֆ"�y�OuF�+�)�|��J9�WI̼X0��n�)�J��g���X��|��6Δu3JUp�<1�y��Y[/5�̭M~7��!�c$������	r�]؊�O�ƻw��O��#Zd��3���Q��\��I�h����ף��3��<������ڀ}ۯ��rf��oT�%fŗNA��'n�k橗�6�k�;�C�30�B�\:�u�a�
<;�G�]Y$ϝ�*�/W�!gǼ�W��Z��X��ˋ,9�H��m	��]"�
i��mF�#Tbnb-<�l��P�{��Rc���lDQ_�zT|h��3MҐ��P�{�鴹���}.���d\?".9���=�*��2eY]N��)��9�i�pr�&/]˕��PS�j�@���J��w�ǔ��[D���y��L�oBF|��q�������e��0�fǟ����q)a�Z� ���+Ze���j\)-$Of�n�U�#`��ʡn
�q�J&�0�䀔lmǟ���q-nڎc��kÈ%��(y�)/=8⦕��Fuh�����H��+��!k���L3���1��,n�[�>�w�!��� l���8&|�iB��TtW�Kx��C$`2�u6�ڢ�x�cSK}Q���F0 .M�#�`����D[��y��S���������bA�9�2@�p���|���R��/𺚯�9G��Z ��x�U��Y�0p��� ����y5��3��X{���-��1�w���t�x��Tj�I�����	n����֨������]}��a��p@sr�a֊�`��8�Ч��`[kȎ�?�?��7��ո�7�$���MC��4��;�:�	�H����w1���&�#�:Q�aSr^X�2�
 .�����]*��7�5�*f��&�1����_t`=`�����v���gUqsj$ٞ�����_�-p��ʗ/�(^ 䊤��/?eY�ls��X���6l?ڡ�����U�~�]�- ���7� �	X"z����j�l���I�a+�z�p���8�!<�-�C�g�+}�*$�/���R��|�9L�ey�6�덜����Q6��m;�d\��n��������9F��r�����*ň-M��,��BC��*Լ���`�IDx��
|x����}�Q�
���w��&qr��.�ٸX|�'��D�^��t{/�a���Ř�N^�/��W*;-L	���i(v�p�D�%��CU�⑙�h3,T��k,�I&���B�9�����qR��zaӮ������(�c7ػ��Ok9P���:)�����t�1����w��a�V�eu�OD���\�_m��u���	i��47˛�F�g�I�M^b�}5A{/�R�,������g�ˆ�~6�/'�K�w���OH��]D�+�G�$K��=�p!���^���?�x���"mFe��[��էiT����|N����E�to8l�l���a2�Z�Y�j���%��ꋊ�q1�KK|䋾/���� 9;�5�jt�K�Dh��B��y;�VJkQ��@��6���H�ÆX	����G�r`�*no�>��j�p���v�>�v?jJ��i��X5�Y^:,���T��R����TX����쥧z �cSZݡ��$�A�S��c�O̶Y��2I�bY���s�Q[k!�f�fQ������'��ǭ�2�W�٥��(��:���\h��l����Fa��� =�N>\R�(��^;,yQ�e��9���6�e��Q�n�A�(}J2l��{�|�M.��vXa1?=���;�s%3�p�}�5]�1�+ڧQ�Ǯk��ܓ�v�H�Z�3z����%�l���%����~�}�8r������� }��<�{�%M����@�P�ɫ��I��8�]���K���gˀ;��~�K�<��H�yUt�8��+�l�(�PMi� @i��qf�N^��j�B�uV#�h�Lk���N>b��Ϫ3½w��S`���,�WE�����k	��I$H9�#�C�;�������*|�5�)v�~V�u;��-6,�����6Cj������a�� �X���3C�k�藶 �|�Đ��C�L�"��KD{�d��l\�T������1�����U�dx�3�@a��n"!x*b��sH��[%��m�>��8��8'?oT�`4�F��eTJ���i�7w}W
Nm3K/8a帚ȶ�jU}y 	�B�zQ\���9�J\���^1�����=~7z!�L�ϧ�C�!��5�O�i����1�㈶��|���T1�Gj�����^�C?�RAA�˃� ���'�7r�Kˬ:>ң�Tb�̆�N�*��f�	nc�.��"h~yY�.���ǔ�A�(�)k̲C�i�&{��N� ���T��|�ϐ�shg��"h��>�h
q���1�>�ϸ�u�Ջ
p�O1�e���d��0�1���ؘD)�"�Q���@
΢�$o?~Ɓ׃-m%�/C�����(vǳ�EX�L)���!6�.y�EF۴�b:t�5�HF����NQ?I~آڀ�5͟���
>q�����%��/���S?�X~.X���c�.�5�-�jj��1k��`R�đ��Ҽ8=R��D��ޞ�6Z��5WU@g�i� �u3<Q�gkX.��	&hqN
Y�+&Ҫ�6oQ��k�VDω&�W�V�4^&�U<Ɨ�>T� Y9H�p\g�gd�*V�co\4D��y�djd�Sn�~��0��I� �U�F�<�����?�1��C��x��ܺ���CC�j�Ba��Øz�1�C����KPf#�[����b��������(��e�+��Q��&�5AL˗Z�R����S��Tż'��]����ܙ�8;����׾l�6mUږ��_�5�l:�Y�]����%�ԗ�����܈l����#�/��AK!h
:[�Ѽ�����:,)�K	 ȉ�y�i�i�� 6~���m�1]��BWxK3��2�8��{�`����y
g���MH�n�}M)�����u�A���xR%CEVn	���k�m�yA��M�~ ��Ж{9�ܚ��4I��ݙܹ��Sd����iZ�P�,�u�����]b�560p�~��-�4��%�����B�*��� �&�˓TF�j;3�
���a	�;P,�%pS0݉o��0�:��(=�&S�Ʈ�@���Pp�m��>����,)��`�p�uZ�P��Zsd�AV��5R#Kg�dӜ������Y�K�z��
�:F�Y����y��n���J.%�N[M\��[�"q��9��c�Q����=��]
`��0�q��F���°��.Ѥ�'���/�����a(Oܓ��h���>A�$d(!3WX�G�E�m�����c)�}{��MX`����ł��3��(��9ҧb�|;Y	F]��׏O)Ht�F�. ���lOw��w�a��@��"ů�)��1K3�S�eI�dL�ol���tEw����h�`�Ӭ �hD�T`�o	�PفN0�2��ϟ�`�҆���z@�k�f*|a_O˹85�������^�K���b���5�(v�a��{56��4�k0K�ѷ�R����WOu�m4������Rb�Oe2�-��_U����JH`sNR�~zxw�d���)J�[g���5�"�Dk,(�ľ
�d���a�X���63�s��1+_��Q#x����4pl�돨\c99��3��E ��w�}4e�X>э��[H^����m�X�^HX�j�@���� 3�0T5�N��-;�}c=�$~�5w�KJl��6jR� �N���#���CI�}��2ł��K��u�YO�&�.�Cm	N��
�>�u'����֏�^����c�ك�
�]k�ź@�ⶡ�ފ&o���c�%�I��EE߯�/(.�5�+�	14����yQ5a�xWU+���ɟ0��7�DC�U$��t�O�uB?�
c������đ�l<X-�������I�:v�Ek�7&�Ď���MfT��p���j�|'�b�6�%OJoG��뇲�%@#F=�u0���9n
�>���\�p'$�f�H�s�w����[?̈	��?�-Mm�HI�(��^F	�$��H�� �����Xڭ�_�iv�:3J�/ޯj/k�݄>�I�(�}u@��� �u�h������Dr-��8����e�Χ�.'<�
����uB��!�-&�� R��[���P�S>����|�t<&&�<_T�P%�M��"�4�gF��T2�h��߲�?I@����dk�� ��x�&+�W�����캐>��Y���j���Tݭ�-�~��5�3�&?��s-��e��z�]�)�����ǭ#��:o\�2����ڕ�{I��4dƨ�o�ծ��_0� ��WO!�A�SoD�_e��gǞ\�H>F���9�Q�T5^e��}<������v�-�6k��ƾ�)��65N[P��$����Aڬ���B�a����(���I�����0������_���3#��&�DH��f�Ȯ9�ͨ
�`��ܶ����1�H�6��|B?���A�(�B�Qp�!��S���oW/B ��J�s�TnLF�g"|d��d�r
|�۹���P�8#H�'�u���M�;yэ6����ʞƈBYF��k=�y\י@�T��X�v��"8ƛ�m
J�� �B0Gl�m��,����:i�'	Q������wm��so����;ٗ~���kR�A3��t�������1?�e��&��[�����׭ ��Q�� ɨ�=v��垍_h��婎!u�]�nG�\7�E4b��}1��ZB7I��k*/h�����1�ɤ=�l�#�=bjV(Q��ʅS^��m��&g��ºz2l�ZZeJ5#����Qx��A9[��rD��1ՠ2kH�)��T� 
A���ɛ�>i�͂O/�K���&*�S�t�F T�7h	���h���E]ׯ�B���e�@Ipg�a�}�I��<��D�i�-2Ҙ�n:�����c�6>2rnz��l���X\'��M�JYZN+��[pw[�Kv�G������R�؟���i;Yx\ҫkE��u�4W�ٖk�����L~M#��_$��� N�����uDQ�D�P�[���Mg}@6�F݌�!�V�<M�}e�����[,�:�d�MM ٹ�sSc�$�����}:%<���z %��R48_2S
&)���E��S3W|��	�O�㥷s�	�~��^�&�-=6c�S�U����XBr��J�޶*���
�(�n"v��a���:ϼXb(�^(Q�ς��
 �yL�>R�YԊ���BG�=Py�'�aŝ�J.�T�A]����RY��pxP@yq1�;ߩ��[%bz��Xn�zgpC��ep������4�
T�0�a23��a"լ��V��?�TZM����&G'�_�����g�����卪�?�[C�1tH�5��aN����\�$�#M�M͵�3ƹ�Y[~�, �wfb�������%$�]����[r��R�T����`§�W,��w]VP����H�"��l�cR2&���Ou�dA�+0��c�5E�]:{dU])�/�J�+a&��m�,��ⓠ�(���ß0 �Q�;�
���R��ݺ��Wla6*{�,�0v�؝���P6���dڌ�M�2 v&���h�{�����!sV�! ���H�$�'��`՗�SFW@��>�{�I���>�9���**��Ī���P8İ@ ��}�@̟>���ꑳf�3$�K-vX��͞������g&�� 5�Cv��f�����eIB�qJț��Tq���ωRŵ�����³��Qr�����WI�M!�,�K��h7<�b�#l�|�tu�lI!���X�~��X�5Ut�;
�jA͈<4!�Z-�ۇ���ԑ���zm3&'����:p�sd6����Q��hε�s4-Lk�T#�4�����ˁ8�$N�<|[t�?j����c�� �8��q2�"�9�f�@`����3�bݶK��ݦ��b�H�wA�YV׾8�[��1ڦl͂S�1-.c3��+5�M�ǿ��(��ZsPⓚ4t��%g&#�;�U��vU<P�ʵJ^n��R���8��բ� ��=��׉ZĚ�jH@XG����������沣���ҫ�u����,�ث����e&b��B�?����*�
m���b�x#�JV�����SjC��[�<���˓��i�W�Q�,�ou�cm� ���@��9l��y$��-�Pq/�l���F���6+d#~�ʙ�V��g϶�89j�����HA8�yԡ���������Z��0qZ��j�$u�=�E�-'���bl�u��4f�8�$F�Q�4�"�tR�!��{�p멪�������艂��3�V?�����^~��Vp�+���R�P�q��ll'��L?����`��' M �Zk2È;ϫ?��pK���ə)Цv��DU�輣=5)$�C#$��Y�c;�l���.}e�V=ps&G��4Nt�?�yM��9���Ψ�;֭��.t5���|r��r���m�[�X�r�mEh�ϗ��%A�!eQY+�@���+tr�������Q��i�������ֳ)�s�;鷋�<T��ϵIxs���aZ�a�si��MRV��$�f|/�4���2���-�8��MB�6*b}���v9����=Ag)
�`,<��	�)�XSw�֠�ơZ�'���2��?Kz�&���U���x?m�s�&2ɰ	�E,d��<��E����|G��u�}�^#�ݲT^�V���r�^C4z�3(������#Y��*�����HF?勿��^T��+O��5�c�?֑�-9Z�$��C�C���>��Ӊ,�;(�ڱ���	͗�4�9	�L]S����T����c��kJץ.�PNA�?8�]̃@f��q��*$�b�${�B��I�x?��-]�����	�RG'e֣U��G������;y�9{�<@e-���8=%����%do�g�Am�ۆ��E��SN�Z֥4��n���k���A���F�1	�bp�~�*(��!c4?8TP�vs��J��\����\�9C��p���aQ�X�֭��e ������O���Q[ݰ�h��
��m5�8� 8}���WyINcʥ��h�>*'`a�?(���������Gr�Y�����s?%OD��]����䐘x��4�j\�pэb�Yb#5&�����ּ��<��j��Ϲ�ELe:D��� ��`!c�ZgOG�KZ(*�,|P�F?�fT��*r�������-"!g>#�,���ܷ���qg	��� ��&g���v��'�[̖�ϟ���L&�80w[K�f������pⅽ�ר��,��\!�v4��E�zx�7�R4��=�H����z֟��4-9����Ș�e��'��T�L�,���op@#*5�a��@�`_��WL��52>���������q����$0F;1��;�))��%�%�9���r��2]��뷆�8��e�J��=%8ko&֦�NBe�`��&�;�� ��-�W��L> �K�Tfx�D%���Ns�1���jiJ�vw�@ZP<�TA�Ɵ�V��x�u*�+vH&	b��z�Kk������6�tM�Ъ�6Q��D�&O�y2Wٛ���<�A�,E��Ҟm�%(W��Xl��pMPՅ)� �Sݶ��}
󦛆��~?���㉀1���rNj1�2&�b��؛�J�R�<<Ƕ�WO��aG\��fP)� 5�+�15���!�9=#��-)]�	����� ��%\���(�R�6�������d�P��g#9!h�ՃZ�������G���\�0lԽPBD8��e�+*3��ǯ>$3q�h;&P#�ͪ��ؿ{"�x��.0+&������(����lxo��d;ͼ��C
݇C���$i�s�qXDD$ӷ�B�H�l�d�)�#��c��U���>D�Y--�[H�:�U�@���m���4����-��1�}E�k��,[n��?��ފ���c�� &��$�pzC�~V`)\�۸�՚[ԩ�,o�ݛ�/���Čo�צ��@oD��=!����?�r3�\2�}���|cm���6{aa��X�_>Χ�Z�3	��j|�eh�}.�|�ͺ+�GX��*���H��q{ME=U��#⹳
W�
�R�Ʉx�q؁� �x��	.\��Q��
�gW�Bq=�3�7@��=�|y�^oTX�kG"��q�x˴}C0��P~��,|�μ7���Y��1����UN�Zvr,�DBV�+�iARxM�GtWs���1���#����i�~�I ��'��v�a�j�B��if1�Z����1����{v�0!�:|�Ιk���O΀vƃ��Uyi���?ȍ���魉aMR"���&��?�I�n��`㝖��o5�nȮv�}s���Y�q��m�@׳y���<�|�'B��χ������$�L��u���[[]O�K&|t!!�F{'�����Kf�wrj�����������u]�b�j\��6��hXo��Ӡ�$mzWK!{��	�P��(�g�����6���^�Am����"�UI�˾Fo1)�yؙG~�1���x��� �:�њ�2!��\o���j-���.��W"7PH�D�$�A������4��Ty��}M�_f�4Op�a�s@��VE�ꎉ^�X���N�FD�;��pɪhu99͍�"�]�J���@���I�e�bƯ�TH�W�Ƽ;̗�:x�����s��EQ��d�gZY�dk�鿉~�biGt�:��i��@�������J<b����4uM[ p�Sm�d�x�{a���4M��@-�X����ꋮ�B�M��0倁:U*��X�!ܞ�t���pU3��}`<�X�s'��w�_f1D�����Om4����q����R�G�����I�w�e��,��S @�oF<�5(��5�?a1n�����f������e�"5�V����`Fd�э�#CZ�x=��*�+��X ҋMr�����y��ҤT���e���U�=�.A���R�,l�rf��:n���G��̘l�m|%ωvs;��,�_e�Mov3���(2B7dc"vJFj+�tdhI�3X]��t�6��,�A��OB�~I}���y]�y�����)Q��Ȅ6��Hz=cQ�cq���!�6F_�����1�v��q�餻�T�x���b�k��9������㚩�(Vj����v8E�*���v6l{�A�����рՂ5�4����nc���-;U"�u����W�	׊q����㙓`;��b��0s��k��-U��:�>�R��%'Ր��M��V]�A��S�&��
tI�����+5bU52p��н́�UBvrlH�w��>]t�}��!R����eg�M����fCǛjDM`y쐻Ǽ�}7r��T�F�:r�*�{�)8e�S���4�u����t�%>4-P������џS��T�Ř*��0����G���u����X;[��I�5�ٷ������Z��(�ޚ�p��y)�c�{ݱG��o�"2;W%���o�kH�|��{Aj�VyT��v/�	[�s}����9��񱦪�^ ��+�萅�dчP�UU@x�Ο�<PM>�?�P�ۡx�D���{~wKI���r�%�%P{M.��C���ʸb��Aq��?��0\��K�9�U��_T/�J�~K�}�`o�ѐ���=0�n�3.��N7`Wu��9]b��0����TL�d؋���)���A��T��-{�X���PUUa����3�5ڑp��n]]����ⴕ�ͽ8P^�\��yZgS�����w�<�75��<�s�A�-@�����4��-�49���3�涢|�sA?g��-�AU�4�`��~�zV<��x=2Dd)���K�eV?��b��ΐ,��hrm�_��XIƉr�{��g�x��/� �(�ܮݟ�'�7����b�%����� RG����uJ
��������2q6�zx�z{��@GO,3ؐΞ@A���.���x��ݗj}\"���������~��߅!`�M��W�G�*�:zݾ�Ղ�"�KGFe>A25��ɶ���<��[����H��;"�����vwEJ�j�e��)�Ix���m$G��N����y�j�u���޶~���߃���	�S�
��ƍ�̈0 ��Z���*�`�o4��úfwX�_z�>�Qt��!\z����U�KB��x(�����<�UO����8�VK�r%�^��h�45ճh(]��f����et��Mñv[0W���1�H�6x[O����u��� T�+roT ��/C3m*�m��$�X����T��, ���^S{<F0��娿���mz�t��\<YN�T�{KGp��F�QB:�DLM�nhg��+�ԜGdhu躮*,��ه���_��S�u�v�RF��
���-T������u�Ĭ�ľ����ޱ ����ޘ%u+r��:���q&��LM�w�M�m?��=� �TSs���p�[,��\��~��'1��������H��s�U��$�ͦ��q'�1�8r}HB�%uX~��VK��G�Z����y��R��*�¹Q��v0�~r5ѹ�"�e_�S�6X�K�HH�"3�d��Q������ljF�U��ۄL�f��^}d߄��R�9-�>��[�O=��q����� :M�
�8y��k������0�g.J�܀��E��-IУ`%��O5���3A9��5ҁ+X��7����ΪP8�o��&��f�J����m�U�q'��֚����*�2���4��r�>Ԙ���!#��h�Zgٰv�D��DE%�d���|��3{\�jH�DX$)pnÛp*�d���.M��"��x��Tc[��I�j�b'A*���� r(&!@u�[k�Q�n_N�9��6����^����0���Jit��Cͣ|+G�k��`63�҈V�]���n*X�Q�}�+�|7o���	�xFqž~ּ��?����>�y�E��ܗq�|p�uEd�����,���`�.�'�h�[G�j�l��%�+�_�t�	޼w8�%��MR��c
��@99-����q/i���F�r��@������~[�+"�m��8���_����Q�8j�@w}�a���<Ѡ��Dڹ�s��2��{;����j4������q>����]Vb%��4(�����{Y ���1�����ٶX�!�q��������@v�ƞ�+��{򿑲��Tֲ���x�Z�Q���l��)�PP����������+c��tE+h��J�L�K��EOY-^��>M� 0���N.��x�:n��q�)d��?�r�wJ�%�OpnY���}��V��O���\4��[�5p��#*a��b��W�>�e���%2{*�q�&��Mw��\y>��hc�o�3������q�oKL��ďa�x��k���4��J"��|F�Y{��J�'��1��q��C��<���l&ޞm|JN�_�]2ު��F.�J�|(��Oa�~	x�~�\aѲB�ۀ;y������D��1I�02��*jN̏ȼ��n�AR$Va�P�<�l֥�M���8��'�I�/nhv*%��O1N���}W�>use��a�bϨ�-�7�?5=fW��H����f	T�\�[�h#�{�É�0-�peD��	�
܏Z;���}�~�E>�9i�x���t��@AN�!3����[�0;�GG���	8��^i5�t�w�"��'3�M���=�H$
P�/Ry�����\0}��+=�D��|����p_KIl���A�q���UD�	�2��Ja����LU���>�A�����a��ݿ�@�ޟ5�$�<	���Ql*B���o�����^-V�.��� z����� �q>}K%�lj:�	��(�������ΑB��TG����#�0~��$�|6���@�A�Ȳ��ݐJ䊌��8Ms�i?q�4!J�S�����N���%r�!"o�+N2 j~�.�f�Mf�A�c�pT����n
���� ݮ7����a��b����'�� Z���y�}0���?@��S��z1�ƥ�ɪ}U� ��Y�~Esc4R����7����Ģ�e�����ţ����͎d#g�GΧ���E:v����v뉊�.�v��[C��L�6"*R�r|��,b�@b�4����q�M��Ti���)��xu�Fb`s;��(�<�,��B���4���*|$��?-�\ݎ��n�vϯ.n������A��`o�ȿ��ED0�r�7���C���'��uX�Е:5z�|~��|m(���#YP�`�F��s'���~��nN�3��{��
�YA��]�nR\���p����Ҽ��yS���3~C�Q�\U*��R|���8��C��E'�jB�sk�����"�oL�ZÊn"��!�������V8�&;"PPaj��`�\�	���̶ޚ�Ғ �&�A�ZT�х�;��'V1�����`�⌟�M3��5�6�{6FW7^�cq��"�P��A��)n���f#�E�/7�yPš2�)����7
Ո�6�C-�����BI�&�B�Z�t{��;p7~�W}m ��\��Hz������΋�h�9��[F��}, f.����5N��C'A�`*|���ua]��:�7��Ɏ[,�8������u9�D>�xg=�,��ݣ��9��,w��^>mSm���^���)����$�]�]��R;���V��a,y�b9U��֣���9`ٞw�x�65�-�C������7Ҥ��0EC�;؇���ܑ��g������Z.�x�=Y}FO]czA��ې@�/�4������T@(��sf~y&,�C����J�MR�l?����*t��3�*�蹕ݹabCj�Zlpn1t��W-��tU��-z
E��¿/�k�lժ cy��N�oѐ�ZUC@���2��_ԃ��t��6�����z8Y*z�4([�� ��A�L�7�g���4`ȫ,�O`�C�(�jq��*����18�sYC��{FP#�`�z��#;8c�ˮ'�0��2��Y�l�I�����/$ex����.�\&�F�0o�����m0�0�{(d�T����8j�e�E�/�'���\.r������2.,� ����#�j��0��r�ё���Yv�,�"*�T a1*
�*jߊ�GH���2~`� �|Z�!4b%&Pn=?t���9��1��d�ydc�sS��m�͊��� E�bf᫢N�58�i)�6�鮋�:*�|�������}�)Fe�c�_$��ýc�9��|U��J�I�$��uꤋ]��ꪹǷ�|����,
{��(t�;+Uck&J'��� Gl6�)=�y]���.F�d�]6S;sQ�#J�u�i`���}N�fޯ̪:^�c�4#��BdVqiX�`�w��^�R��_U�F��rR��H�]�YM����:R2��ӿW��c�Vՙ0���-/rv���%��1�ir�!.P�\Y��r!tK&�i$��ک$%6K�Xb ��&�I�Fg��1oF�ewv-7)����g{+u�~;�ۼxҼ4��Pp=��Ф�q2�qg��Å���Oe�ZbG��|�R��)��(��1�WXԟ����!� �		�����*ׁ��,H�t�Է�j�o����fs�i��R�X�DFZ~5J�t{5M���H��AŜ�\l��KМr.�8/�"5h���5o�B�,XN�{k��Zb�R�O���AO���׽�j�g�f�z;�ø�M��U�����W>��.�a����f}����g�B� ���1�2UA��]Jm����|9f��`I����Vs�;��pY��/��l���ekM^����z\��[���:���F
bg��(���+�6�)4W���`אַ(6Y�OF���UOT#�62;N5Z��4g��WC��Io�wy06��^% �y�����+75��=ʒY@A�����ڷ!B3�,yxt_e
��X`��$إHvG�m�Ck��޶�����'��h�����N��I�49�Tvu�m�Lx�?�IG�v�;|ڴ���V��ۃ'3|s߀��s�!��9��I��x��>HO��0�u����O��&A�c�Y�����f2О��']t���BlBed�}h�$w7v�r�)�iR����!�r�f��������� �
R�4�����/Ա�h�P-�?��c�:��ҽ��� �c��i~ю(�E�V	\˸���Q!�u�� K�����o�G��w�X(+۵i�據/��)׸B�_��"�(�Y���;B�/���܏�jHOԳ{��+	$Gl�F�W{a.Q]+��и?x@��*�q���	�΅�D�������0X&XB! ���u!��;D(�g��V�>a�@x�Ll��,{w��Jd~X��p1vC�Hn�\��oM<��bJe7a?��s2�f���rْ�J��m����53M��5-�_\^`x"��!�6�"V%�H
~[8Iy^�
4g\��k��N��Bm���l�.�&l�S`{��W�n��*ѓ��	����iԗ�ME�<��ߖ}b_��M�H�NT~`����lK=�$�JMC�C���'I�[F��$��Y�����ۭKs�+е}b��X=u��k�F�J8��߆Z��Ч���@˩��M��o'���3��.&�t�г��k%!��C��r�(2k��>��C`�q����՚�T�|���M�i��COEM!d�G/#��1�,��E�8.�[��:��6�qU~�9����b�+Ɋk3�vh*�B���6*|m�m�;g��&�#���������1W�Q+$�]{Z9n�e�V�\���S�Ao�dɬ�D�I��t��;f����%fD���5&(�	Q��!��9Zs����cZ��@��S�EA{���|X0��	E}s��R��c�U���.Bo�0����1�3����W.�'����<x��?�͛�5���81�*��t���dT��x�x��\6�}t���ݰ�'?�f<q��$���
Ɂ�	�ҧ��w�,����gt/��OB�ݥ���v�?6���u�N��!G~�N�_�κ8����C���>���GA����a*�(�o�鲆m�D>��A�3[���m��q�D;=3��9�����n�0�>�l����x��y�1ɫ�ZYN�ѥzǅ gK��~z��ý+�|"�,x��5�T�-�ض�ހ��C�A��Tk
�c��3Z�T���O  ��wޔ:�w��QNq��%��z�����u�-��)�
&����l�&�ڎ��kuʵ0�H�/~TS0*��Ƨ;�jO^/>�����P;"�{i}�1�HD��
���$���M5�.�-B�:��W����}�@��h�G�F�׺�9&�֧ ��Fѣ	��a�V��*:\�f�H�]��"�@�  4Z#ǰ$������ɇv�!$l��zt��5�E<o�yX8�XeG�{|r��ʖO���j����0��A�be��u��5?y�4�ܙ���σ�^J���5U>�@LC�9�h�0u���N�m�涠��5U&�=��lJ�E�{�ɓ�e�Q�j*��oأ�I�+h��3hh�G�*'|�����_͛��a�������nU��w:K�G]�u�������V_Z|y*޻���/�O��w����<�u�Io��N�-���6gN�r�zN��~x''tct05�X�-�Z�R	�K��>bs��5�!*�IR/վUd��m۫G�W�Zw�� իhf��V��S���ĉ��NҾ�\�n�N�t,�s���V����֬߰n�i�h�%���IS�R(It���Õ�#a��Gn�Ɇ�J���a����H!�aS��fC���%�<:#����E��._]����G�����Z�l.�z��	�RB�B��{|�&?��[��`HT���,�cS��|�9��̜X)`�w��4��{T�2�2��Y�×��Y��!Wt���_C(�c��(��/E��:(�:�~�j�f�s��z��ˌS5軔1��6P�:�9!~8.t�����d:���^���.��19��2EU�g�G 0Ԣp�a�ɝ�|��\�AQ��g�<��\?.3���3�Da������v���,�=l����!�r��?�/`.W!��-��Js�ce�w�r27lBc7`�_�"�-���q�U��.?�w#����D��qA�Jٯ��Y3�����π�����a�I苮�^;7���!Z*�N��P �	A�${�
Kl@p�,پ��5��ދm�ּ���+��T�ay9�i��c02�@cf���Iv����	A\e�z �q/~��d[M��'�v'6���៞I
��r�hU�Q$��2s4lN���������MI~�5�IxE]m��{�d�ְ����MjF��	�ݱL+#����PW.Q��k�-��m䠁"��n�B=�a�@hH��]2�	�C��Y�F�V��K�����'I̓ޔ��6�y�P1
���IA��bo��A�V$9���n~�+�C'���Q��3�+��H�!�.��3d�$Qo�� ۚE~wUT*�I�-%��˄#Au'�ޛ^�B��C���ڜ` Md�^J�)Se�8��g:Zӭ�6�|�$D��)�*/�H9��k�.��ui\kc.a��$Rd]�iRP�TO��AP�_�Y�x򛘙��µ-�rwR��3�$V��7��?��PE�[�`]O�&�TW�3�=�_��fu����[I_�[���;M����9P	�c�p�0[m	9�'�9����*u�ԝ<	��>[i�xk��	�:��.��4|C���.�Q��]�f�|�����j8O�^����	d�8�rvu���
:e+l_�`�pr,��=3R%�-;R}��'7ZH�]S��K��ֵ3�d~"	��'->�v����ү:��3s*��߹��`mح�o�¨�2�=��!���4��N��M�m�/����=�6}iǶՀ:J�E������� �Y�3u}^�ȗ|��s��˸@�v�����J�2K�A&(��p ��Kֱ�<e�4��7@��,+���4�nB�HZoY���ݛ�߹��|8Q��ĵ`h���3�f��',	6y=���]��m5]�5�:��:{6�S;�AX֙MJ�L���V:�a^��tW�ƟB�X˒y�:楎E3h�=���z�!�w�w� �(2�i��g��.aW��Ř��
�Wk�N"�݀�W�G��E>�&<�o@'�: Eu��J��8Q"����|fw�|���^+3�<�4�009wik�}��I
��ͳۢ�L�������Lң���X�oDF��=8w��%�$�{܌�G��K�l���	I�s��{�1c#�)%���!GHf�WL���6 �I䪊5"����a����y2M��!��.SK�\dD���[��ԕ8��_"��7�HV��)"���Z�m$4��4~|���n�1�F�-ƆH7���#ć�?pB��ݵ��_+��ڒ��B֙p;/��w�(�t;W�q?�,
LP��(����O�ly�0��@}��NU4%�_�{p'E��-uV�x��䬁r+����(MZ�	�>�\�@�����ܓ3a�(�+�Oиѹ$�k���N�yG��p��_�/���ȶ0Ϻ�ar��
��k4�;pq�T�K���s�N��pD5r� b�������V�����R{��2v�	kpS��`�\��E���]����V����t��\��tU���z($Bm�A���DY{�#S|����X�;:��k��D��$�iӴ-Ȧ��ɾ̃�vDd�}�F�ֺ�5�=�9��b��l��^8C�uTLbV�-}f
P3��^2��*r�C������qfG�H��z+���#S��h&���O�䅌o����y�XieH���2�{���1U�\U25�L�+'�>⦡Yu��*^��;���s�C� �U�i�6����s^;Z;���������>� ���Dy�?�D�Q{g�У�A��H��/�}�
V�&L`�����7�����ߚ
�}�#m�H���w�ZN��4�:����u�&!��Ε\P��_P���>�0J����. g�wm+yW��99��/
��'B�9Sp�����z�S����y�x{=�B��m������>�5�`���
����1�)_���j�������FNb듽��T���J�Mm�|����1�A#T��8��&�g��Vh�eU��M ��A?�(�2�b ��,M1���i�Yr��A�*�#b�����BI*�S1^�O�~����|�1���{�����e���Rj���"���=�(��"���K��u��ڹo3����*�"%\&a������vR����G�y�y��ϑ����k��#ܔ�8�7�d9p�s�;�t��&���~&��A�Xn¾���`����s(�jx��'��B�m����y�ҏ5W�j[n�FبY21��	�5��s��Z�BŮ}I =��Ϥ�~�&s!Ok��y�|���o������C
�n�l���֝�����&R#��6�RkK7�S-��� ���,�H,�-���2�ǧeO��d�1#���9�>�Wq-f�E9oli&-��61�}�p~��as��� ����v�����%�ʶ�M����]?���-�H�HF��0��LNn�ޝf$���g�4�9W��v�y�Z�����]�+���+ʑR���N�Wԋ��G�)H�K�]��{G)a0�W~.r0�v�nYo��	��-�Ҫ]��uGw	�½�ߋ=[Mù�0=L�y��%&u��Ÿ�'y �C�� Z��ݔ�O��i=��'_����A��ܨ�k�},���vm�}�M�:��j���_ec�#�F�Q蒁�HXD-��V4:c8Ċ�R�d!2g�	�z���윞��������)�$�����|���L���-P���C(�P6�X��V�^��:��M)`)�U>#w��EYȢ�T�m���ʎ���l��N�滒�IԨM��HgZ�@�o��8�5�&�ܤ?[&z��J���Pr������ǁ1�����喼�VM�yr���z�'�{+���y��e�"]wMNM�*� ����n���7��)+5Y#�TѪ�h6^�02�8�`�<�\x�˫�0?40N�����]/G�/�D��AЧg"�AA��IE=�	x8���&����@+Y�>5i$Jw\U�2���Q�o흛25�V�"�l&�"*���#{�c@�@\sA�mt�hMٜl�f��.�l�ѴX,�a�N
�`j@�"Q�*�x�,��m��s����~�`8��rw��P뼓��o�j�\�jY%f?�����e��`��wd�(��Ǻ�t����M��X5��c� 8��`�(V  ���m�}�.8��(2�{��7�fQ�PZ�v/�|-C��#�8�2��~���+���f�Og$��O����	�{���6
�-kĒ�p�2SK�"ʬ�lZ��H��9&R��&�� �\�O��e߭j��'7�DǴ���fo�|o�����B)nt��ƾ4A��*�*�Q�>���kk�C����[�d�Բ�Z񊋡�>D���{�Okc=P���z��s��� �/H��)I:z�ؿQ%B 1��9�k��@���<���SKEl����2M���N��i�z���7�/-�X=����c<���OT�-\$�=�c�6�l�0����w�� ;���Sm-�{�M��\��t�i4�Km]���k���nQX�eY<19�����pI����������c�[[�çS�ƒbVM,��՝\��;���{m0^w�:4Gy웝G��<|eu�F_�������J��HZV�V�i{�SJ`=�c20]��o+��l�66tm�>����[͢K>f��cnC�#g�Ɩy�"��2��wa{�����*�95~�wm��7 �3ws�Ms��>��R����]}-k!���
��B(��ts�Q����3�Q97�p����6>�HoFv��� c����� �xhR�_Y�^r�U�&�Ew:������i�,���i���8I�єE�����������Lw�_L
�ЮŜZ_:�
�����-�X� ����,��I7�Oq�:��L[P��憝�i|YF�}g��@�vo#܅�x�p��m:7)�ᠩ[^��F�f�W1�e^���P�~�}X�L�.!��j�m��q�f
MQ��	&X�Q�7��ft1-[��6�p�X��(A��y3h�kR���z��8�x2B��W��=���bހ8����^�g�)�r����b�j�Q�}�-p� �x6�
�jB�)�(=Vs	����%�r��4��g��M��{a.,�Wqcp	�)�>��<ĵ9q�W�w~gJO�#��n\�����H%�� c�Q�:��9�'h�̒!'�{�kJ�����X�����zBT�_aްb<�c���g�*���\Y��{5�C��Fy�
���?n�Vǀ δ,3Ćd-���1���jcy���/�4�����#���9A�s�HP��3�ͫ ��ٹ���%�݉f����~��a�)I6���/z�&��n�
'�<#�N翯��Ī����+����V	�/�>�"7���BjL����D�*]ɹ��"A�Ź+��F~��H�4�-T��Nv����R5x��k�.MtM����p��w}�B�����|�;���c�Ê�aE�5&|h��-��M��8�`!X<pG�q�,Ͳ����U%i��Ն���%�5 [9q���	f3ğ���JcS�ş����P$��6 j���ۭN����~��?��E�˂4�ς��|��:�.'Z�0:�N�ih�Y�ơ*^���8ĦG��s�{�<q
�j#@�"�|���h���tH�(�Jk�a������W)>�`E������AQQ_�8��c�k���v�1��4:wK��?ǹd��Co�:,� ۑ9p��~F�*A�:`�=���|1-��� �7��/�#<-�m��+D�t4�������[�{���1����k�G��`��%)��L�p��!���x�?g���4Z��k���f��9t]��+��E�Nv��$�K:��&&�N�S�
��Le'��x'!��	&>�-D�.���Z��q)g�]P����Ss����� �E�5~�������4��_(�x�RH�JjD�*�,!{koy�6�tW.����7i(Vg6�ռ۵�KWŖ��+C����Zv'�$�A�ܡ9z ��Mgj���4�B���� �_��-P�����"|��l� �+�+��V�w�G&�-:��L=ؼŤ\weC��xӣ�Ͷ
�ױy*cs�M�D�8�;�YV���6��'��������&(Æ;1�>sB:U��7�:�ޮ�3}�E�þ�K����"�w��f��N"�ᒹ7\2������;<�B1����XJ��Ax�׏G���Y	��E����{����9����f�7�6���	ÿ�@Y;�������k1e��S��L�j���>ѧ}�����Q��x�,N	���k�ۨwR�犖��o��o�$eE ��cƥ�q�Q�By�_���{�qt N�ձ������;~�'�Q�j��,� ��op�D������2�K�%��7%|RJ	w��4��k�4%@L�-W�?��� o�y"!�s��!M��	�>���V�MT3����U�V�	��)��O��*��Qo���ͭ�[޲�*�q�w�'�g�[�H.Dw�n�	�$�@u�ndzJ���o�o�l�n�A���+h`M���Es,��C�tqN�:)�M�M����Jx�R��?ʬ�I���3�"t9�cj�a�$�:�Q�Uox�C z�V�N�.C<�5g,?�֝�f�W����(��΃ m.P���N�D�J��l�$}�W���i�X> ���'�y �`�١��r�o���-g�N�����&9��d���[gy=j�������g)R��Z�t���3���'�g� ���C�ĀLT�3^k�4�+���������p��c~_��H
鼎���r�"�3�?_�?}�h�K�^e�rz<X�����/<MC� �:7j���)��a����j��W6��Ō���R��?ƫ�Z*�[��E���V��Հ��J-I���f�4�{�$㶺ֈl<��Vӧ��΄}��+����&Μ�	�|3��������mA�K��ځr��᳗]<Ƞ�������7�Jy��ylaVUZ<�}�wK�;]/�l�j�:i~��eI?�Ȳ�Z��C���������A����| )����j�D�6�U���ؕY\~�&�{�p���L�H�[$���1v3ꢶ.>�s��S��j65(xEXqD��<���6`O��Ңk��q[ȑ��$v*�/�������9Sw�+�Q���N�8Fz�MC$�gv�9U,؜��;e�T��G��4��_��N7BBaM'��-�UsG����H Zh��L����^����t�H��[]w��i@t-�$D�g���-����@�+�vϙ��	2Ko�1p��� �p~��9��5}]Y׈��ʱ+B׺i�f��yt���i��2X�S��%F�f���àD��CN�_$�B�"4�A ��X���.Pٟ����Z-BXY�曄5֣����+ݚp�v��]�i׿q���X���K@��"�F��*/���Ȗ��Wt<�s�3ghP�L��
)AM��㘌16GL��U�D��p�e�|����c�=�)]�E����Wyh�9����n���U�������([Q��3U���&�ؐA�7܆��{����e5���gp�[���{�-��,�(�Bݞ���=[�����'ǡ~�Ǧ��w����߂����h.�Ka�D���c���c��c�F��\PA冬���I���I��H�>�G��	;�ڞ
F�rk�Y}?��&�܏w�VS�7o�G������'RP�s�T��� ���I��暗+R�b[���p�+=
h�'I�OOy��n#�,zH�ʻUdQ��/Nu�TNk��c�=x*P �v� 9p�:�f�v���݇`X�g�y�U��vO��B�
�U��1y�A������d���!��;o(���BĎ�M����L�f7����N����mx/E�Y)���t,��/y]3��#/�c�s�ӱ��g�޸���)J��m���!�7��n�S^���t/wv���I(�Hekµ0�W�F�cCv?��7��"�z���`KzF�Z�#�4������W;�^���H��'�M���za�u���C!���ⷸ�ܠx��,��%��5ņ���o��T�"s��coP�g�t��>	��$���	A�G�k�F��,�*�?�9]��G���s<�d�mb������l�RV��T)�z38fD��aD���ܺ��'DŇ
��-L~�{F�%���~r(�$7�����l�6�3����١��d��ڌ�ol��v������\�ЀD�j_�xM�Kt���n�*"2�i��/���ˌ�C:�]%پ�ԗ��z�dS��t���xv�Qin�����z��e,f����)�d��߯f�������~�]nh�dW~��am�`QIabȑN�_Jg+�V���H��(IԪ�W��@�\�k����qg��]�=��U��j���:�OM0M|�'
�҈R�[۷��[ʟ#�X�]�Л���^pM� P����fSf��c���Ԫ�/B t�h8Zc܏�r�L�����Ug��Gc�Q�^'~<�#ϒl.�y��	�4� ��9�0:v�¾z�9���*�0�~-W�f�B�tZ��.Uwe�����2�(:����=0��C;9�yQ���w��y���*��AA�1��`uo��u�V��!:"4Zw7��F]p���1��e[w�Nc�J��I�P�\�N����ClX�}����.-5>�4�R�
~����6O�R;�'�N����Vh�I��*�aiXe�-���Gy^r.g�O��:���j�J�Z<�Y&���45>NW�$ቇkD��n��+- ©�IS�n�by�ϣ��2��$��9Ƅ?�]�s�6&�L��E��gcooδ�;B�����R��t�MRT�����\�眉[fͰ3;(b���%�W�(�Px��+���x�`
��������q�2[������h��I�]r�57%������Z6��|$�'��n�I�(���=J���L��s�HĤ�����
չ3�S��6%_*T����K�5��]Q�䊫�Ko�:�{b(oQ�ϋ�r����o�O��C���<�-����`�Fj��Ia���s��%9\WE��d���߲���v�}�؛�\-!���_�+�37n��kJ�1:K���~	��?@!qQ}��+69�<��ΐ\y�P��R�pq{����\���w��Y���1/j����_S<����Ӭ��}�	�y�q̢�<�T�"&�	B~���#�`�J��gE�� bwQ�eR�������w��=K������ִ�����\E,7L
ƃUn: q���a��j��h��(�;������N��@m�DJ®���{[0�pfq�8e���φ��;Y���XF�Gp�)�g�.-���`�@��*��b�"���n�Jnܕ��X~Sa���쿑F�螨��lv/��������� �7����Ft��4ح��ݺ�][�³ݫfU@	��p<
��:��&�0��2֡�W3�F�0��o��V-���o�IN�ж�JRI��:�9�6�ܣ���.�R��!2kAn�`�Pkϐ3�c��;���͙���l��GBD/���!(�x�/_��vZ��
��d-pW�d�sO���&�������z!Bn�[Dr�;���a�B��w���ߞ�C���;���-+����pS@7�G(��>8�R�Y�a����e�cHJ�X1��kb! ��$^A��-�����;��U'PW֜��4� �؉�7��&�U��*�'A��'9��Tﲨ�8Լ��P��y}��x��7R���KМ����ѣ����%b�+ӝS�5;���k���КW��Ѣx�E���\&seݷ�ɰ��=�l �[�� 4�ل���orFg�5ԷJF����Ҧ~4n�7+i� G��0�&b.��BX!��?J)�y�wuu���HX�qw6o�^�ٸs��fU���:-K�=���)��%�u�n7�D��)0�� /ڲ{�̀`���|���sJ��^s��-n�����E �j�sEF�Ĭ��
��k�e�~�y�am�_��u#b�.;�jW����>JZe[�ʠ�G�i`�Gd�م0N�5ADx�^��8:�8��J����4<	�F�ݱX������_�3�����朌W��<��S�[�&��XHu���B2�Ĝ�����Vh���ߌj���v������*+�^��	�8ԑbx��i�Yh��O������<^f&>}�;}f���4(띬e<�צ�)�ظ�'�E�*��)"X�
�0*z��m|��q��� ,�*LT'5���]\J���`7}�]��O$V�
w�	X V����K�pD�K��I��TW���Ķ�KH�#�.���	�:�q��#�5�O��q� H�&��t����tР'"�@;el��:1�7�j��W�6��En(C�J۬���5�'���2	�f�C>|K���>3��)ۇ����{��p6H�j�9Im�QC��̥�YK�Я{~�ӭ�9K��?�g�$�\}ܾ!ڀ�f�M������f�l����_��ol�;�j*/si��r&�n�����n�j��Y�){65��?�����P����ZO���[1�ڸ�w����qؕU�FĠ��f&)$�U|�x��Ow�s�Ҋ�@+sJU�}��5#�^D���HqJ�H3,�kPv�������ÄO3L���]OL�8Qu�xԯ�
:��������o�G3솦bf��$L����d�\3�kK��۞v{#�;6O)T��&�����ŏi�qlnR�����Ā_�g~ڪJ���A%�h�Ȳ=y�:���$P>��H�"@e��7�}�y���7��7�g�����s�����c;!;�P;����+�N�훂�^���Y���u��J1r_���2��x�w�����K����vN%f��n�W<q�˽d��a#9�+P�XzN�$��`:M�c��޸4�X���D�Ys����L�����w�Y*������N5m~x�WBK/���O᭱����kxʨ�r4�Ҙj�!@<�H*���+ί���ёc�ԝzP��d�)�>����4d��Nt�$�nЙcs�pT�R��5�O��Q+��c�@�3,�=�2:3a��{�����*f&R����(��>�%�qS��x��H��Q��x��E��r�"�\05ӧ7�V��� �����|M_o�����Љ�ȥ
7�
�� 18r9>�S�n�x�ܲ���Lzsp9B��r�~@M��������ʛP ����&s��Y��j󗢧9�h�u�ԎEMM��ǌ��L:4v溓s�^����\M���T�ȀA0eS�"�e�"�+�-W�f*!����&���d_bG&胅�J-�1�o�

�k��[ac,4n�˩�v-���3�Y�Z�3�ޥ��T2�)��<�� \��-������٪�[�/��԰y"�2�攻x w��/���uZ�Q8�pڃw���!S���:��E���}����ߏ�ѵN<�&f���������{��#��&��br�F]�fh1f��,7�_�鋖��mRAh1!�%8Lv�୥�|�9�$N��snV��]62�&�Yv�!�Ɩ�$ĺ[��w�����ϳ����~��Y������8Ο�C;L�+��9��R��HY��-ɴu�����ߤɝ�bO�:���Oj������Z���ʧ�w����l?��xp�鄈t��� "2<�$T��1M�6����I7�	��P�95b���Ez����U�bm��7���6��OV�Tx�I������$|��rƖ�z�q�i���V^gq�7�W�1��s^ee\�O��|���d`C��Z�Ó['��ς�
 G���E�`�����p
��Íɢ�^K�'���),f���=�a��N����ۤ�8��+�Jg�-�܎��LP-;���;�	?am�=x�*�;ER��c
�U����)�r��	�$���!�x�Fr�Y�p�@y�иVQz�o���?�}s�ffR� ��M��Y�pr��ø�x7�e�R�s���5�(@7����5U�4Lz~K5��`�BZ&,� P��I��K�{�͡FS��LCK5mL��P1 P�°?�uT�`Ҵ��	7�#v�T֘#`�+�F)��T�XJ�f����*"��r
R8�Z����K�,����b�����0�w}M��}�0�X���3��:���n�1bUn�����8;�)�l<��RC!�ĩ$���g!�w ����8�b(��%�_+^���h}�*.#pY��U��a����M�L�������������V'y3Tj�o��aJH�qc��n��2��icjK���>��B=E�X�uƄ�7�4q�������Yvu�B���奶L��)�[���Gbhn��i;��Ǩh��P����`>!t&vU�0��қ >�}Y�MB��:��2zWA�.	����!�uP�Be�vTCKN�N"l�^X��h�;A@渙o[XgdZS1��O3�G�N:D^/}�/R5b�������N0��y@m�*��궯������*�A��V!8�����(��ԪftYl �%��eK�+rw�G�"��|�٦ʡ�b�ד] וp��<~���Ծ=��e��/�6��{I՛��'FtV�hy�)�#�vVo��i������G�Ԕ��B�~�8�d��=/�G�G��̘8w�Z�6�4�;���ǣo��3YG�{G��l��!�^���/kެ������	�_i�n	:P���Ij:w�E�ʨ�#�Re�,U�Q���� F������!/��mU�/|Д-���0k���>��vC������p2�01�\�����]�>7z�;�*��B�i�ͺ^�:H��|h��a�zueى�;Gyx������j�p>�!���W����P몷�������rs��i]�
=������:�⾲���A5	��+r`Zd����ʹ�O��ſ��=Ir���i���Nn��@�{�v㔐��Q!�|r�N	R����F�������~���gQ�A���q�`�G�O�Xk��B׻�laM55UCd�6Ar��od=6��7[}����i��	`̛线}jvYK�L�z��;�i��<������ηt�B�Be���[��wh^��'�q ����;;^��,}J����gx�H��ZK� 6�J�j��x��V���v���gŧbH���^�Pёȕ;�Olm�N�)[�gT��8|�ךI��H����6�e"�B@�f ���_�����V����6G�tݝvd����&<=qy5���8Ӝ�:!�z�a���Y��J[�&6��m�m)���#�-$�y�['߇�NO��D'��WXM�ƅ�kO�i�R-/L5A�T��gSZJ8*�z�x�_HƱ�M/��ΰg�w���@J�`ʵ�8�m�)?�]tI�'��a'�u]O8;|>��઩6�  ɗ�<h�׮(���7}/�cR6����~��[v�X	B��:Q�C=��Q�&� ��qWϼ(VԸ���e}����e�~>5`o���M0�)��BJ̗[���2��L���AM��qX�X
��y��0��d`���c�(�pTg�Y�( ͙K;3 �*���P@�
������5J^�)^
L�J�����E���g\ֈ�2�C!/��&��c�_��W�]g{M�l��!r-iM�4�����>�Ov�x^[T�<i��3b��s1(Z�U{��3�ƺj�HCG�}�C�O~�L�`%���l��e�߭��`�`�E�_np=���'�p���ѱ�Ar��wb)��j�� $yg��f�Iɉ�0G�^�����b�|�bپ��䁫��#���u���2�9@�	�e��Z�n�A� 䓾_��gc�I��=v�� 4|�s�\Z�	�~=�765�@�J�g�o{$�d�2	\JV�Z}ǃ|�MX�s�����"�[�<��f�Ù���L.f|_�>`�Zn�7<O)�w�Xh5)�~ϲ���(��� �hHoh�HF���e(b�0cf�ӥ�M�+���Q�p�R�ryJRo��S�<���\#�=�`X(9oy���-iG�0���]�����{�h�����x;Bwl88=�b�ݏ��o��u�y\��o��7��=��˷n*�������V����y�f3�|�0���Y!�wX�r%f
C���l�w��ڨûB�)�S͔�����7�����r��ǩd���$�c����+�@&�(�@h�2���*̥L��/$�>{��	HA.���)��Ox�m4C�k�篔GN� ���������z�Rh>su��^�T{䶳�L_s�%���R��C������B��H�=HN:9_ɿwjR#l(��D�q�:m&%�1Ջӹ�
+�������oQҧ�	��א&N�~�D!��k3J��@�Ý�D�a���/���T*�Q�%1©�i!��d�7k����w�h=1!�S
�g-c�g�9�-p�-�V`Ƥ�����xǾ�c���I	��0'��vo>���S���U��HQ���:ښ�Sp�A�JTU@Z�0���}-=k�5=J��sۣ�3�H�����$�9F+@�A,����TDR���}u��f��9�����Ꮻ�~*%�1���~GCMnTbe�l�n��	��y��@�f�I�(N+�/!$J�5� j���暽դ�n�|6��*�%��#�9���t.�fYs\�I9O{:�ۚ���}�����|3��C
�BL�_�&����v�cs�3������s�醹�ݼ�Hh����oy���Q��o*�-�8U�"s�Ԧ�d�k��6�2���9p�r�Pl���yq�&�3��R�Ջ��wB�,$A	r����[���q�ilU�@�d���+B� ���,׌[=r�@)�ܙ�2FZ0�,����y����:��9b�u�~�0>��Ev����E�g*ؠ�}�h����H�vP�˵�9 ��e�sP�(,.e�ʃl�ϼʐy�h�X�����H9I���h����ɛK��t	_.s�<
`}z���H�����x|f+K�B`ṍ��t�Rx��N��ڃ�G$��br�1Ԋ�"VK��~[4�X��Z�;>�迵S@���}.�OPv�����@�ZnD�@Z�jQ����p�t��� {f�
��� �&2��R^��A���S���{���p�e�B0��ϰ��\n��\z9�{oYu��kc]ۮ<����%��u�+�Yϳ x��z���[�r��۫�-fKh~��n0�f�6�7��; ����4��o�ږ��ly'Y�6z~fc�1����.U�y����Y~�����-��m`��c�Xu��=x`��׏����l���zM�y(�2 ' ��A����z�y8��#�G3��wE�e�����`#=� ?4n�"�B��(�f���yc�?�����}��A�2�u4c�{.�?x��]��pa�U��ð�=*���wk=IE�-��-��wAA��(nF]�(Դq��
(cI>}#�.(]�tK���rQ�J�s���s=�繞S�kn�Տ9�9r��څ�L�l�Iِj�IA�{�v�2��?ԍl#�U�{���# #��e��N��G�	v��W� "��=7֮��B*�d[�����s�v��R!��*����*��$���^��T�^�u'>M,��^�<�I>�*�x왘�K�
������XQ�?-�r��6����bt���9���b��QB�q���>FQC;�P�����վgX��*�/][�!�f|�@A��?Ê�t�`��o�ϭy,�ӁQ+��{Q�a�#ĸ�?�c�8�p#y��_�2?Z"JӮ�y_7TH��}��gr��@�K�[&�	��a��\@E1���w��"q��:3�B�o�DLܲ��|�����.t}\+��8E��o�����(?�Q��AKՙ~S��h�
�w��9vE5����Ϛ�^!Y�s�?:F�q��i���[i��*�_A;	Q�r������*��.�;�$y_���OEa z���,��' f���8bX���-L�췽u�1X���Ah�1����1,�
�c�����^t*%5F�����}-���������~SJתa��K͟�W�B�H��+�#v�xq��׋x: R%��gi�׹�V��읥�NϪ���Cc����������;O[#Ra��Up�[�$�Q��Z���Sb�o��_�G��k�v9M�R��%�\��#�k���hK���i�-'�E�B�������`�&̞px��phWu����"]ڨ�@PyO�~p�*9��~�
��zv�[�=��Ŗ{b�����Ãn	���0��Z��'�X�,Ў���X:�p&�G��t�1S'#wA�8�)wʩ��≡r9+.��� c�U���.as�,tm�7d��:\@�b1��V�5�S�K�w��X�����}]H��9��M��@�Ѓ�:)j�ıj��eB)���b�J�̭��P�����]��׶�e�R�q��g��곾���A�q��9v��>ľ�r�	6F]��p�p��5�Bʪ/������&����vi]�-���n�*�0^	*Q�����m/T������ �Z���t3�>�r� ���L�Y4��oW��������k��Tng)\�n�@=�B��6��n���;�΋lf�>hj6-!�h�:T�+���� �C_��A�ۏ-I)���y������$}�kؘzs�q>���[�"g.�ӳw�{Jpkx5�ȗMIF&r�.`���cw��!U��P�N'Z�F��$����n�M�'�0������e�l�
Χ?�N���BK�44��9�IE�r�g(h�T�ò�C�˅WB�V�ݔ|Wx�8�8C���X����w
�	T�0]Դ��Y��N��>8b���F$��Lgh<���3%��P៷j1�fF$ܩeߋ���~��+��lM�C��(�B��Y�r��\'sd�mǉ:��f���'dX�V�B2�H��𞊠N|����eNpKu6ʶ�r�����,f�mD����p�K��%�/$�sg�/�� F̿��
�ؙ^�2��XY�Cp"�x�O���F�#�\`����>�H�p�7�-^�!�rx�tpe�P�@o�T)4��Y#�a�]���������U֙�w�:u��
2F��Y���
dF7?�p����@F�ʍ��������/8Y�`�|N@��B�(��OQ��aHn�i����~�=���+��b�>@T�fuFҮ���W��d��=v>f�X[u�e���G�!`��XM9CP��v�	��kN���Nq`��U	\��Q��2�3�O�D��Ԣ��q�ߋ�ѥ3��᱙*ҳ��@Ы������W|��`�UK;>��p>ݱ��mm9��NK�Lü�9�2`��B�s+��q��3s����TE���f'j�1�1�gG{rZ����t,�$u�H����pY/N8I�6�z]�c��� :E������nb�B��A%�|�?#0���d=�B�h����T���3[st���d`w��g���kolZ(�7F�h�A �_��i�����ao�mBʮ���j�a£C$U�� �5y�F�_�e6�0��F�NGz��\DB*�����$ǡB�h�u�F�Nd��}N�Ki�q$$VF���e��N0���W@D��ex�MMD��.@Y��2˗å�e�y�p!jZ���ܖ���pK��r�G0�uPl��?�����c��*����A�į�8��z��q�􂼎��(���6u�:8��f�u{B���B�C4ϞK��'��)��b�6�g���o�� ��|_S��� ���P�Ō��A��~%����� �������\їY�m�t^m�̮��)����2�?�7�"�%P	,�G�F� 71�iQ����]ޑ߄]�m�c��0����a��.�ܒ}���#a�K��i�@Q����p��}u�$0���Qu����m5%F���|8�����C�z)|��n�,8��`7�xw��Q]��>�D�W����GO:U�١VH���@u�M>�4��R�-cx=M���ݙMH�b��I$+g�1��l������ Q+��ә?�y���<4	!��z�K����Hz��ə܊�n��+��SbX�����OC���8eP��3<L�I�[���&s���fS��d�?2�����ֳ �d�f���Ӈb,d��esƛt����v��ʕ�qa��W�ul���Q�H*P�~aK>��\�(0@
f*�`ޢ(:�v�/��S;�ॠ�o߄
�Y���oF֬cOHz��.���L�®Ԙ���(�mL��N��M1����v!�9N��UsC}�������p iܗ�B,oS�߿�X����9gZ_oG�p������`�>�pDlM�l�1�h_*���7�A������_�d�,�L��3HG֯b��|X�F���-�c�:���?tA��$ ���}�@1gՀ�0]���5,��Y`7�LB���"ӕ�Щ����<�|X��|Y�І8Gv.��:k���17JW�(M��=Y[b�р�>~�9���Ҫ��R��8�pPte�E�����Ψ7�2���wvZj�\�
t4���tv`�֕��XT�,C���	6�s�>Lsf�l�0��M�T�j�c2r6L���ҔcU��j�2�?��P���� 8��Jk�V�]�)��N-I�����»A�ŧU��EP��i�|�t�l���{U <����QCOek��n1�qi2b�w�d�XN=]�E�~lM�^����!�����|� �u	�d&6hS�i�˜"�Ӓ_�3�tw��.�+�v�0�r7_�o�s��<���x��<�+Æ;fl	N�F�t��R�ğ�u�xw��V*y1|BTx�4��4�е�h�1׊�=��.~������k�Qu{ �Ag,���zs���c�R�ͧ�3����`957K�-�S���-e��C�^�=@v�y{tQ�̘q�M$I��Ě����FK�Կb��E�x=�#Ǥ��h�ֵ=li�	.߳ϕ�M��H��/CAnh�g�1���O����������S����|}z���Wy��j���P*��4�����P��v�d)��eHl�5�`�*��`]{j�K^��\&|�����\�9�9J3J��{կs�_��t���a]�گc���}w0�#���7��g5@F��(�J��6�H�Pwl$����~i�>�~�-��k"�V�q8<Pm�`SEr
�S��T���3e��dʡ�"����0O������WA�(�T���ϻ�,���J�����=��?D>M�9F�//bi?�����i�w�N��Wz����E���-���":Ɋ���7G\�f���Rz�[��(uoHjW8|�sYW��T�Y��>>�|5�/�nH��;�KV�r�2�����!���۬��/h��cUD#����_ރP3\��{� �#x���0I5ў㞛��ՒIHyط �J�(V �q�o4���,H:�����U��rn����N�ӛ"B�g�TaZ�y��Dp�K��-���K����	u�^F�P�z��)������ϋ29Sg�́����Y��<�f�>I|�� �Z�]�	Wݽb<1�['�9Y����rڏɱ2�v�J��h�@�)HI*��څ`@��7&凋,���g�����磰��l4��9��A�
������;~����؋�m�w��B|N�6����c�Id����ro�y)ˇB1��/(6��AU���*�-
�f����.��3L/j�v�-�]Q78�/P��!`�j��g�Io	Խ�����@8C>�E�����.J����V
jdu�)�����ۊo~�D%�0:��%]�_��1B{$kV�5��I	�E-i�z�i��l~���d�����WH��2�,7[�g����w2=�L�vKd�k�g�׸���dI9�82��������^�߄��m+��T�^�B�T���3¹u�QaOwAg�~Jd%�`<.mPR������	c(h����\~fꑞ`��a�xZ��,/�k��|�T)�!�h���s7@�v�@���� �b�V���VIwd��[�r��9���C2�A7y�i*@�]�ٿ����H몲���ܱ�sHm"	�x X��
�i�T�g�\�&K)��J����_\ ���=f���<�d��{���S�ܫ�N�v�+y�������q��~RRS��3ɖ�.|~� \.���^O��i
C�5�i>�!���3tA���ݰCt���W�9z�8b=��+$���O����|�a]�i�v��Z��h��ן�~F�6_Px��g����'�vA��lAB�yc��p��!��;�̇L7g�������`�1#���xv��fK��V���\X����⌓mJ���==���(<E�P�&�O}��=�S5p�"�z8dȒ����Bс��&���`#���a��4��/=Ϯb\B;{�7���ܳk�w�>}��b *G�P��"���V��+���+ȧ�x�am���
jW�Ʊ�	CRP�1aZu5	qE�m�g'��?�<V���8���)3<�齷�2�Z�zc񿔷A�AXUΰ�/f�Y�Ow3�zLB�$f�i��,�<mȄ�;������%������Nܝ�1����t��A+��z��C�sa�7��aS)C��P�U���͈�'3H�hbȉJO_�<��.�~\�#��מ�4Q�
U�3R�Op��G��te���̑��5���3�ح{޳��"3�ոq�Q\���5�}���cE4���=�Z������}�32+L����g��O:��?����zx��ު�J��5�ln��b��%I�'�k�T�{����NHQײZmHn1(�]�"AĘU+�+䙶�9�.�MaЗ�#��gߡ�B�sĪ�l�
M2�ӛϻ4���h��xÂ����o(�t�_69���s'm�}�0l/§��=|�<��ɋ£����� 
���\��KH��I<=�C���G��Nŀ�}��L �����#�f���L� #K����<������C]��Q(��N�_��� (�e��	1�v��E����*���[��>��XĜ��׬d��Z>��� -bЖ�u��=�#;�t�͛�C)�EᲸ��i��ld��(Z��!rZZ�Q��{�s<�<�߯��5)�ڍv�Q����'#��n=w��ӎ�b3��~@��Jq�ۧ/�����J���H�qb�j��%�N!�w'[Cdax[:$8�TPg�qd�ٝ�u���&0{_@�k�!ڋX	S|M��FI�o��n���SWS9�7/��NxԻ�0��Fj�����<��E�'zI.ED`�̫&�3;a C����X��ד�BL�/�4�ԧ��_aЍQ��&g�~����{h��k��eΗ���!�ګ���ͅ��}�,du���O�/�V���#QP~�o�Wo_`�Q52�a(X��W����@�jq�� E��T���e��>eo�� p0�\|�uJ��0o��{"�����<mr'�yοf�^��,=L�G|�l���ex$��遁��~��KҠ��g���з���$�Zs�p�c4s���ZS^޷Q�!T55=�N�))��
��B���=�2}>6��^�Q��~�5�����^�G=H�L��7����K��*��
��|��;t�	R7�n���(	J��ID`�5hE�ԈҘ����-̚�bL����t�+1?��~�u]�K�9�Ú�+���I^M5-����:�oM�BbW;�Z�uL��5��iK#¦�p��~�K�Mp�����0 D�����P��A�� �����(��L��U'������w��i�DJ�`m���ob��@?���B�	�LA9-�\��Ms;�X�
 J�tP�{�@��
�m��n6��C$��O*�����"�����6�ND��ֈ%��@�*L�b�r��S"5�-sC`I��<��C��<3e��Y���g���0��֡Ɇ9�\�%$�Ѻ�
蓢	G�HA~�3����5������	�ɲ�, <E�T}����Ϳi��_�߿���j:T��p�oq��C�#u�W�Ľq�����:9J�Y5�E�p,��n��x`�4>�5��"�v��z�x�+^t��2�eD�v߫MF����vB���j{��hZ+k��\�t	������M�]��t��i��V�-�x����4�h�ۘRm0�J}w���_n�K\7j9I�]�/T�x5�[��f�?�Ңt����lB �c��#���n+a��S��=�����k�&%X&O�P�d�8Ybs9N{Ӡ�#,��������6$ꉦ�V��/KX,�,��pe�"����5���ŭ� mt;U�'�
9�)4�N�x3��RZ�p1���>�q_b2ބ�3��0�0(�;G�B둙,=>^8�1u9�T��q��d�8�-�r�e��䦶�y��V�ߖ"r���F�n0���&��H���<UվUy'�E��C�5�%_E|l��9���0_h\���T���G6B���P�����JY�
=)�o9��^�l5$�������b�����_T[������u�C�蓯�rbY�q�s6j�C�@**��*���L��}�P�*�J~�ž�����~�s{	��u�n�̙Q�$L��5_��w�����c���չ�������jA5�+fN�a(���t;Y�q��-mP)~$ړ��c��S4�<Iڼ|��3����o2����->}R����;������	�xf��ck,�F��N� �y,v������O{�FA�DIȣ{��&�N��3V��Y�����I0��8Ej��F}z;܇�wO7O|�I����xc���tSƨ�7c���cmF?���w�k|D��v��7 C���'��n)���{�謼��{>#^�����y���s�$y>���>�RB�A-v�{`5*쐖�/�G�sU��^)t��V	��[7ĕ�+�9����CV�ޗا��н_n�Jn��`��e�W�D�6��C�U�n�І�,�#��,1IIr������.G"s3�,d��Z�{�+뫵�'�7��G���Z�4a;�k�M3�A*����p��p�y(�Aa������������^G���2h�ۍ��vHp��%W�u}j|Qw�a˞�h6���0�E��WRGX��U����mT�mM7�)y^*y�D���/Wna��GbχOy+*�ʜ�� �+���"i�۾U=��'x�)	ݸ6�g�1��D���6�z��K�R��W�܊M�kq�#�>)d���[��*�͞q�j�N�z��Ʒ6�}����-yɴ�Pus���5�H�d��{C���뒎O����VS�M�4h��-āھ�(^���b<��m����qq��NV��,I��5�Ū�:���\m�|�yc[D�`9<L��,���Br��(e��a�鱞���G�9�ؠ�~�2Fh1F�lMN���_�����஼1W`�^�L��f24
zcs��S�+�<����F��};fR�͠���>�#salS��l���6i�0"!��26�~i)��մ��h���ׇ>��#j�K6q#����%����/��*U�I��{HΏ50����X?����%��	��c)`Έ
�[���K��.Y���w��$��f��/��p��q�$xK&Kpo�<?6n��usQ�([q$b�}��z��	�H��,R� �/�J�7��.���ս��8ξf���{�?K�CPtm�?]����/�T�5�{!Ʋ`�Fy�@b�95a����J/�\5	���������6�w��x�9��KX���3��ͯ�l��Yys lr�d7-u����� fQ���u-F�e�y5���6偳�p�弁Au�g7֗��!����D�l�aB�YlΟ�b����i0~ƚ�y,�
�M�1ܨ����*H������=Z����E�+B�n���M�B�^@�>��F|b?އ��X�A��;����ԗ����8�`62����W�(+���<?R���y��j�А��:�@����Vq�/@=�F'��YYR&��v�=���Q�>/\q�|򣿾�p�!��d�M�L�L�۪\��:!�r�czF�n�'�+��b���ԗQ����a7+_oP/S]ݹ�x����?U��I�"�{�������n),�l{j]�z_�d����A�Ϻ�5�$�nⳳ�(�s��|���P���X�߳{x�R=J��:�24CD�?��3���+�;n�;�L�_�rc�=w�,��l���/C��M!a�E��wƞY�Ln�y�-��'s��vBo������X���x�����VV&/n3tk��{�����-aqX/��=ď�?�ᇵ=9Q�X<b*�kE�J�/�t���� l����~DSӿD��6x�#h.�$5[��Г�=^1�NIL.���h�5���m���z_?��mx8���#`�g��p��Y1�Jl�QQ�-���cc�`_|�^��9�lۼ})Ť�>i?Wl�?Q��Ƀ���8��R`�w.'����c�{��GT�O��Ȩ&\ا)&�!f(���=`�Cd�'��(����B� �76�0�c������ZB!���6E��E���٨([�#�N~��z����"��Na�w����d�⭸`�����'�7�HƄҊ�0����g?�#�|��*��L�;|o��ڨ��
��U6�±�F�u�T��\���K��	�i3�q�ڨb�@�˒�'W�wl���������dJ�4�s�Gcҝ��wn,��<O6�V5�����F�k�{�D��Q����3k�`W(l�׌7s��Z/�1B]�k�����ȂE�#�L�܁P p�����u��c�?D�)��l���{�xz�-��`�-*���}Vm�c�X���vdޒ_��5��Fvao���z]���>���5��`�M��i@	�A�!���L���U�AK	f���83[0��	�����qH"2��K��j���gp�p:�(憧ML�!{M
cm�$q���-����xZO����[�"KX,,?fE�~g`jG�
f�`(��}���)�m/󒁧�>cH��B/q��t=�C(x�J�?M�K�V���OX������7o�^�k_(�2��T���K*��;����RR�k�4
�zTXf4�߹T��>P�9������$�1�a"
�8m�y`�?&]�w���Y��XY�

¥2��G�R�I��A�0��Z]v�T�*�2E�VH�kj�v�l�-.#m~F��l(c�{+�й��O`�A���~#HA{>�N1�HY{�~�;e�J�4�T�tI2�	��/��h��9�d�v�7A վ�A����#n�v��V�Y�W�r
��0 "p�X��'��w�jj٪cL8 ��=�[��h�|�F2��=�!tz����s���ѭ�g%Xu�g���4��i���E���_�;H�^H����9��oz�?�|�
I�#�Md��N�P��X��%��/A3�Z�L1�2 .�4���N��4~�R������g�����RS�gPr�O�%	�������%g��J>��M,�vn�Iƪ>j�2~�����AG�s�
-a�C!jF��oV����8/Totpof��3��#�#kb��<,�.�$ۗD^����\@����_(S�Z����5��m�.���H���]��#!�ؑ��"�S�J�r�
�(UO�?�<��p�':V�B��Ynp��.-��c��}�U�P%�w���O� /�;D\+�3���&p<a�F��$�|�פƿ��:�t9��E�67&��P!j��0x���l3��b��j�-�GerRr۟��znq(��H��B���J�%B��o��F8�e�������` ,?���i���r���h4^[���L[��e�^�߀��M6�9mt_Nq���lf4�?�ΜA��ƫశp��� �̪aއ荙 ���.�I���#p�l6B����0�wXo�X��+�7��=e��3���&�ˈ�7�<J��߱_�����:� 3�ᔽ�'`sWc�e�@��+��L����p̰���p��uB��x=����ҮЫ@$~a��ƃB6%����W��H����Eyy8M|\�c'!û���c�.`��{cᧆ�$i����'��ॉ�p��.��!H�9��,و�v�g
l��{C����qF�����y������]2�I�Lp�>&��e��/� �b��4^�(�lB�[*�|k�ɖ�'����Fʶ�f:�ź+MM����<��3pT��f��H����'��.J[��R�iOծ���W3T-�F�7a>�Om�?��.�@,)&M`ƫ�75h1:�f\a�Y����!��^t�<B���0���2(l.��Y��%�����#��N�V�C�#R�r���l�
 ��B/X��Dܭ�4
�4�#d^���)췆���|��B0.�3�^)�,|LX>�e��է��*�o�&�cS�5Q��q���ޒl��9��ٲw~\�1�󣃥������S�w��xi�9^�f�|,���.,n- "Ѥ��Qc6C����rۻ!�י�W��0Gw�~��'�BT&�%�Æ�Z�6�T� ���#�wIg]tB5��*:��� �֌{.�ã�D)j�f�c��EzϖIF��M ��_�^��X�4J��4�i$T��@��Y3����$�&���z2��[fcU�x���W)�t��#�K�
���BE�f��6�2�*��)%E��4Y�Ε:T�����-�}�]u�Q#����M�����@;�Cj�q\��.�\����;���IEPe���rY��J��X�*`�'R����#��Û'�G�MD_�E�r��$jK��Ч9i��$ko�^ׇѡ����{��H|����;��54�T�M�]���@��ᢑ���nF9/�����/�|w�K�E.J�֒暧_����%GV���^X����j_
�[L�N5��u�H�a����#+=pv�8R�i��OB��UbLj�*-��w�r�����%ݜ��$�� }&�q��-�o13~��鿵����<�P�!�)o<�{��}}��������2�
딪>��|�wL���N%����,8����	<�♚I�qrMc[/D-�z
^��x����B��ⴸ�r�O���.;��,E�i'`P/��O:-�Ɇ�(����診�-k·�viXq�kQ0R�щ��I��]�ᠠ0�@^8�/E�V]τ�������4���{��F�#�I�D�=n@kK:\�����\��1^R!���_q6z���9���|�����j��Br����\H��I5T���؍��QvK,��
]�Xa#T�č�r�\<8�O�D�{�%_;����R}�Fh�Ҳ��?��#�r��͕a�U�ӱ'Ea,�����튮�m�sp���%${'�� �Y �w�Z�I4r<h~S�0��:��w��s�&qX-�_�g�(��|)ޮ�_y��=�i鸌��䠽�b�S��d�2o��Į�VI ^Ƥn�\)6��~���]�YO�&��&���p;h�
�d�$���K������.���k/�5xO�����{ ����H���yd��g��z%!D��\J�!7e��7�W:Z��2f�+2S���	�} ڡ�����|��5D�_�� �y1	���/
�4� n���70@�s?X��w�#�v/Q��_m�F8��{��Ӊ�.������҉w�����f-�)a��X�f������1[�"���u�Z�%�Zx��g��}��$xVA�����=��s�fD�:a̒���tZ��N��pyly��?W�O4r�\w�H���/ٯA�K�(�O��j%3�'	�8n��Ľh�+# �G�H�G���C�O�>y��,2�����M������{Q���>v/Z����~���:�Z�|�؛� ۢ		�!�~g��QLA��,V'{�hT�������teQ�#���C7�$ N]�z�N��Z�j`a��0RJ���mz̝�.F��k����B��}}��+���9
��3�����q�O!�Ku���>�VaR)���K���yk�õ%�ni�����j�-����Z�5"�W��l���+�?�ր����fL-���1-��b�QŞ����� �
�������к��F� v�Oz�'fi�C��u�ۏ�$N��?6�XW�]{g��7-��c�pP�Ѹq�/���t�
��#F��^�28���y$����Yw����;Ӂg����s� &j���i�r��S�B=�w��-?N��b�(M�ٕ-� �;�9����57��G�ˢ<�g��@�]U�����Lr����I]�����;N�j�{��l����ʥ�����)��7���q<J᭿��k�>c��*�2��⢧?��������Ю�9/f,�ώ�N?�5�q�ITc���ן�)@|�%���ك�@;Ն�k�a$����������)ոl)㮎⳥����MX^:3E�[{D�Cq|��NԐ�	�!s��hM��<���~�J����fB����-��=�Qp|R/�WcH;�o�[��cSbi,~��n����dT��D�D=��*�,�at}T��B*�^�.�r�B����7%9�%B�\��2_����P���\ -����ͱN�4")���<?G���7j�L����^�]���oZKⒽ>�9�=��+��5��K |�^-�1�\���I+�gt^���=Fy�9"�z�F{I��M�Xve���+'��A-x�p�����bF6�y;�!�F:HP�NTP6�r��bs��u��z��\���7C�!Q����t�4^8ͅ��	,>&���g�'i57�t=�
2hQ�9��a���wH�z,����lΑ�,�&�����|���� V���GY:cn��ֶٹ�Ω�&zuG�4[`$`���j�4N�EEa붗�iD����HıCJ6���¯YE��\��m�)�<���"4��b���6So�s��>��h;�V3յ&|9=jɴ^��)����#<B-�}�_�J`����W�׹�����&`��)	J>�8��La���/\������O\�<�B�?W�5�J��q�?e�;��������=j�1[�>���9�8!�a���+���G�]O��z11�tR�w��ۢ��`*�0����ߔ{<�P��H�p��&8��v�ß�������$��v݇m���,?G���A`�|��]o����쌄�m���Ҫ���XE險�c�g�ˠǅR�k�(�_v]ړ�R�R�G����I�U2��7��0�dHĮ��ϔ��BԔ��'��������6�o�:�H��f�3_6��G�bCĿ�a�������$Y���B�ڱĘ)~AZ�ɞ��h1A�j =�G��E_��t����{Z�Ӭ�][c_�@U���GϱIʗM2�m�L���ks�p D�������s�sWb^Ƒ^���y�? �<�m#C��y<���ul ��׶�����ʫ�^�~�U���deX=��1�hsp�ە�Щ'��Z�/YL��J�[�HT�F4��H�fq�+쾋0tJއ�"ZΘ�,�����F,�68�t_y�C�(f�ț�б������I@#M~�8������Ƿ*aw�m{�n�ԕ�	�UXN��2*���'��2��x���J�,�kŹ���`�[v�T�4�GE?�mj�ᾆl��8��ZTg�֕�<���V����%L�s)+�H�r�8X���"�y�+^�7�� ?�GǸ�?���˸���poS4z#q�g���8��ψp�����4It�'���GJ�:O'f	��rX�4�ga��-��LO�xj�w2��t��sh~���x�矖U_�ܥ�C�ǩ��v�*�p���,���x�M������v�UӐ�W@N�z�L��.;?�!M�I��#�ڰ�"�ko�J�R�B
��QPq&�n͙��{"Z�6d�w���H����UV�Q~��8ٻ�}}\ 5����v}͙!�}v�I���+�*�������"_M�x�:����A}o�þ�������^9���R���O��J����KG�~9��!!|� ޾H�^P� z�eȭV�D��A�Dn���r��~Q�E^� ��J%��&=��m�|�9uF	A99������닇el���e��aߛ�B޷:�X���������*ߑ[�[bX�y�
���Qb ���]p#�v�v�,�$����*eŘC)�s���oѹg��MU�����K�f�٨<>!|��y����Oz�\�lN�/�ZZ衅g�Π��:�����U��Dp�ǣ\ٝ�@����oud�k�{>�.N�It�����00\
��S��R���3V�f�St���*W�R��
˂��g^l�B�ߋn �Ube���%��%�-s��'(x��D)�5V��6��7[>3�Y��k����{�	Y�M�B�1*��0�t���6v\�L!Z���,�q�[��)I���鶬��&άߒ���z�#�����5?\'����F:��>�A��^e<B۾SbCz�j����6��G:�/U�(+o�U��]�FP%{"�k>!rrp�TŐ l ���)�[��C�d�:y��n��	=t���Uhҧ�1�_�?w+��E�����)i�f:����!!(o��Rx��Һ��O5.,�p��!�� �e$���m�����,�0���@�&  0t(�}  �{>�sA��9i��<`5�3 %���D���߈���!��
W�*���������*B�>˅�Y����3=�d�[�ZB"mw�f��oT�"2���W��AgP�6g�>7�n�Ѽ8L��c:={��ņC�4�����̩��3_��s>����)����5#6��� %�Y�/���#9�#}.PLb�+�,��U�V���#e��Q�A��� 6����r��_����B�xs��8,()�L�zO��Gh
���W�*웳���~����Ĕ4v���̴�+F��f��m��s?N�x��v6����wA������)�X �aW�l�4�F�r�tL�'�UO��T��T�4�T#E����h���_�p��[��Z��c��P�0qa�>v����:�V�d+��W�v�� ����e8�u�>��������c�1�g�K�L#I7u+�����_"'�<N�H��O�?Pjicr�_8�*�n������<����k�F�h�M���쭜;�=�qS�$�(K��ҵ��ힿ@�kss�M�������fop¶�"����{��_;!.�Og�T�άY����P���V�߱;c�f�]�&)��Y�8�+��$�^�����q	c���p�<zq��Ȑ篂G�yƵ��	q���[���x� �#�(�����։/7B�~m"eN�|^�2O����y�j���x[��^~�ޗ/���e�����2D�@A��~���H�T�P�ga� ��>��8�uO"5D�D���2�����������mN�Y|2���F���񞔬�ioI��.#�����P�JW�Z�[>�>�E��ٸpDo�p\��ܹ��	��N��(����p��R�R6�]�
m�0bU������|�޸�]��Vr)Rb�`�2#k���2#�7,�Cf�7M���IT�f�ٔ������,�1��c"�;R: ��b�k쫉�ͭJRw������ �Ҥ֭�nz�`M�S�js�����Y�M�=�gl�S���a���<�V"�tg���L���(���-���"�Tp2��Ux�4������h�iw��O�:��u��`�+�aL�ѓ�QEz�?[6���u٘�02S^���ا��o���(v�#�"-Y+���~�@U���o��6��.��B5~,F٣��)�Wt���&���� dH⮾S�"��g�[õ�-� ��\���«��b��Jv����[�Z�����+�LA@��+:�<�ԍ}t����>^�FVX���<�)ŵ��!���i�M�	��V�J�o�n4�)����{w@��m�XD�-��y�����m��5��u�g2"��jFWU!��e�V���H�(�A���`` 7�>��0�0w�Bۥ���Z��15 Ť5�?��`�t���^!��Q7�Iw��I�-�^� ��z8���u�A-S��C�Z���.�5Z��!����_�'^Х"m_�-�zF|��e�2ŚS���~u��!a��}<%"x��̘N11�
�Mq�R#]]k����~a��{j�\p�8�MX�n]3�3uf{�ul"��� 5�?�!&�T�^��?ک��D}wA��3uI��D啖΃]&'���@@E�Fw���k��I%�Ea'lQSX�q���m�yŪf����D:A��ҳDf��ԚŠ��y.XpC�"߼aV)�n4��}���9E,�� ��=p���%f9+Y/�ެ�R��G��J�~.k%4Z^MM��HԹ#���l�*ַ���q1m�g�@��Q4�d4�w� N#�ތK#���	0v����X|LO��	������x�S��Fd%B���*�h��ף����E�p�Y��u�.@`�����7�#���8���k��!��q��pkt��t5S؀k���e�,RN��[�ض�$�-�n�'�A[������Z������D`�oԾ�	�b-:�Wk���y�d��`U>0,i�cɣ�_V ����X�z��S�H���o�DPJ+�bYU�2�9��)Ͼ5�
����H}��m�\�澼Zm`���cArA\|B�4=ʊ�]o+��).��>]? �'���=�%���W9��PB�3�x�|:?���Y���R����_Wxz+�<��_t���.���K�Ӷ��)��m �GkuM�b%�Ҟ~�T� �۲;e���>��':����	c�MI�T�D��WQջڼ03^�a�
<Cӌv�?#<�t[�@n����)[c�&��	C�����9e�5�u�~H�(��߬��1�����6����W&C=��S:(�,�] &�9����Z�-�Ec�]~��5��F��w/K�&�^�%���%e'6�@b4����g����O�?c@�Q-�}^h}�b���b+5��`��*F�B>���]�ox��jXV���mk{�@6�|c#�c �����Q���B�����P��[�'��!�[��ꯆ\#�/s3]*���m����eD�Mi�����@3='�>�Ш�G̱ה���Z$=�:���)gS�{R�gi���Jͣ0v՞��o�p��_�WB�8W,�~�����[Ch3y9�o/��<"�
�-~��y�ۻ�$7�}��������"�y�
��%�������	S(H�l�j���?Rx�?'��fK���v��ȭ���'���w�J,8~Y��>��کL>hi�\x�X=ſb�7���a��T9v=md"�de�F#a��������`�R�s��|4��f�]5U�jS����;�nν���NZu������r�<���\=ya�ei��"�>@���4�}w.R�У(FX�O����ֹW���V?��M]�m��������y�>]ϑ�۔ƍV�M'CW��7D��|���w�a��ӄ�,�fv��U60����I�� ���Q��9r৛�����-��~��@�x�G$8�]�ȝ:5+�Ͻxӡ.a[� ]'@'g��@�,�ި���2	nP������6��ܜ\��m��0�[�{iy�K���ԕ�;LF^Bvz��#��c�S��r��P�[&�mxLTfj\cX�g]���x|�={9l���-G
�gN�\[h'`X8ŭW����4����6I��静!Gˏj��A/�w�WI�6�o����P_��0���Jӳ	q	G����-��+Ȫ�c+y��Us�������-��e�MT��'�bf6��8�
t���sE����s��*g�����0��q4����	�l��4�L���g/������r��Iu��@LoMЖ��!Ʌ��#�t[]��w�35�A�r. ��/� ��E*�,�z�A�v����8�1�j���T�p�$r�>�Xw�/2�⺽�'o��M?X��{]۪̐G�Ui�{'���<�vX�G��9	f�Rw��H2�g�������jG2:�D5�w��\:��%�qx\��T�,���嶑��/Ć܀�^�3aI�0�$y�֌��#�  >����D;���$���]{; �|��]����p�O���D[�K"A��w�����3��,��ȼ��)���#RXi�D��W\�ʻc���4��`*�#5gy��\�V����:.��\���)�p"m���̐܃�/}�>����.Z�x�'���α��=���?Up���tΥ)�z�Y��Έ��Q�ћ�E�}Y����Z��&NFV�*6��E��
����7��;Pc$=���
����:q��RU%:L��}�����Ĵ��(fff`�M��2K�)����P�R��1��X���i��/��dtg,4�L�*��p|츥Qߠ^L֞N+�l���װ_~�����}k3	�� R�g�<�
p��g��]("[��H��Lo,P@�������OH�?� !#S(S� �KxC.��E�JJ�%h*E ;���j�U�3��	/m�	��B[���WE��Hv!H�'�h%��HR>�u>[��J�}�ey�B�Q�Z|�A�.=Z��������n?j	�4zt؈?k$�{5u�M�����t�Y#2����uͲ�G�\��_-��båF���"Gч
�& ��ӷLa�0�]���I7����<5�v���\L*f��@ť,Wĺe�S	�;���gB�N�?$��%>}�Ů�l:��z��;Α��~v���� �D.�`$�D� �/����{�~���٭��P�F9N�|����x�٨<"�?�/dh�[S�g�,Z�����#�^�fs��j���_��1!`�"jw���ߋ�}$��T����NǼ�_kH��^v�E����[N�9;���SKybϽ�rﱩ��N�T�p���O63����nC�X�I�a�x�tT��׆<�we���ڿ JO�uI��?I�c2�d��6I�B����,K���%l������2]U�`��;^��(�l~d�5�+O��7�\�&s֔��n�#ǃ��Ӑ|��Pȵ��E��~��#�Wa�;�r���8��k�i}@L��Ow	�ȇ�VU���,����L����8^������ 	�	�Tv���X��^��	�� �����3��/\*\�g`dZC�B0�4D�l����{��XV���H%_�s)���ƣ�>�t�r��X9'���F��P�B@J�)ÙQt�a�X�l�mv�%y����Q�_��2H��KN���(�,�.W���fD<��)܌��~�ݙcY Uxf3N���'��w-/1�B��*חp1��y"��I��{"�C1�]kEj �&Y�:�ӪX&�8�E,$���*�LP%	@�_�V��͏�W4z޿�3�q�w�.� ���ȸ�Cж]I뎠.�NOKhF�@��>7`�T+�[!�&�9g�i׋��R��޲�Wlsa�}6LlVvS�������;�D�����k1������7��2Ғ1�
R��|:��I�|d���-$k��jal@���J���E�=���)�	����}�I�6�Z�1%�~�N�9����s'<��w��_��05����L�eF�!���~��X4�du8���J��j4�{/�9�[� WѢ�4�R)gЂ�=� Ƹ�@J��I�e�'yP�i�֔˶��bsW,�:��#j���x`�q���c�6�$����՛�R�s&�=�.[l�d�����U�2��tRkuD{�Rg�vK+�$�(��PL�^��J=�S�^$P޷i]k@�W�}��d^h��{�
8-��uu$��@�#i,0���f��;sP�T�.�ҏ��5�1!@���rzo�d}�)zo�K�>'yk�TH߾,��D�����2�M.Mk^B�8M�۪5�f#����p�zr�-��JnSLk̈́����̤��������y?*M����$������8�mP��R&�Ň��p��']C����&�b%�'k|��rl���.�B D����M�y`,���Ɋm22}�ٹ���m/6lm�"�lhyoq:FG,�lBn\��@ȅ����MM�}��ZOtJB��7vY�M��¨�!���rG���q�Rs���1YL����l��-A>�M2{os�������\�8�ՁJ�' }�v�i��X
p�M+���� <p2�ք0��\�>���5�'2��=+�s�}h��H� ���ٶ�({���'Qcs�\	�,�D�V��ae������_ �n��sw��=�����bg��l�ka�@��}R�)]WA}������QAUV��R	���
����PaH(�U����=���ʏw����lT�	t���kP���_@�ҽ�/ȯ|��kI�jc��߾�`^j�sz��X�-�Jy�������Ū�OKƒ<�W��6���� ��H่Z���x�J�L�����^��F�N��_����N9ө4�&4OSo�$^����q�����r��iѽ�Q��+��I(i�/�w�j���&䪸�Ĥ�+v�糹}���C.�e �&�%�j�&��=X��@�zypΰM��;�'��� ��a%��;�S �������v��k=�K�8���_��N�0u����"(���,�:e�D����&����9�l�wL	L���T��߾�ͰTP%{��Ք+LR�7��r¾�~O!$-}�0��M�1�I�Y��N�\%���WU�m��^���F�~��L0���s���� �^�[
�l��	� �숀�e��g#À����lA�*ٚ��A���\�׹�"zC��&�#��`2R����y��)_ n@�
�K?��Wxװ�c����I��5i��u�f)q"}�a��!d�y�<���!�AP��v��T�����y,Ιg̝9���Mj�z�t�Ӑq#?O�IE��b�g��
 y��h;)�:�z�3N���M���p(䮢#l���
�o�0IP��:��� &$���*|`�g+Us��tc�@O,�k���S�˃W�>��i�`�ƌ6hRe��>���8�\Ȏ �
�۟��K��__��P����O���I������?q,Z���\�\���;�I���]��8tߝE6�i9�E�J�=Q�V:?��B�~�l�s¯g�����gij8A@�ks4o���I:�?fPeZ,vnhe�%��8�Ye%X�4Y�9�~�q7�@&�	�����L�W��%D�pL�I�B���j{+G�e�`LiS�xx;Z�����8�j�mX�w����3�J�N�$��wSH[���%�? -�!�x�Ė=��V���C�1tQ]yoL8�5��3H���J�V���"��~R|2FЎZ��e��%�|V
P���B�F�%��>`�7q��#��o=1u\��<�$�����<N:B?� <����J��ہ7�����ߝ>[�CyT�+M�������3��/T{<��CGZ��-��>=�qᘠV�;���:BΖ�u�VL%�}"Y����U�u�}M��m��`�� �]��iL��Q�H�9�8�� ]HZ�V������I�������N��o9�����'t����K���׺�� �1z0�yŌK2����%u�D��s0�Nj�\�4'�s�����Y��|@:��v�Ӷt��
���p�e\�#X<����^���
6�`��@� ���%xI�Fp~o�9Xըm���/�^R�=��4`�\	��T�Dg����A2:��!V����#+����k����HRA�l"������1�
���S*G\`�w3'_����D5m��ڠLH$��E��<`r�;!���e����Fw�p���/�"�-Ͼ<�����@�uh�0�>�gt`F1(�����犪�A7ج��l�1za�*�S���a��k$'���@�0�e��=H�u�tH�/t�6@���u\ӕ������W����H,�{G���AZ�S������vr�Ij� �@o����-����{V�7C���c�t�=a^u�b�'�U�A��eƢ����_����Ve<nAGȑ6�"���,�(���>���,@�R��Zp���dTg����W{
�d�Ʊ��J� �����7��W�1 ލk��يQ�=	r�R0��f�|;T���J�k�}�No�u:[R<�2�<x�mG��ֱ�C�c�<�Xt9ff_�5������莡w+ⅤV��H>I�2�]5��%DD�l�\h�92Q=N�k|斵�fQQ%v�l$�~�>g\�ɦ
M��� @y}���0��)W�mA�e{č��V�SN���=zqLw�Q݉w��'����["|���GSBH �4�ؕ�S�;X^��SRNޅ����&ɬY��,keGqʽ�<��Ŧ>:� (h*j���(�ɍ�7�$�����G\�_� �Ii�H�j�p�ǆ+�
�������~2��O��M��E=W�"�M2����E��.�5*�KR�E��o`{�?����ԛ� �L�S��Rʁ����[�ʹZL�H��ٖ���w�AEU���[�W<Ǵ%�2x��8d ��jt&�l���в����+��.W}Diˑ����D����@�6�^�$N��P&�P���x�Y9�V�VX��zK���}�b,���p����� >�?�.�����k0� a�ۜ����Ы��XG�1Ʀb��k�X�����W�CQ�/z,����o�J�Wh�w]=�3��;�#�b����7A�q��dxG�����G�Ȧ�j��+��w؊��u2b tYe����Ȓ�9�xZ�P6����^��2ߖQ��5�<`�k$U�0&��(q)�Bi����~�����A-\*4��T�����?�#68�5�,o	����s���"6r����l4��	�m�����[--��=CDMmc����������b�U6�V|�R���JiC�|Nc#�(0��Z
䊡xO�AW.�;�A��=
Q;&��*U��v3�
�� H�����U�"ˢ�(��-_�`&[�v�K���գ��!���_��<����#4dD�Ū8�>���炈��=����Se(D�^�D�v��<��!ާ4�g]�Z�����T+�P��m4r(�OLa�f��yq���u-_^�x�A���"�1 M�@�3��7�i�����C$��e^7�3}֋4tU�F��q�/�Uxf�;��.R�T:����U%(�S	�q���ŢN�K{xJ����Lx�D7���~	���@�k�BA���]JR��I
��6�򾪊�R����oV�i@k���U�<�nճ�u�W��u����ՙ��ߪMo���aX�ʲ)61,��V1 �y�?��nv���c�C�E4�Ğ��Y��������6?�V[P����v�@H(@/*��՝j��4"l������*7c��y�wP��U�)��]��'��6em�9<d��P�լ�W���&t��"(D���Dwo�i� ���K��@��D>X��4���� �(+�NSlW-�iD@�5ۃ���ϒ�]�{��Y�tx�̌����n�lDu�H�Vn� 7�� �r+M8�ߐ�ao��H�I�8z�*8�o�f����	������~r�Q����6����&�?����>`Mt�-wP���xLv�!� 'kE��,�<�TQ��ua�
h�&�eJ.TԂ��w:�L&����QH�m�=�d��it�S(�4�7�[���&୔��һmP)�C?�����A$�=�DPE�C:��Q�\����뜿��^C�3^VW�1M���ahj�-�+7��E� ��&��h?{�2sD+b;gO�'l��uX_��J� ����آ]���|ߘ����㺪a3J�$G�֘�p��n�
�:�V��3�Z�l��@���i]�&�~��߲���u�NȜF�j~��mqa��6�z��v�!,�X�>��y��C ���X��u�3�+@b�MZx���$Lw��c�^V�C�s�@;���:jg{�Ct���@�(jg��J߶�hv��#��1)�A:>Y<����i�PC����)-�EP'�;�eķ`�W�G�0oY�����]��72ӿM������_�p#*/'W�.�����`�M�7孍�W�'��
��,^������ X��GXܾ��Ri K�&@g��E����'9��������2F�������o��G^����9\Z�?,$�D�ϡ�m!����	MQ�K�7tm����������Y-L�i�I9=�cD�,�t����C���`G�\�:��Y�d��+D�++��Y��Z�w/\ck���Q3��D�RQ_�=��N��V��SZg�w�����qXC��>I���)�s���$&�^�&.�e���''��#@4��I0�,��^t�hyv)! w*��
�H�\�`G#�X��8��U���U�Q��jƾ�������[���i�cï u燐b�#-;Wij��������>`a��yf;�eSH��<|jw�~1������)n�4FZ��g��Ͷo�������W>��f|�)�����5��a�-Y8BY��S?u�ﴁ��6�!h��v��!]�ecl��@.����
��К�ݤ�B� �$]:PQ��oz��e`���k�
�:�աU5t�g� '������G];�f��^+�q'&������{e�mMu8���6�9�A%>��q���wVa���i�?? �������Ɛ��$M`qH�D�յm�<��!d�;"��qS~��$�bBt�)?���7��Jq�O��VA�5���Ѫ�.Lsd@� �E�����1TY{�N�g��t���d��`Fz8�<��sLYJ�8��s��}��<~~� kGʼ+�;�sCzLp��C�Y҆���1��O�� �<�y�L46�*�{��"�*7���Cr,��GF E^��Gn�l��I��Y�vZ�am�=Z�n����v��N���M����]�&m��c+�(�yzߎ�x�(�S2�8�5F�X�����!��s~\�@�H�x`E���^jל����s�w\w���(kn��V$��5���d��֣mSW�R\��&wj|�����Mz܎�[�s���Y'�nta�)K�R%!g{bD� �zl���n�m�8����/[V��?��C���H=_,�r�����:�Y�a5dr�5\:v�RG2���}\������J��j�0�&�E�0�&(�f���B�r�s>A� R��S��#�"gF�Ӻ�`��[3e��@�S kHp@�����@Ei����G��pזb���E,��v��#��đ퓏���C�š�-���c��dʍ/�,� *�?�{JR2Ia0�V�m��Z�~ 6�	5��J��ֆL7�E��N�*l�>�m�!mk9���+�3|mT=�T�7VZĪA3�!�*9�8'a�H�"0Ha�Tq����2��]ᐻ�~�Ѕ��ܩ\V��vW-���VF:E�vuP�^+ŋ*n��<V�>_$spv�P:�ǉ�i��Y%[�~i�RG/��E�%BB����0C��Ӣ���XK@��3
�ˈ�MJ̽�s���g��|�/�ΌFG����qt=M:��ٖ"���:�����'i����B���\���8��_����Y�}�7H��ԋf[φ ��Z�s8��P'�Z<�$�����0�>)2��^k�W)��Q��	B1��#RU�s$&6��x��bn����%�b#�K�%x֯�������.�y���{���A�J=rs9ļr��C���!�u�&C#����� 5�ͧgZ)�ZO�Ե<S��C��wz�h�7�������j��}Қ[G�M�7��5�zX09T}1IX��x�	���*��E�m����e�ٝ�	���ߴ�2:8@H���ߐ�E����L�Z�{���m�&��j@�]dKfw�]F�%����u1	*�;���G]��i�P�D�h@N_ ��©�t�B��V����WU1�?�h�]�|t�՘����B�9��oo��#+1����IlM�+P��*����~�8"��Zq�4�HF:�6O��)��3����O��r��� B��q*��*�a��R��[ec�!qG���3�!mi����~��s�D�&��!c���N���b��X�����q��3a�jzV���>Z�?^xO_uk�~��nLN^��G�ag$5��WO/�~jV?>��Q���Sf;�ٔ�|}�> /��ހ����_�|�	"ٷ׍OO|�<F�j���kn�RQbG}��U��%�C
�-.�b�N�ۃ����w�w6F;ж������]��d떗`��*f^�=M�>���ս"��@��3�'T�}�>�C� *0^ �k��tĜ��
�[�I�����9q	�K(,A��
�7�m(��9���(|pµ�V��e�4Zb�)L����(���34���%G���_��,�E8]Hx��vOk�W'�%b��B�n%r��1*C�yu�Vw�:�
rD�L:قH�8H$A[��w�a2��9t����1+b�U�~�C`"!���*/�_��� �Pk����t��h,Sܢ�X$x��l�+<�H�.>n��KI��Z���K�N�[�.���y+�;�ŵ�5k�f���H��l��Z7s}�qw:-��nL�J���nS٥�0a�9��&���V�dc���6T�tە�O�V?�< 	O~;�#dfL�T�4cD5�5E�V;�kL�<���}��W��)Q�^J&�M��YZfc;�n���(�2r@��ac�(O*4�U��� �d
	�-��q�Zَd.���d,Mȿ
�Eܣ�9�B�\0��/�4��2����e_�
�O��lC%*���_�+�ť>:�g}��~�1"a�Q؋*���U�	��;�d,�Q�r"N`<�V�䤮��9�bI�шZ��C�����IBgbe �՞�d�9"�V���Ȥ���E�%�!NCX0�[����?e���!Z�|�&��4'�}$�&G�=�4T����P�k��3x,�@���|9�<
:�E�ȅ<����e9�P�g�3�0��鸵���T�q�]="/��N���$E ۻ�n�j�z�>��zS#Q	/���-.���p�E2I������1��2��O}�6��x�ѿ�n9�K1�2�>!6��~$O�p���9���bB�LL8��׈R"��}�i%�1��A[��N'��nHy��N�[sv���M�$���/���-�|�#4~|����?���=�v�������q�暖�ݕ?-hNoHqi��|�cn�K��?|��!��DbR�>e5�Չ��?���1��Z��'�X��\�b0�*���U2؁���k��p=4=�`�����˴m�&H��O�ty��:Ƀ����q�k��G��e-̇�O]m4fc�`Кt�+����|Ot!V�Lq�L��^	3�S�v�#�I����k)x)=�g��^\� Bb��s����Ӥ�E kM� �J�f!���M4<2�-_x�Ӹ�=���������Hf�=��7t����KB)E=�\W$������m׭q���w�e��}"KaV�%5v|��>L�c4��Z����3�ii%�#s,IJ�
p:�8\e���:	�eA���P?��v���P�Dj~�'S�d�**��F�f���������J�����h�?��"��Ɋ��2�4�}kү��ʇ�+!4�Ɛ��1B@��mhL�m>�T��dvݏ^��a���Ĕl�cK�����R��;�^Kj�mV-��Z��ө�����FY�W���FY��8�)�`��0����54�tM.��X��qc?\�P�pN�_���*�a���#�����=���5ػ7�H���X]x)��V�n4[��_���s]���g>�k=��<�wC~���֗��N���t���fd��j�S�>�N������p�6�{ �qIU�`!&ʈ@�o&L^ީX��������T�!|򹡻�ٴw��C��B�j��E!~6�0X6tQ�e&#����[��uJ����> 9n�[�[T��-x� ��������L�]D(��Ii#�t��ێ���|5=�3N.�.�q9V���KS���/�<%6���/���^F�����\�"ȵ�I��tm�֕9���!��E�	�e[*�g)r����y9��B�=+��f0+� ���:�a�0�8!�U� ���[/io�9�?�}<�U��{�ېc���gnB"��a?�]
�1U�b�5���,�݃ym3�<��,�MvC��wA�r�ޅ�G̎_�y�g����~���&ƌU����#�1��ZԌr�)x����D�b�b����h.��^��`#^�=>)F�<^~���O���kb+���\�)�Po����.�#X��Y��邱O�ߡ��p���X6�H������V��u���]R����1C��w"���w *>�T���|���>P����}��X3�K�hfD�`2a;������X�@2A�0k3z��c8��""�,1S��쓙��թ?y�q�ƥ�Y������9_mQ^�W��S�t�U�7��D�:ŏ�}g�+���� �8�����%~ ��B��Y/�Fp�Di��j��CPi!����/�	_X��NUb�`�A���>�*�/<�dZI��6)ug""�dh{�'i��tizN�8r�)�\�S������-'3r~��Ռ�.�A�ᐚ��p��a�T�P�����2��d�N�8SQ�X�Z�fjw%:�B�;͡�y;����c�K;6N�y��Iں��Q��,���dxW���Fȴ�=�\ �ͦZ�3���4�GC���*�)��1�ņ\�W���9E�a��L|�l�Xf5:a�fT~�&�QN��8K�[>˵K�m%�O�f�aq7�P�Ӟ��rj [nΊ��/K����%I���B�J�7�̈́�����bw����d̮��P�֞�ʇ堏�"�N_�0>�׳w
�hI���\C�# ���5����+�ٰޜ�'V���J�@�>��F'�>�Z#�ΐ�5'��������^=V�=�e�'�)r�koZu@���k5Of#6���)H�i�7x���ZS䜇�7���jPo�2�g=K\����O�ڑق����s�>��J��#�3uo�����U��A2nܦ]@AB�ݷ_'���9�#l��c.C\��Ì��?!��흞3���g
�l�fI^gNUF")~3,�` TW���H�q7%p�s�M�&.�v��I!�C˛V3p�ڳ6-��U⓹���O��u�}��x�3+��{�Ym�,�;q���Y�l��0�M/�$�J`��e"ٓ���QY�Z �M/8E�0uV�H,�F(H�WS���FĬ0:���PD�$��� �'Τ�I�{�ݻ��li�
��5���բf��P[��<G���\0�N5ٳ �k�G���n⠋�D%i�����&��t��(�$�	�(I�����r�Y�JMB��D?���H�~f~-&k8WC�n̩�њ�{�Yds�!&�
���R�K�1\?1�H>������o�4��]�a��jjm�u�C�Q��G�~qہ�7��t�1�gᬡ7H�����d�1������2ؘ�r��'��2Xn�]���޷ۓÌ���r$�r���#_����!&V &���a�/p�͘�f�#_��ٿ.�,iP�ޕi��)�����U/�9�}��c�rf�s�������_��R��Iv�֡lw�<�{����H��<���kW���[���x�w���6�O�8."�>%g=v�O;�A�몱N>H�ʸ�=�8��؋:ֱmA�p�J ˣ (��0}���8�.�)��L��2���}���L5!���n���ȇ�Q�7�����.���iFY]�]�C���ަ�,����[y�<�N"�a���֧o1���G ��z���˞���A#�&����[fn��'jJ��1�æErmGn�L��{�����_s���1\/�53���F<p'��´GX��0��;Z���]�^'6H�#�J����z�NԃK�B�^�/��9;�J`��z,2���	5��Y�2�����.dyo����~�ѭ@aQ<Uy��mཧ��c�������Ԝ�n[�i�qJ��&p�}�_"�	t��O�-���j%����A���3M�J&���}�,�P|I��Ʃ�jP1���Ǡ�[.R'��^�UK<")�9�m���kb�Q�J�:i�~���_�*��b�t$����c>����J�8	�����lH�9����y��d��i��&� �C�����ފ�p�kʳC�A���=��5��}��K��M�����S�����@Wn~2X-kj�8�O:�p��RO��Ds�\�Ijۦ��R˶���#i�6�qmx�
�фz�`6���Eo�j�,fX�?E;����� O��jthʉf�	|/c_7N4�v�gLڲ7@�P"���jG�Rq;�J�D,�7y�;�`���OAڝ��+��5�m/�?wّ�����X��7욳a����$�Q>A��n;�#E����4��â����ǹZ�-�g53OL$�E�����3�y�R��}f,1#�1𫿼x��P#.T�G��m�|�_����U�6�2��1t������B,N�SCg���=�����L�S)\ŧ�O�3H|C,�f���?	���Z·?�-|�L�KꏙI�J�8j�>X��lPl
��R�}�fo�s���G���_�󍈺eYư��м�Y�_�.YHmũG�,��1LK�0�x�Ł�ez�_ ���w���Zw�"���2�����cRF��hi�rHD���F_�G��uL�%+��Oi���@k�4r���cXɢ�Bsh��c��/[-��8o~^(�)�_@5K��PmU=חc�sT8���v�׃�[�C½�Q=4�#iy��x5��l��t�g��M#D��i��U��zgFa��}�З5�h'��a����T�ֳ|?z�~�{�rf�f�;��lg�r0�v��I��v8�H����qe�[�A��%wCyX��� ���V���V�i���VJ�8��M��J_Ӛ�0���!ܲ�1�%�V�$
�
���(n��>
�Q�W�%Md`p���G/�Ո�zћ�@HY��邫�k><)�,#����� F{	���Em���(q�H�n���
���A�R�N�ŉ�Ɉ�`��_}�f�oDV���i�O�I�L�R?R���<��ҳ�)���ƽ?�r� ̎�`� D1��E.�{�Zs�c������Z?��C��e'ƽ�|f�ܧf�;c��o��l�Mه�K��>�)07ƅ�>�H 8:E_���K��?���Fq�Cv-?1�=T$[��q�FV��oV͡�Q�!ҷ�� wM&mu��V~E�h���p�oy.(�@�rK
޲���Q���p&��BP�P$�<�2����~���]9�i�߭r�����ٞ����ł�?�n1�Յ�Z�D���.�@YTx�CV������
!C��	�".�ΰo{�o�G�#�$̎���쪲��
����@D�@��c��LG����
�,@�dV3����I�7U/�!��Gu�XP<r;��:�~I��s�����2H"��N�� �WwE��^K��؝r?v�O}]у,�(�~#�����Y=T|�;P�`���p�M/
��}�lF�K���q.v�T�f�Cv�JU��������$_s���_-_�M�9���E=�����|bݮ{�ǢsRP���9�p���X�z��������X���l��'��1a���z��4�`@��߻,�)�#�,P�H|���[�򘛁%�v+���@�ď�bXi·���V��>�0�jm��}
���o�$Y�����	3���fП�$�U��/x)��)��]��B�/^&�v^���Z�x�R���9#����.Za�g3>��r���e�Zܾځ�n|QXX* �?C���[gy���ĝ�D��8���2̺�����3䩒m��W�S�-@��8%�wz��=����¶ NyT�#Af�R?�؆�5����!t�uH6�oa�� 5�ō�ŗ��B���u���'}��s~Ўj�8�����8��P6�j��|��?�����~Tǵ����*�%]-�,n-�P��;˩U��o��mc���[( GZ�)��$��plm�ʌ�S��˼1Q�a�o=9��>���*:����g1��e&g@2�q�Ȓ�� �N�r��l4��t�1r	�	3�Y�G�%��ϰ����*�,��D�)�W�x1R�Mp+v���؍��j�cV�w	=�DsV�BG>��+����hOO�G�vk��]Fq��i~�FgP��^����V8B�/��v����E���K�Ѕt^OۙR/<�c�!Qu�}�פ�w/?��,�UJ�⼧�z��	�k2�X�GU�E�SR�[��;���ݮ@�����~����d�����Z�T4�fG���*nM6� j���ݻ�_c�\:%84��3Pl�+��+ҿv8���?��PK�g!�C�Q�X�:�*�a#Pa�MX��U��6(�N���|Q�V��5f�n ����E'i��x+J-�]3}3&��j	+,���ng�\4�+�}�sHf��؉ʇ���}h(��Y��,��j���R���A�3��v�'$M�&!W��z���(�fT�؎q�^w��Lhp����_����j*!��F��]�xL��Z$2�vQ� 1��w�MH�`*�Rb+�WJ���𔠑P�$�;u��t8���/��?8`+����q�Y�P}c�#��),��H"�s�Ԩ��@��R�>N��8?�<�gm荗� ��R�7#>��X����`����G�=��ۥų�p�s&c�^b�I�5dx�U��#��-�A�lcؑ]�I��oOv��p�'̉���U�L*>YV~z.m�%�x9-���)�!�_�P�,���b�Yu̧��N����6��Z4�@m��|��煭w8��lIHvD�� t�� �Ĭ�2��F�OqР��d���$�Ft��@�/�ϻ�1�y�GQ�����k�YO��xDf�*��
�z����K?%|�����R۩\aky��F�Ʀ���'��+��:Z&��q�����؆���#��n�6�O8�2NM�*�$%M2"6<�N#�����-Vx�t�D���5����(L�^A�C4{ã�"G��# 7��z) �o��c<زUBk4Ɠ��,������U�o����4:q��O�bD��7X� �;����W�"{��?������Dk�tC�po@�G
��\�w�!�����WИhՕu�!�D�z��<�
���d��iU&�I��u�+�F�9�T�*5�nzh�U˃�t�ƥ�U�$L���g58+���H�]ĺ�I>�V뮱�2��+[��DL{F����!s�{�t(�EwວnӘO/v2#6J�Wo��)$1e'�s�Z~�"(�J�%��g87�ڻ�Ͳ)�Y����2)���q��7�Y��2j��T0x�������f�,�ƥI:VjAId���0��Mu�e����(kn�w������@�r�zn�������n�	v�b
g�n� 4��Fj���)X^�Y�$p&
����c��P�����й8^|���v;�>����K�|�L���8�޴kN�^��>m�b7?��m��z�P��
���'�pD��)�X�e�5�����s�/q��4@3r'c� ����i�Q6����� ���<;=: ���-U-������l�m\G
�1�w��w�Z�}25W˵5�Z3����E8�NqbM7ou/�5+�ׁn��_]��\ ��1�V�/0��	¬8���e����k[8�ES�wΙ���e����*�&�|�x�ҫ�|�(d���}V[�����Ƴ�~.�zX7�Vm�䁈r�����d�T���㴍EKD�՜sӬ���@��naj�7��>#ꖍ�[4W��)[iIr���d��LΎ$>�vI��Z����5zB����A�	}��������=P�)`�pR���F}����48x�J�-���j�6QL[%��M����偠��3]���i���y��^%�%GX����A/�6��¢ɋ9����	�dR�����O�A\q��{�J�5`A�|!'�+����5HG�3�]��n�zeN�Q�!�˵� �]�<��Wh¥��p��x[L-́�5F�3��^(.C���]��s���8��cj�.�T'��G�S::>+�7T�Z�!���vϨ>�ӟ��\���F��5�@�R�M�q�E�V�_$0g��c鈸H�r_��^q �$d��p���HR���&���\�LeE���It\�e�+�ݷ�M�V3��Y6�aӜt4�zD��f�K:��|E+9D\�8���v�Fѝ�ߟ(�}@����P%W�*sCH�e�gr���R�!T,��d%�'cy�|��D�L��mx��:�lW�7��L�n��*����������e"
�,c��M:,�#e���,��ɋ�.�&�H�Ȅ���}�/��YW�z�SGz�`: ���־��|8iTYۢ"�p��;7B�T*���(�����݁��Z��f����3hH����Ԅ�.f��C̵�)�����y��Ğ��@�@�w�;G'K􎆰-{۰sP|>?�&�VW8�Q��zCd�3��Q�HH�
��4E��c#l�����#	���j��!�pzAa=���M����Y��#��33�2��?��<�;0�p����9�����@B"�h1��_`��� �S�oV�@�ЌW����Z�	y`6�}9�0Q���4G'���f�= h��̳�(<$|��t��:1I���Ό�=P�Z2c�'�r1(N%�vF������-0�Sp	�����fn,8�j��IhwG��Ъ�P��:A����+?�O�)N�����6ԋmL�
NĔ�C
�b�ɷQ]��b������QF�w���\C� �.�[�&�3��F49�5j�˱sX�1'��q6H5}�2�cb9�}3U��~�"��i%wP�J;���IDD���g(���oRd�W��Vkz_�8�nry��9o�D�5�iY�|�P�hp�ռP����fC��ᗞ�t����ǫ�u���rF��t��?����6����ϵ	�H ���gz$��1%�<r`�O�r���v؛8�\OP�l�kx��:9�G�Wh2�@��>sB"���f1F!�(�Ɛ��0>�V�7k�̈N��闗��>$�UX���A$/�@B��������eK-]D�#�\��e����!�ݾ�P��
$b<pg�ت�3��~����\��y����'3.����>|�F�h?o����R�Ҷ���G�h��sI�(m(F�9���>��gx�G�9�pI5�3��f������i�B���:)$j_Ĕ���ce�?f���_P�R����5Dޢ�ejA	�� 2��	�f��o�V�vĂ������V�^�+,p�5>�x���y� ��?���2��j�a�7�*�kZi���v�ڱ,On./Ex�4�i��6�8�1�?#��:�~ˉ��س9��Ikbb��
�R"�� s�9�&�z�D|-{1m���	�&��;Z�7�c�]�I�ަ�U��ν&�5E���18cd�x��Q���g=�v�'U/���I���DAV�&�>��&h���`y����a�����-�-"����m%?�����UZQ�B%�T)v��(�N2*@/��i�UAU�^��-�x��+��Iٶ2P��x��j�Q��ӥ�|5��`�5��>{;�����5��6[���C�Gҡ\����j������c�m���ڙr�����W,.���q��5�6����T��0m"������]�K�g����>M����\��T�.J��l�aVR�j1�+W��Ό�M�ts��UZ�#s�����d�W�9{Ǟ,����M��;�1�tr�`��G:i�϶�N�)��0��ڝ���O���@��j���v	��?��2�+�L.���<j��j��7;>�,�$��T�W�x�ztT�Z�`h�6�#��)�CK��tÚpT��3������\G�\ ��h�o����\�͌Ɇ瑠���0�Ӣ�$3�0���Ҫ�셗¸09���' !3�,�O/���NIx�%�!����,�G���_������H�&T�%O�;�L�a%O��|�	�Y<�IqK�,�F�Yq��x۠�lo�k�L2c5*>���L���S� u�XBc)ќ��!@�~����;㴆;s�{��f�_;��(���U�x5�;�M8�숷{��L�~LC�	�'�lw&^.ʙv���<M愿�0�ضV���P��a�k���ֆK�u��ts�g��%m���=�qH�|�' Iex���[#J���&|vL,�,�.��P�'�����mg�7}sf
?�G�~N[�qo�+ ����,�c��ad{�)FNk�׮Q��4wO�*n����ou�(ga\y��r�U�(܊��8�Z�FKth|�(��l<.4�(�Vmp���z���T���I��J�R(]r�B݈�����
I�]�g� �|C�_\/<VFǏ~�	7Z��9=<�		I
b���a��8��m����h��;�ؔ�
+	ɢ��9ca�N�����;Q�@�%�r:EZ�!0ύu�Q���6��"ʫ3E�(�B���Ğ���?�W/��ᏺ��<�y�u[b�=��.]d�K{���9�ǯ�;���~'m�Lg���Pʍ�L��X�W�ʔ����7�B�����a!ל	[��k.u%�N�i�;����s��b���&ؼ��߆t��1�{B����y7q��Sw]9Gɓ�"��D�@V�z�����7=�1��RW24ؚ��բ*����6�1��C���^��� ř�s��D��n{ZbLb��R�}U �
\Tc9y?<�5>`4��"�=�J-����fjRŰ����8q�tL�?�&����8�~�M���IьTE�p��D
�݅s��R8�����Hs���Ǔ�2ӑ5�f�!e�ײ^o5i@�|��u�TV��n!P�,C`��.i]��8�X|�i�H}��CMe�q����0���rl`΀Bf�L�����#�}J����`u&�\p�ݯ��bJq��Ň�=�7<�a�h�+����˃�Zv�IY������?	?Q���FV�RsSmS�k�PUQ ���ޱ~������gJBP�s;��}�Wu鬟�W1g[i��^��Ձ#���4j{Q����XB�UxF�����\`�,L0���������������<�1�9}Eɉ��V�bACI!Q-�q��ar>k��B��S]dC�fF����Y:�����nyQK{�E�@e���8`�b$e��e��e�W����z�j����6�h�=� '�(�������Z��Ո�{˗^�����66�f%�(�^ݕН��Org��&/�WI3+VRV��Wcs4��v�	��j�Άٝ�ͻ��PDCs��lĿD�`}�cRc�#m����@���/����R��^���69U�<*�F�--͕�>���4���&>���Vf�zg�7�еI�5TJ�-V�JhJH|��/H8h��F�[L���"E�}�t�Լ/%z��1��_5O��)�A�2�I��{(tȸ�u��6�w�Tx(1���LdV{{6�n¢����JU�p���Y ��N4�\N���N �$�2�`�ROݻ�+��)M�[=��s����aض�LUcTZ+��.�/�!�)��MYE	A���`��Q�?ir��e��a�c�\eZ�@,d"9��������ص� ^����{�9ŀ'�M῿)Z�磟���6k�;s�<�:��ַB,��eb9Ƅe��&O��*uuG#��Ү��w}�[����8���_�(���wt�W�����^M	����(��N�4`u.Q����t�"�%F�M�},oQ(uNq4>���^�$���̮ټ�����wt���@�!�=͐e4&�̡���\�Q��?��^�y���F�H�f�W�L�J���r�K{�l�(�����lƊŭ�
P�b�1�yTN:F��H�h�"L���UI�YHt�`W�����T�m֦�4T���O:I
 μ��_�iG6��w�%#q=!��.�B�5�F1-�5��<`!��"�R�A�%�/��!W������N�+;<A&?�)1X묯��8(�`�$&���!�Rm5��Z{�p�7� �?ME��i]�@B�&Li�fn�p@�xE(@$(�%��[�ոs��.0�I��j���'������y�šWK���x����:޵ �c�+b������o���e���Uހɓp�|K�}�"�i�8���p����1i�Z!ڻ?h�n��	Ƽ��o~6/" �S�e�{�$lh�0Ɋjs���C�,	k����ɫ��rԋ��w�J��ʩ\��#�L//l3����[�8�9"�H3v+� ��/.�o�y�^�=�yn���y��Jg��mڀk���!&�bsO-B��������E4��Z�^Z�����RT�tAZ��!�y��h+�j<4�R�V�B]����Z.�!wx66s������p�v�9+ߴ�R��,�t�w�3@���� b�cz3`@/��Rf$"������	���sAE(`e�"23�~�#ޥ��K1���~Bɹ�KA
)督!j�h13�ô����*�{�67�"0� '����ݯ���-]���z �nU�1ڑog��9Cx�$�"մO�DR�1��BUYNoO�ak'�* �ot�`�	t���������g4W~�5�-�V*A�����2��GމŁ)A�>�˄�%����I �g�h��@��NB��&��Mv���(;b�,?jс��@���n)�2��f��g%�|�;i�����}l�x�Ԝ���+�J�(�C��e"�C�O��dJ*MV��bU�)�>56X��'4."�c	��o3�z�7ݬu?�Ph\k��cEQ4`޿�dY�T�3���������Ե}�8��e�DptAZ�(���U35I����K�����!~��d���6�}�����ϩzX�jD��-(R���/�a���Mұ��|i�w@}�q,ЪBn�������ihT��~��&#�\Щq
2��m�S�eI���D��K�T�$[��U��Y�&Vl]{dLS���]��=	�:���QH�sti'�rzѭ\R.P)¥�H̙�C9����DN	�H��O�:��(-�{����mk|؃�dS4�g�F I���#�-�S�39��>Q�������w���g$�����~o��Z�/\��\�� w�4z���"��	���ؾ�0��3�g4ֲH���F� �O�2��������PI����҂�j�C|?�N�T3i���]XO}S5����E]Nz_����N�/=�ΧW��G��ێϦ�(YW3��R�D $�2W��`���w�zH��/ŗfVY 9�����	�N�B&�^��ӑ�bN(��5�3"Q(��Cg�7Ș�x.u
���)���
]o���Ӗ���+n@U�$	��>|*�#� �>B��&m�z�h�v�������'�2b��v`H/7 S�3�u���ɫS�Y�Cs����)�Q�S��n���՟�hlN�u��0�i�ŇM"��B�fL�#�������;k���S�vI���rh0+�aۧ���5e��!���{������7I��
ƖeU��wǑ#+� $�}�;��mlg�{�C��-+�J*s<l,)��:�x�N�}#D�E|#�J!��D�k�6��UX;���Ԙ�?| )�EDj �z�!�Bzg�M�)���1�F�D&���?P�۰�{����׬�l����9���b��<[}~���$9[`���b��7�a�Ը*�Z�}�d-���m{��5��'Kc��4�i��@��w�'�$Jh�`��Wx�&�MA����D�)�Nl�j�Gc��=�h�	y�*���e�IztͅK���Z+�O�+~�RQ�b��j���4��(����N�g42���47´��'��!̤޺Awٿ02+S� p��s���c]�#���5TxY�>@qUZ/�t��S�d��qܵ�E��5
�����&B&z6&D5�E9���*��.�B5	Kg����Ĺo�Q�dj�D7��٠���x�V6I-���M_u��Yeh@2��{|QO����		\�����s��/��_�èD�[�Y�KS��<��z��U,��y.Ho+}��+F p�s|��G��_��r�y �`�D�v�D^�������_׈�m�F��m��% �Qi��vk����{�Gb�hS�Ɋ���ɿ�Bk%�#6G1�Y��xXd�Y]%jFDt�(l�A���@3׾\�[�̿;�������ǀ�3N��YZ4i�k�ؼ��5��8��Ǟ ���U��"�|���dMW����S��٤��"���;�}N|u,J��R��0�Z���{w|�s��� Ml��IG��X7�����G~��Q���r�Xx�=u���De����y�Q�ȘYg��?��@�/#p���:�����S��Fr_�g�괫���kK��:����*{�cQ�6?>��Q���o*M��4��9ڈ�?��kF�Ő�����o���[?˓~{�c�)��ur2E�yc�A��Ur5��s�a�t'���f�|�.=�U��gZ�($/�"�9�6�@Bt(�g��0�q���?f.l����6����tj�AU�`O�Բ,�2�K�}4bC2V�ɝN�;|���&w����J�Z��Xw8�4��@�q�6ߘ�Ե1s��ζ@j:�a^R�g~����o��/�TL$7�od�"&34�`�M��} &<3-y�m{��k`7@�|'�q�P�z��աc�3�D�V>�h�!� �r���"6-�ڠ_���I�7&-���r���?�L'`W��1$��o8�F�l?��0us�����
ۤ�<(�p�O�(A��q��Ը�MI��BF�k���<��}�N��"��y<j�g��}i�m\����B 
�D��]h`��g ���Y5J�����l�>��~�:����u��H5AF�[w�	����`ڿ�dX��Y~Ȏ��,�ls:�M>1���kq���y��c2ӷ�j�s�0���ԯsr�0Y����-i�E�I�9��"�ޣfa����_c�[=;�.u��
ۂ���hK?�	�F�9rS
�Z�Ȗ��+�̼����=ᑘ��_��?�/+�+�X���ǵ48Id4��J�t� ]�g��KF$�F�1�p���mBP_!Օ�q�$%�9�RqG`��D���~_��1�ڴOoݽ��u��U��/.� &�t�Yk�?�2ѷm�v�rs�-�S1��|�f�@�<��|�H����;�m�}��vi2/eX�`�ί(�ṃ����}�2��4+۟a���X���������� �U$,����Y1j��c�{�x����2� 8J���d��[[�'����*ߢ!����G�R�CN�0'�R�))Q��~���j�^���J�e7�_�S�i`��Q*�y~�T>��_s�d�2��8m�}�ެZ1R���i���J4{A���[��ʐҞ��������&���~��
O��l2������㵙��C\��h�ց͍}[�<�_��Ҥj����ǰ�����tj5�]hX�{Z�";0��!r�y��T�4M��h94J�q����B���g�"R{���Ȏ�b�;<|�b�R2U�b�e�U�aAzT�����(����]���!6kҋ{��L��
�C����P�5�q�Y�J���̈́y=*	��;��4�I ��ҹ%B��F��Ҡ��r���=��Y���Qa%Ok�2^��V�R蜂���_�;_^��/��u�Z�0�[�t��1�rR��f[�2��+	{��yE�}do�2�}h,C9*�_�
�k� �:��2z��1�$a�1�(uy'�����V�9�V���M�5|�A���b m��m�Viwmn�Ui�?�f��������!�@�{��Y�2��F���"�_�H|7\��}R�ڽ�r�:<#֗7[A0���O�S	=����!K:A �ST^�)�x���0�9�sC�!3�zs%��x���>���z�T���ǂ�%U����>^-8���#�
��F���&��\iQG��;�#���@��ɶL�N��s�g+.+�79i��nz��c�$��1%�_u�ܧ����� j�_5��5�-��\%e��C&ϛx�3��Y��`��!+�:�]�7
nRf9@�լ�L�^������7N"DR��z�e[��s��mmI\ej������g�l�* �LSwP��/,K<5�"����*��};A���\)f�Kt��Fc��U�w��x�t �۪�X8�&w.���:���dF�j����I�x]Yh���ި�N����X�<�9;���Qb�lkP��2F�K��PG��|TQ��I���ş�'�)p���j��IdOZ�;Ut���:��/��U��X\�ߔ9��4m�/o8� 9��#&`7|�`9)�T��H^ɡ]�LW�-�Y<�wz��N� ��=�,��E�d�~K��'��A���W��P��\
}�#5�ag�*7�{rO��P�Ww!�ZMi�2�S���W�A��.���S���B�� �*r����є�>	�Aoޟ�����{�,��
�g,��P8�2��=���?{�i�����֯�AF�d��)�}����Ei	I%��ٿ�H{�J�P�d��y���wd�P�XN܇	������?�>8Le[�hw�7�$��3"��ǎI	6�����k{�%�� m�r�(�$ᕸ#8�oX��Y ��7(��V�q�vu�X����*e�T%�<�IYص�@���C�{��p��t}9;�� �+�c�YEp�iof*�[����컗�m�l��E��lՏPɒ�3�+8�T':�����0�5MKɩ��M����5�Lq�˻���o�[��ԙ�QW&������[��'.Үe�Jm�|�(��C�)]⅑d��󘖣1C���]�Mo)k�Q�tF�~�@�󁂳��+@;]3ݤ�Ve'l�fN���W� u�
Z\e�?�~^Uo�h�4�	�V��	b��벓�̝�$�h�'}���qo�'��%���'��}�+��6�8�s��E��!�(gQ���c�7#Y���@���h�Do|k�p\W��7K� \�e4X9?xSѨ�>y�qX�m����6yDe~���Aù:�7�̹A�3WY�Ќm�����wtL�'�xӱe��K�IT��Q��σ*к���&�f�*d�����u�[������Feأ�"���k6�9���\�я!С�|���)��>�W�-c4��Y�=+��^�'��-p�$?�m
��}ۭA�&wm����]��������/�4�7^�ݐg�O^��h);���*�W���<�S��Nv����ƍ��U6�-O�d;7`�;�-��zA���
|�( ���e'�mQ��L@$��.O��A��
Ԝ�����-�
�ѲLu�������%*�����Zdvz}���k��d������Ph�n�Yk�9�C2��G+=��������K��8:�������N�VZO\DY@R�L�q(M�jY�
\��^����"b�r>)�E|X9��A6n���V䜃7f~쀃^��B���/Y�OLy��������^)���}�ޯ�{���֥�V� a���)�0m�0��8}������V8C�Ҵ��М�Ąg`,������K����M}n��?�;�^Bp2��c�꧓�T��{�F�G��yy\L��3��׿�:�2�*/��b�h�Ȱ�`MX� S��
�ԍ4��+��@x8���r\�N;l�u�Ey�6�ٜ�fJB��#*6���L�1\	�% �9�ڭ0�9�"�!�߹�������"�5F28�`օE}�q�Ь�3��\��|MK��3d�!QWE���s���%MFK4�l�h���+=�3�L��������i�S'4d��wV�oUR�TL�>��Ě8�lLm��'m}�����v�҉ro�,@��ڠ��q����2���Z����[�0S��XZF	Ib��M�V5\=K��<������ЧOYe�a+���{���N�,�PϩdJ|��Xx�:�\��Л-�{����cIm������a syR
�-�����/'H�{�&5A�覙�'������/y�j����em�e@+�_lo;pBAw��j�@��D�V*���o����6ȝ��C%δ�ƀ�Yw�꪿�̌v@JF���$cJk�k������S*}_��i�Vì�We7<T�ñ����X ݮKlai�xGˉ����?�KE%�TNR�e�K�(xa��f|�\RO�UŦ�ޖ;.H���/O��w�!�
�� ���&q����|(
��O0y�H3)= ��n��J����.��\��з�w�m32%}ȯ�*s�,�D��Q��VxU��s�i~�H����s�7�&����n�xHfK���O���0�A�͡ M#ڹ���U�.��` " ����(=B�}��tQ����D�ry�8��Bzp�j��ی&��F9��p��L���v�9-��Π ���w'��� <ؒ��׬;���JI@f��Ӣv��40�B"8�����ݤ����T�ij�p�I�C{�c���C��>�bq.��vpf{]K�
�L��ՙ�e �0��Fb�c�cB�Ǩ���P�Y�&)�A�b)�k�>ɪX�QFzN�<K�����%`��2RJ�p)�zph�I�6 �BM�v���wb�P� P����!��4;	�4��S6m�u�R��-���9� xҎKۡ`�S�t�O8�41/�/�M�҅>ޑ?��a��������^�դS�N��B�m�`��bl>�4��q;*����VMuj��0zt$������Y����Y�]?�*O���`��^�<�WU�'͗��֌e������/�`��� �A9��j+
�wa���{��;�k��F���%�!g�j���:�$ŏb>+ʊ�T6��Y�D:;�ߑ��Q3�R�f��9�u�+��\�歜xl0��c�V�]��˽_����
p��op� A��䈘��1d^XB��i��v��!S�q���i�V��p�g*D�S�1����'c{�F_��I_��5�届߫p�P�y��f)���N�K雨����[L��3�f���J,��҉�� .V�>a��d=Q��aE�EU�ȵ�wl�J�a�����o�Z��r!�GP4�g�6�=LtJK�l)��plg2��C%5���kY�~�_~|������f-+ù��C��H��e2�h�f���^�	ˢ�K��Y��j��VT5%���Nv��GB�������L"f$�c+�OY�O���~`M�DV�e6����(=������l?�+�)N��Ԕ�7��#vB�OD�Z�1<���Wذ+���A�� 6P\ o8���y~6O�#DH͒�OV!18W����M&��̜:�C��Gj.�륃�0��ՠ[�ڡ!���Mv�1[�u��ň}�����?RƦ����B}��o��]KG��/�z��+���է�`7� ��>�X����w������\�e�,���	Jd'i܆�yɛ�AG#s.��E*e��7�o�Z}�%��<�@�����7J��N=t��Y�!6mu�Q�
���bδNj> �8EYE�~a�����m�#���R⮁�ӭ�KS�jF�t��2�|��7��Z���#�n�o,͗ �M�"="�$�����%e�G
˕	���{���'�4�y�������K �.�(���W/�0�7�5�jJ�2�����Z>����R4=L3�u�e��7��������(�=��d�ug1B� ��������V}5&�<�&0<z_� �#��R���)�˝'B�`�hQ�
�	��#}$DW��Q���-u.P�U�� 8���I�pD��kTJ�@�������X[�n�j�x��{�\U.| �8��7~�N��k��7��!�2W^ ��D��R𾉾'�4DL�{���{�9e^�9��.�җ_�)���8'z�*j����(Q"|��9ա�P����H��J�f�JƂJ�bz� 4'b2�����Z��r��v������TFN�8���ը��I^0�������p�|���6�2Є��-u�p�4"��۔�p�y�6����3��s߶��ɐ�1d�6m�E0���W�����ǵ	���)1�hm��W���M�B��ǅ�鄊p9gy���S88���,�y�w�*���lv����"�jՀ����y#���ûG�(�"ʟt���`��b�i�g�k�2��)*��!շ���Y� $ݰ�-%���J��Y{uj�w�A��]��N)�Ii�u���J�~�s�sr�"0�_���h��%J�VgYSޔ���]Hn(bAz	@�\���6��'��������r�T���=0��>}p�&�>I����J���!7������(8w����[�B�"�{���{�A�2{R	9ɔ4l��U��H�j>� ��GJj/�Ck�(�N����2��q4�R�w�8_��F�T�l��p�c\�>��B����v˾�>?�q��,��><�˾29;;{)��I�/�� ��Fӣ�5j�2i�y��g�\PM(t���:.���6���z��J�L���~u&t��-�k@�Y���%��������Re�{<�e<-a�gSJĀ�Y�_[�nzL��K�8n�u�nJ�xM�-6%R�e7_C��Y���`ǡ`�q��(��pƒ�X�5#����fϓ)�F���[ځ%(���3���i���i9�x\���E���Ka�@D�\�x1:���0����Mͯ�@1Ӄ{	�'�hφyR"�xqG���`l(2QR�;C �c�	H$��̹4�<���=�=]�=>r���T�)��Ȓ�p��,R������ @ �[w�u�����,B��o���60�� ��U,���|~q,�v��@I�3�>� ��1��3���h'�b:�P�Prm�K�-�ž�^��M�z�����&�R�Jx]�*�?Q�>p`�����RA��>��d��x��۱�4�c�C[o̶H\?^/�i�U��γ��vvM{cٕ$�&��
���9T� ���J.]빶O��,�8�����{8X/�C���a^���Q���h���`�Pѥ��E��y�R��lc(mA��7��;vr�y��s]�q��:�G���?�7j�/׳-�%UDO��3���7�Ė]'4�����r�V�x7?��!n-�Y����P}�khڝA�$%ȷ`�׊�$>�a�{�ɗΗ��8jގ����K�An�b�F�iKg�C���]H�UPmԆ�9E�5��V�36�ou�.f ��4HT��믧���U���3Np�݅�2�U���� ���E_��٩���:;EK���bY�U�{z#�hS�^��̺9�FU��vG���v����E����a��z�*~�[ ��d��M畗t�m6I�!�'�#������N�(��"���	�y8 2�9�@=��	�z\�%�7*N\�E!i�mk �Φ�e�ػl��r�KYU��h�ahcQ�z���j��A�Q_��θ�"��>=ePpM��������T�.:h�:i�Zm�j�!Q��Űz�?�IO(�H>��B"7�(]�%�!��J���Mo�Ëh�b�F�1T���[XU��#�c�	�V���*S7�Z�p~dbv�x�;ܙ�������//fk��uG��NAw��x
��o�_v�T�
4
�;Ҡ=T�l���a� R����sUD�ڷR�ؘ*	����1RV��A��*���4il��p�K�rB�"�^��]�$�G{&�{�@��|�h��s��V��8���3��z��_P����h&��\���"�YFВх�u��z��Dk���o=i��Q���Q2b���٪������y>�t��?_��A�@N�K���sp��~���������ZE��\JGj3��ඍ��g�:ͯj��_{2�1|i�4Mv�Fjt&���8��/|��v�8�I6
������u�J0|k�_���*�M�#�#6��Wl���ըn�3P�﫳��+�|����'����ᨛ����S��ì��F�m�K�Q.�*僢�@�|m�E��� �[�����J/ܸ���d!-�:��;�">�wJgv�Ǿp��K��o��>�qW*F%�Oۜ&���{^6|���6td�����3]�n��{����An�`� l���+k�Ї��𑱽�e$���%�E�����P6��	j5S[O��:9��3A�N�˼�fm��`C%K�ē-���Z�ؖ�7��/��������*k��.:6�A�r ���c��M���_�1d��������If]T�V\�g<��D��>�I{l�pݩ= ��6�� �<×W6H9�z��1�FO�֩M���O�6��h�?������@xow/NTRj�Cy[#\ӽ۳���@�PL/_�Y6k�#k����E֌q?�9Cr��P���E�e�1�2E�J�sN5;���E��ߡ䒎���?]�ZI-G�}:>�Q�yS'�1�9yj1�\�4.v.��1��1e���!X�6^dD��7��UR�v�F�D(z�
X)�q�ԟ:KL�@��3�7� ���&c�@��?�5��ʝL�aeq���$�&pG��:x;��_h�r$_�k�OP���9��Jӕ�QL����r�������V	�4-%�L@`˨!��e�!eV��R��'�NwM�� 9�}��A܅�ܹ�B�roEl��D*��li�sXu#�z3�0C�=G��y��C��C8�j%�8�8����ҏ��ٯI�i�3��ѐd�ó�V��������A,39��塡1\�?
\�Ȩ�%<©�75d��|�Lg�-�����:q�K(�X!�e��g��f��D�7Z�XO�B�����>R�l�~�i�4n�V4ӌ���b�Y.��zv��v�^]�K�]��m�~aD�(�c�i3b�[��P�1���e,�3�~bv�	�b����d�c�~�+�hM7\���7�x����'�&�^2-�Z�ǎJ W�OB�"�vz4/�-s�a��~��uR�'w���nu�'�L:���mE�zW����%�0&+
ZPsQ��!�6��h/G���8�\��L�k���W����Po�C�p\�0-o[���p�g���P��m��=�W0�p⑫�!�f�$(jê=7�$\�fp-�˰�8��e)�w8��8���8����QR͛yaA�ƔJ�U�>ā�@ @Ò�(q*B�l�I_sD�R���ι��!�z��L�  ��m~ \�h��[��-Il��(� �L�8�����С���Ebd�b�E^�|�ɕ�}�� �WRi��`�ۼ�ܴN�8s�@�e��K���5��
OR6s�r�WW������w9;�$8i��Դ��)��� i=� 7ל֕�S�7�H��9��4EB���՝4��ss�=�X��hN�L�Ni���pZ��}�:�/���78�ga.|�߅\?5�_뽙��=i'RM��=?�P����<�L�^fc�W�@�T�gH(��{';#����^�z�����jF�W�ew]� "��u��&S0���T�a=' Q��4K~)o����$*c�^���x���i�/���aG1�g1���r����� [�>Y�<�^	�^!C,�����AM�wU=�h� %�<-n�R�����c�Yrd/�A������W��}�kﻗc�y��ln��FL��$�=�)㐍�]��wv\��(�)O��}��L�3D�j�bN���!�j<��r]J%v�F��_�qcf5qGĪ�\�Z6�_{��a���g�=�H�a�=ױ ��õ\�xk\;X�!7L|0[-_�IY6��g����ˆEt��$d���8Xec�JL�q��W�}�/��Ǘ����t�����8�J7?zo0DG�ߛGؿq�.�?2q����R:�#
���iy��@�RTVb�TCC�J]��Q9��n�w�/p,[�)�e�|Q�T=��f��S��}Gv���k2����|Jēg$t� =�?Vb��N��N����ޟ!N�8�����}x&ٰ�ur+���ώjؒ����/���1
��U�(��d-G>{�E���w�������-��V����B�Z� �en��[�$���^����l4xK�,���)����#y�*��׏o���QT˩�\ӡ�&3߾����7}"���R.K EHA%	���I�L�#6W�%B�h���}I�|�F�b@��b���$_�%g�@��q'�\(œU�-�كB�l�
�Zr"ϼ;�J��MkMHDW۽*,`��+}_t�~�ZU��W^�A#�v�ڨ��}$	jM.��'�=ؗ��ck̽A˅��'�u!���%I��B��1��n_���f����R,�W{�Jg_Tk~�1�{�46��s�D²��ȼ���	��(��K������៷��[�,��L/s�7|��kr6��.�؁�@�֐�]	g���S�$����o�q�]<������p�R��m���������`��/�w�D��s~���!���o������̖8b�D=E��b�����Q�o��S
p�A����gj�Oژ�(�Y���#�dX���@��m��!s/�`M����{����+�u�,Z_�f�Nynl�omc��1$�ʷ�ݫr7��?b֓_���Wv�=�	�;�C�f���eu�������[~��Ŷ���X��8��0�,:��9�'�{����F������]��|��@�:?�uJ�C�i�Z��}|�����U��9���{�)D�h.;�sBIJTC	?yk�� �0Pc2i�Y0�/y�n�HlQ�T#�Ŀ�dДK�[A�%���ܳ�10��jE�Ѭ!�0�����6��0��W�[�!k��S�#�1,�_�(]�:O2l�z���`�>�W�O��S:!2>u,�\����s ƃ#���V�2h�9��B�S)��������L������YkZ#��C�J�<���7�^��GU����~���7�J[�:��B��߷c#4E�0��ڈ?*4�:�罓���S�,�ٲg<�q�X�
�,_5��s�u2�Fk��p��0�쾾��ÿ��J��7:6�S�x������u'h�@�H���yÃ2��� ��7p.D�n��ױ@�#�\Y~��]١ޙCժ���]��m����j(0��+��#I���^��׃���}�߫�@�Qn%`�nS�KbӦA�1}n�+���Ds��t�+7�Nd�n�c���e=���Gp��q�b{-���'EyU����N|��	I�x7-(�kO ?KѴR��� Փ��_���Ɉɭ+y(K�X�;����K�k����Xj�L"ڸ%<.P��&�yH���48)!� 4�&�^���H{%`f��Y\2�� �����,+�	�l�f}�U 2�#Nc'i!�ư �����x#�w����`ű�joc�qc�κ�oև��j �yql�V�E��������+M!܉�����jQ⇦& ��1	��Ś��|�P�rf�뇌N IKx��a*Í<s	��-:Űj+.��x���X}�"��
�vGs/c[��@l�,�-16�ə)�.7�F�IIo���x�5�
j�0j���~��G9cJ���z�Ɨ�t~(������ߛ��Yp��x4��u��(|�n��N�m؆s_Iy3�P�B���wk��h�E��:�W�"<�8 ����GY�H=yݹ��vP�pïߢl�k�
�c1V��i��}):����	��9*���n�A&��'_�`����Tp�O[~�b��6[D
̞�[�k�f�x�ֹb˻���<>k��53�9����h�˪af��s"f�`�{�`3�iI��n]��	@�E����u~�{��]%�/!`�M�Q�WɈ��P��(t�B���񯆢�YF"d��]A�@Z#]�E�&�"�g��T��p�a���kÊ��
xZ�}@�y�R}ߌ)��?L���-������	�^���#@�mma�`�"#~RF����(�D�Ggn�~��6�㆐kD���d1
�@q�Uۯ��]� 7Ф��5*�V��/J��LUy����W��{��E�� �|�������?���e*<�����8)`:�U(evK���Ԋ��J�,�5�Z���y ��ḋ���Ίl ��ǀ=��� H>fB#z𒣬�m�MJ��CR�.�>9��Dc��M�>��|9�I���������L�[�3�Bܻ��*�:1��$H2e��[c��gX��C�ނ
������p0�`�X���f����/��d�a o�i;ɳ��^�����)�a�3�ۨWC:�.�m��u$��h��_���.�7��z�@O�,�|Ԉ��h ����(�?�Jh����+Jz�@W�ǷTH.�;�ie2�#����,qKOҹU�\e_|��*�����g�m
 5U��0yw>�Y$�,�����/�ޠ]V 9���o+�W�E4&���ˊ.�VQ��>{�����2�����yhK��>���:*gH��哿V,2������1�{���ʵȵ�7���r?T�u� �*�f?b Ql����^`#�kb��V�B:�v	��j�f�ڛ���\o3���(&ҵ��\<y.���2���x!�e�Gm7^�Һm�'��9}���`tB��1㙬�~�{�����/���ׯ�Hٴr��Ȱ�$�0X|8
/�uVޏ>�;�'#�F����g�q/�92��R�|6`d�����Y:㌢܂�5��$��e���,Pze!��u����!r^0rK\�"o�bj͢wѡ�*�r�9_�rL�e�u//5ѩe�fI�[1�؁ڦ)	g�q������ڔ5Byw�gTUG����/�hAѽ�ܱ�x���|�H܌O��s����(`���U3�~�����	�-CJkY��;a��p�lL�>�t�wԳ�*�oƀD�"��ݗ�񊋲+a
�b�>�m��L�����Wm�=g$VU��`�#�*�唚�4������@��P�?[����!���؊I�K|����� �F2E�[�X����J3^4H�Yd�Է�M2Ǐ� '���Q�RIb���DH��S����$�`��Í�K-���Q4���q���=�*����ݤK�^�T$��Ј�!)�6�>������T��X��*gb�B�y0.�BR��.h�r�l��D��+�6������o��ٖ& ��Cr����JphL�-ym$�7��
�����9Ƌ^�۸���D>R:�}�m�������$��]4�R�0`(nLH��	?���D�9c�T�0#c��`7�a,� o]��7�h�+��-�ߨ	{}r�<N�˻˾�0�|ȟ���9vCeS�m�PۧK�Q��*C�]��ݗ��K� ����!i,�a�>H�뙵�IڞX����
�':ī�-rk[kD1�E�����P �c���ߺo$�fz6����+�l1b� ^��d�G�Dyq�H'�JD���*�_n�z�knhA�&]w���ݥ������
"�a��U��������+W��I�r�Ac��t���ӽu�0;��_8K�b��ÕB^��*���Jq��*��{~ċ�k���BI6����~6��U*�b��2�؃�S��I�H��T�nD���^% ���P�p�úcq�����$j�Y�?�5y���"!��t��c�xt0@��Ug��"�{L�t��»��D�:k/5Z�E���L�{�ǰ�݊��<�si��#��N`��F�h�4W`|�&�dNY��끣�6�3rr�bw�VA�;��٠��BiP��<С�n�p�ԽA�O%�s0��^F��
�|���C(�}0�}��9l���9����n��ށ��D�+�,'q�l�i:�0�	<��49���.���=�^S�� J^A;ve�%#�ڦ"�%!�~ظDa�p
��ם� ���&�p$�ܲ}o&]v.X{����MPG/�Ӛ���ic�5C���3�E;�|(�!�٠�p8�-E�y�NŽ��J�\�V�S\�L�BJ�|�h`��O�����:�m�p'�E�OJ�r��0�e�t'Z�gu*���t�
a)�e�/=�5RZ�&-�3����q���j�;��z� 3V(�~'��f�JFn�
QW6O�|<��������n��J�+'�pS�����i����dMI����W��{�I!�[�rw3ß¤�c*$�Zu~]�i([R>�)�2W�?�VC���I��n�,-��ʁ}�	=�O)����������=c�1O)��{��I�������a�zd|��&��['I�x�T|�5�xA�p��b�%�H�(#�l���$Ɩ��^k��E*�q��Iq\�[�ti!�r��Fb}da��H!�����@K�e��9Ye�����=t�q2.>��f����}?�U��~�֔�RMI�g���k82�܎���s�<�R�?�_���L+��wWעS$ ]�U 焵���6o�6��Ɵ>C���Q�V�M8z��U>��B���_�ח����[ ��⢛���Gٳj1�R��h#(��B�g ፬)�
��Qlr�"����`����&�:�+�}�ǐA��&�a��>�
�28�A^۪۽5R��<3���|�V��)����6h���
NXo56�N��∪\����˕de���\�|��Ss?��\7L�2�+�����t A],� U
�Km3��(�U��;��u����kF �G�0.�x#q�������>A:��|���Sw:wb�叩|���$�Ԫ|,Q��I�-���DT��L��k�c���2����@-d������$�p9O��@v�zT����ڏbу�	�Q��B[�ۿv$�D8N�Uy�v�.Ә��z��h��[T<A�[�T�/,s��ӏ�����z��J�����k�c���	N�d[B�]�,��7\uS�بw㘂�v�X�Ԥl8fr[�뵽҄*��^B���/��T$s"~��,�X������L���5�y���bf0j�K�J�/?����Kg����i�xG��R�d-2��X�|�m�9 ��	E�u��kʋ�*��ݿq�k�:hp"�̆�콰(6���.�6��#Df�9`��B�u4]~�
`,� u}��K�0,3O?]�s�8���c ��;��\Q/�W�S;����f�q?+�O�T,�!9es�c�����o�W���m��	-�5=�@���U��C�}�b��g��YL���� �V!_�[�.�VdU[qBE�*���L��L�s���l
ݘm���)��-��<�X�x+DB���bYo((CEHIDz��d��M�i��sp�dUw��4'��$��L9�<�	����qy���3���qȽco��q�~0n!=�"&�8�Tx>O��磹>�j�����^�L���okr5�����*=����Ɖ$ު@%[<��ҧEg	龓q��R���R��o��b�����l��=ĹMk�8^J�t�#��z�%P�PO8KZ�nz2L�(�8%6���rEM<:bl���#��]���<�SjI��R���������
�"�L�y��RK܂��q���h�w9P���}J8l�~��W��<̑�S�5|h3a�$p�gE�=���^$��o>@X��U�4��l5%<�a,j����{����ʃֳ/.�%쐄R�.�R�u���#%�~j�[)���#&�o^_w�ºy����k��;Pő��fRťhb�C�)��S���#!���a�XX+��g��hͬ7��M��1`�n�	�xCGY�<��>WP:g�R�v/�K�s��	������%�Wꑦ�h��������.�)�}6QRc���-UĽ�Z�!���0V�d���	竹�K��8�����;��x��-����B0�Ŗ	�z�x�T#Jw��)�k�v�k�,S-�bT��������5�\a�7P\����%���"2>�|$O%�ңs�ߚT����acn���o$vMR�Cʊ�?Ɠzﻟ��Y��udl�
����31���E��*(cPc�N���9v�� �+Ar-ME�3��6�n�hhK����V9��>���:�g>p�ؾ�Gm
�i��(��Eؿ���g��
D�[��cm��:+��w�	�*�Ͻab�K>Ն6*t�c�F�Ҩя�?y�G�[�@��cB.w��vN�d܂����k
g��s�t�f��r����ڝ����a�܀��P�K*c���%�]�]�	���D0	��g�V�,��}{�����Y���l��5X,����it�%�N���:��[T���'ê�����#U��X�cݓ\T�������ֳٿ�r�d��(����hF�UV�r��$�[9���Q�	��G�ZM{`C�I��2�c|o�'\�ܪ������|�מb87����%8�P�ǹ����/7`|���&�y
��6���rdS`�ܱ������ӓ�H�j�B^�.��}�������4Ӫ��)o��� l�1�G���A<١�h�6�Fūa,���2wC��g��TD<u�����L>5;�N�R.�N��X���0�)��ѹ|����7���^����������WP��-#�x��;� (^��TIK��v�N�"8jt�.�\�Ϣ��D;F;�Y�5�d��¤ 	��W��z!:p|�z��0{V�Ê�h,�J-|���;�����A��/o��6}�Q����!��2�V��'@~��@��WQ�ߧ4�:�(rD#�ۢ4��,eT2��58$7JMjhJϗ��wt���Ju4��%bX���Y��Ŏ�g]Y���!���K9�x}��is�1HT����\�-HD'+�G�{��KK�a���C�ߔi��Ь4�^����-��M5��{�֏�B��.�_d{D|�d�O<ǜm�)�Z̯��>�4Y��/@)l�~��x�����E�Zo���`QOgv�h&��(L����Q�.��1O�۞��I����p��(�A��`a��g��]������aC�t����]DV�w7IXH��� 7�&���b�:(WF�͆}�r%�EVfY�n#�q��|i�ـ����Fu�o��EV����#ظ�������'F�>�f�
柰�>�s����~l�������0(��	�n��r��P��,��2
�T�Ģ�upHދ	�2����6!�7(U��G���z��v�����t9����4H�[���O_���i��u#1�D<�v�L��eU+���m��VnB�V��q@�ss'�ǚ�q~\Ĩ�z}�?G���@x_.��|\Z�q�dK	@���}�q��7jG$��9L|��R������Է�l�C)�j#"�q~4i9��!��A|]k�n�PL)!P�I2K��(��^����\�<��q�$�)� =�Ỹ���Q��BQ���S�(3iw%)`�Eb����xꒈ�!:V}Λ�q	�L��da��
#H��+�$�s��ګ�7�����������4Q]�����f/^W-�lʓ�H��
�V������G����쎛y⋛d�\�[��;�ǞK�ԟ�N�^wq���Ґy���Z�_U�Q���fBZB�5�+��Q^JĶ��j|���x���Ø�&k,�����$�V`�0�z{"2�V�d��)��a2�ǽ��_^�9�
d���kH� �ˊ�k_7���>I�����*-�q<�������++�N���/Cѕ���������Aōy''*�Q�-�H}&]BZ� 5�=6���~O[��^��dQfN�3O�=���~�/vj���+y�v�TWc��bԳ�5��1�dBN�.��6��u�B�b��q�j"@�d>g�ھ�V4��✻_˾�ѵ�e��X��wx��OՕ&r�6��:��zd`�m����>$8��35��<��jƨ8��ɩDc���J���}y�+"�vsV|��E��$~��׵]h��?��������lw�F]L�V�w�"�d\ݔ.2(��(�G�@�x��6� xA�JP��BW��`�kb���W���4�@F����}R�:U_Ckzz�DۍBV �Հ��l�)TJ���4H��8�7�+ '�.�,�1�AJ�������l����Lx�9���26���ۼ9��ɤ�M��#�5��>v5�
�È��qӺC�B�^��!��bm�t�Ŵ���hм��Ҍ"�>�%4!���y#���Ot}���yi�Кg�i��`=�y/)&�D;s�l�8���8X��WS�v�/�^*(ah���;���ToZZ�'v��4qNx
ȖYګ��>��A6�s�X�dإ�Ҝ%l��@:|ces��_>X���Е�뎍n-q�����L����rv�&��^7����y�T	��oc�����
Qt2�Jݟ��v���xx!΁�*�KE~*�����9���-6�Ѷz��)���d_\�M�%�a�7��M��,e���g��KRcl{��*J��Ạ�$��=�F�d�Xdʛnr��yi��)Ͷ��|����h%��rHq؂�h�_1V)����ŶC�/o~U��د߹�Ξ�ʂeM�q!�W�R�L� w�����" �[�W�෕��"��ɥ�����u�� �Sl�1X�	�Z]�*�A#
?���s��B�=O�[�2��8҃�\����]��OԱ5j�L��KNӔ������$�
^%�;�H��}*��C��=Ϣ��ar*��@4ʜ͉Es�s��ɱaiwOk�T��x�QY�1M�	m�v���c43�L4ɠ�s�1HWQ�t�n����o�/��k8)�Kt�sĽ��$���b�R갇��I�A4N̮��B4x�F
^�R<eC~V[΂L�D�[;��@e���cl��o��/̅L+���"]I��0�cT�[����}�Yy20ͷ?��D���Y�����a&�)#�$�X	��l��\3��QJ�(��@:�z~zs���C�FV�)0�au��c�3VH�-�9�C�Y?�sV��Ȩ�˯Mi�t�m��6�-#8U�P��21bC'sr�ٔNhf��3���(�{�a�s�9���@�{�5Q��t������2R�u��k�;G2�����lR\�� �9@#�,7�����u�A��չ��0�*��Xu�ytj�F|��u[����k����P��� o᭼��@����m���ag��ɞ�{g�{�}�l¯���^+xV�!����2^3#�J���u4��(�tV�K��)К��J��f��	![P�Sj%��H�m����2����&ڶ���l+��p���ۅћ���u�U�%,ȥ��"ى'�d�,	:]@(#6͕1�+�n<�A	�+�I��_�_�j��wg-������q�:̭��L)�H��/9�Q�Ӵ.ӹ����htH���?�އ.�淥*z�%�ư�PS�A`�w �_�	��&��Ր��6*pK��q$�1��x�O&�w��p=m�[���+sI�!