��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\���V�fnvx��ÍG_;�ȅe�~�>���9�>��Y;�0G���O����W��	��	N<?9N:�KTd���Jw�*��>����*_�sj�n��2�|�7��i����L�A���Z�*n�T�����>3�/}�2t�݀I��T`DoGc�A�Rǎ�\p��B�%��3����6�p���7���VN8��@6����0�{d8J���~��y6.����&^�㞾�z����O��\�t�!Wm_ZYZ���gk�RQڮ^�����<rT)Z�jЊa0B��Ҽ���V��0K���Y,=�����3[W��Z�/��QhG=����o6-mhG�9�yy���SG:�X*��ż�"{�ԃ��8-��l8\��e��:��Y$PT�İ�w�1�XO!��Y\T���/<�x1�ndЍ �����ô�\�����x�߿ ek�j����}�չ��E�)�K�u�AX�� �U`R0#)<�?4�vf���a7y��`�6��嵦��vF�I����L�J����J�W����Fi�yObĠ@���̥֗�X�r�ya8�J���'��*���JZ֭�V��;�-����ܚ��a����.ُ�<���ӧDԩ)?��,�MWs�����8g/B���j8�����]tE�jE�6��G>� ��XkJ���qN���]OX$Y$g�HmQ�����/1^)%|=�g�ɸ���b�\�W������TS(�E�����&���%5�B�\q�~��C����Qv���:K�[?�ž�{*?Z�6��<B��g�e a!��6N+�L�J@:)_�d�a�l���)%��i{bv5�E�����Aw `�%a1	9u���]*#�*ט�}���\�����"d�����;��{PѰ��K�*H���������G�-XC�et!uݟ!��iWX�[$q��z��2JE*��Y ;�x�߃����a��9¼�3�� �O����ÉD���� �h+��\5eF�ڒ2q��֩�ī&�)�k:W=�p�P������`(��J�8�yD1�ã�]fG���}7h�=.r��%Xn��O� ���t�s�_�����'#�Q�a����Z����ɬe����떊�b'�����ә��W.�[��ק��+$�K�6�d[��L�\�#v=��*� 5�V�ǈrʙ>���K��l�����h&�h��⨼�nI�$cw��ɟ z��c�p���3�&�͗��$s�Z��<K���o�Sv���#:�s|�Q�|��1�Ɖ��C�&�-�[X&C�4�>�w��� �����G��;�A����R-�FRqJ���;����v{l�i=� �-|�6���Q�'�)$������
��i=ݒ{
ݕ�b�x�X���&_��)l�m(s>~�Bu��r�c�v�8�ﮟ�y{ҷ�x3ՙ�07	I:���2���1����3�U����e�%���fp��Nc<���G�Y�5�����v���@HA.�{r݈�O┥�ˊ�l�Տ8�+��6y�i;1>nЌ/0k�����	��m `��d�1 L+cO����F�gۥ[����#��s(r�V������2�h8 tZ�1�r)]�_�Dz�L��9�`J#=���~.��	�����M��?wci��-�,}���nS�ldq����<��y�E<���e��+���d@��#ya�n*�n�,�M�b��&G��#qm�_Gئ	�?�6bML��b\����Ȍ���|��?���u�XF��Chb@	��;�Dpb��n�ʖ7XY�"��|����P��O)�t!*����T�,b���"�j�M������17�m�Ha��M򶈙3�v
^n�� ��yʠ'��1���5�u@A�3\Ր`H�����m�bv��WM��?��ҭ�X��j���øA���X߈���$\�V��c�b�1 ���[\�c��Q!U�A�ڎuI<-����9��?qtЛl�b�Np_�Zx�_��u.%|�R�'7����_C�62�<�&g���(�Z�~V�E�&W�R>P�v
���qɻ�I{gQ������p��n��}�=n
�"�e�;D���~=m5NG�C�N���3���pn�O=��Q����>�>��I��U�>��Qg(����$t���3BW���-|e���qg�Xb�$���ӜjD��B&�E��$e�:�3���RT�O���}���)���	З�*�d��7/��w~)���	�|o	=UD�6�U�+w�xa�Ф�
�:� gn^l�(+��K�;�dq>p��M��y)�[��|�xB"~q[$���c`�I��{�x��rk��:3��W2-���o"#��{u2�:�B����g����R�x�c���w��ǹ�gvY��>O�J��XbA��� fY�[�t|d��u��B$���x���ƚ���%�>*u�	���=D��?�~��`F�6)@��`}T*v2+RnZ�%fks6��
��т���0S�>,�s��>e\�iX~!�	N��wy5�J1�>I�DA���^�����:[b+lE�iQ8�c�����G�:��n�����ɐ�l�����m��h&3t:���`�\v�N{��M�6�^1�^S� �<���v|���=$u��x��
�!x��#mq5WJ��=녾����V�b��"@��{��O�L*��@��a�k�<��WS$7�|�:ӕ��P壦Gg��P,� B����So������� .�.WJx�	?菰
i��z��7�ww|2�/R�����M�\��Y*4Q߮��i�0ߔ���tЍ\�2�LȺ4Z�"g).@'���m��ҡ���䫢	L���C�H���y%�!s�������ٲ@pd,���$v=+ ���KT�	��S�t����WK����[�x��*�_���h��;��^�?x������ 2/�t��Dj��@%��	����%/���8(�q ��Ƹ�a=,��e��yo!��ՏU_�}��.��(���Is�c�] �X&K��o�şx����}ituj�ns:�Xe�t�s�{bok�:ܣ�ʵDP��Hsj��f0��i�l�ytufY,ޤR>;�ů��pIɣ��X�L����ԅ�z�=�3�tPs�yQrw�n�x}�ߧb>�(�P�v�S��iF8�tu/l�w�9�+!C�5^;0������k�7�&G88�C�����M�χ���8�3D��-d,0&�����`}����b�s��赤�ݚ>�ÿ;����0\���2�㕌Z��׽}���(�������F���7��č:�O�9}�#�)�i�G2� 8�0���� �;��|���̶�/�ٌ�R鲂Ol��U�e>����A?�#Y̓�j2c�	������6�@m26�i�rrH7�����z؞�gd��?��#�'��C.� �������6��-���]_�e�t��i�G�A��د�l��4CQ%-��w	ߚO��1\���r̬��*�0����cV�O�&XiQr��[Ns�����=f�dҭ��j1��B��8=��Al�@���
bsڛ6Y`[�2�z9��Ѡ��3�@;˖���xM��=w�9q�,lF%�b���鼮eN�*/�hR�7�D����@�;�GP���cl�1��{+�;�e�570v�T&pZgʂ\L�֝�£1�v\'�Na��Q��+�O��C�y}�M-��wSL�"kA�܆5�� @g�`�Cea��?�1�S��-��V⟾^t���3�tR�
MWڭ�ʌ��(a�[	{��������}��F�;��#�3l��<�˭��kK- ���/�r��b;�ᠣOnP������ݦD�-k��ޯm��|OB.�?N*�˔ <����i!��ƪ"�nI.ۆ���Eo|���Wo0z�.���m8}�t�@E�ͩK �syF2���'b]�]ќ��Dv9����a��V�5�@/S9X�k���M/z�z~�]�,����9��k���s'+�=fF7<���Z��gz�zx�rA��JSδTuZ�\N���e�o�7a�t�[e ��?j�����o�!u�?Fp�v��'���g	�)��g�HD��P�\�_��z1�%:�˛�8GIO���;��QЕ����q�y,����p�E��!�2�h?� �EXţ��A�v���|ͫ�զC����+�8��z=V��2����7R��۬f�6h)uw��2����k`]��>�w:/����R�I�2n\�e{gkC����d�� ��4ΫԊ+٭�ϓ_�*�|��cI�:�?E��m�}Xε�2���
Q�aM[���g� �WXϰkӨ�О�:�5���(?F"￰�����=T�»~�qӵ`��Q�	����ꈾ��0*�.1��[�L�6����{L���4��̫E�r�0��r��<�O���ۘx�d|���˷L'��9�o6�Zl~�-7�&��+��QDh&�-�l�br7_��M�q�x�E�]��R�@5��Vh� :q3�U�+* ��(r��q��	��8��,=��aДL(��+>��M����s#zG�K�������z]#ɟs�Zs?�CU�j��5e~�Th�#�	�C��w�{��YQ��d0��D���~	NL��f�r��Yc�sH?1qo{�lP�_;�t�
,s�% 9�:x�S0�Cx|�aj��Y�"YV�N�X�Z��d�3 ղ������^������A��yK9w����f�~��Lc�Ż�-�K������CR��ˇR� �*�}���Bo�3� G���^{�����Ys�M,L��ƺ��0�liۅ�+�Ƙ,i�������5��%2�^��9gk�Z�,t�p)���h��D�Q�ؚ�W���N/&�l����M��S z���N���Zf~�_*���_.#��W}�����$�P�[v-��5Dm	��� �����9ѡְ�8==a���h~:���ǐxz��!Y�`-��v�J}���uV.��t�(ؘ��id|
��)�b�ǡQ�}��b�k�>���O�r_z�Vb�u"�e����~�����1K/R�_�R��DE����1��)ZIן�c2�oI��
L�*���%�g���V��_)�M{��,�`�]*�����.:�瓍����YJ2�&����Mbt�e[>�mo�T�	���w L�Q��V������]�]�/wrG�fG@����R�sna�T�}Y)�!�t���=���x?�Ӭn��P��o����>�%��S����'�i^�v"zO������N�rPO>E���c��{��������"|��*����w��K`/��`2�a��(�ó�D9��?��ѻ�=��~OR�ظ�:Ș$6��~��d���R_8��Ma�������d�8Ҿq��.0֖q}�=�g۞��/�FR6�������T���o��=�������a��~��B�{�	��o/����W1KJy��E�'
��^����h���T���Nt1�x�"�wU�=9����m��jg�6�~�q��63B�lR,D�H4g�{���ҝ�Q����s�(e/P��b���ŝOE�RQd�%.�@�\�K��0��N|���3v�	ӏ	��O�������|*�CFH�x��u� �i�r1g�K��6=^�``
���;�+��f??��@���A��|?:��V��ILo���cd���"Q���5�_9��?՜��i�x�Ph�Q�`K1yq���ݞDG��^�M~���9�Z��~�m��hd�̼/�)���q1~�r��;3B^�~�Y���M�4�.���c�8A�Q��Ɲ���bXf�T���{��87h�LA-(C��\�b9Y]դ�.j�@���ʭ_�A~78��,��������U���Ԭ��0�}��(֕�X0х����SQU�o���l��e�����4�>�,��:y�����W~��՗�5@�/�8�Xθمzi��#n���SJ�`�%Ngƃ#�#�����~ũ\��ޫ+uxҠ��[������*�5��'��A���^�HL�ƙ�$�?�k_m�	J^ʲw?
u�/�I�}�=�]7����L���hC�<���(O?]�j��:, o�ndo��W� q���;54�H(�����eU5h�+!���]�W�6��R�6~���S����+�~ԬR�Q�̓�R��W#�E��SB�\��=��@�����OD҄�U����yþ�P0*�� �-?$�>�:e���u)���l���m0�r"�*��\�+z���=XQ]��`�� C�%|Y�(��2�"ج�B�{���pÝ�IW��tn��7Y�t�H�3��
8m��`�A���q:��{rC�O�R�-+wJ���yH[NAw.�s�e��ND��4}�n�Hq3�${�q��.����s���N��^?���	/����|����1�f��'
:)�R�bR���S9�x�Ѐ�y�<V��4}짏��$5#[��η붱OHB%��=Wk�c����N��>� �(h�:ԋ�dJ�KHw�I=��[��@�d�e=*+ݹ��H�������;s�,�Ŧ��MSZY��/K7�?���D`B[����I�A�=��^g�`����砓W���1UΤ����Fa�٧�WT �Ɗ�q����VV�t�v\m�Ak/p[�g4�FU5i���|��Ø�N 	��8��jԵ��b�<��N<���X�s�պJ,��^A"�D��OƔwN�9rn�\�&�G�7�� ���z q"D�H�����K�~�l۞�N'�����T��G|5#�"	zTs�H�a�M&+�����ɕ�	�`�Ћ=F��zhس	��6�B˯�Y8ұ���@�i=ِ��A^乩 ;�Q���"yIt٠Hj4�o���|<��Z_��c�����|�q�>y}��uB��۪B̈3��u��_Q��w�;���&ڛ_N��{{<	O�+��eE��6�ә�)�f�j�J�td�/�Pqj�E�dX�m��#���A;�Bf1�v�Do*c3=�k ��w²nل�ig`r����U�B�@֎Up�v�A��K�?&�
�Jw�rִ��3�L끓8�T>��[�8��z'�CC-߃Œ��v�WL.�+�do���3{D��P��HR�7�	lvH@��}�h?����m��7x�7�'LW�9���ь�q]�p�	�{�gѪ �����r�[��T���|��� q��m��L �C��54	U�v�+1���G'o>qݑ�����M)n��w�[�Vπ�Q�.�8��ưc��Q(r�/����Mr$�T��ʪ������Z`��(my5���\�Ɓ;�]��d�[{-�4=�C�ڨΡjZ�:�F�������i�@N\�@�k8�~6�����xe��-4��S����a9;t�ﾗ[�#߳3�7wyf ��ʰG�dJ=[�XQC�*�'Y�'��Z ���+�����Gx�eHmm�uh�iL�d� �~V�Q����:no�мfы� '��G�p�'�[J@��IDP,��-��᎝����|ˀM�{v�Շg"1w�S��%z}۲�6��tᅲ��ġU~�����'䱽�f��Q��
畮�,����U���'s2K�ݕ8�tR4��?%�v� (�ҩ ��<�1��c0C���#���	���z�����]&--�ZW"�l���/�������I����c��XW�0=XgumC��֭]_w���S�<ߢ�6|��8�埴)6�Gr�f5���I_�D�����L�5~0��N�f�(����?6	y]��+�+n�����w��"N�z�Y4Q���՞6x��09���ܞ���W���22��4��u�I����z�^n���]����A��W�Ź�ʽ*�((�K��D��6�ʑ��E�efN4L�3Y��D�#^�D��a�ާ�4GuZ!xF't�:!Ǹ��s��/,x1hA��H(I�+c\[ ɟ������8w���Fz�q�5��^�Q�/{����������]��?������%hE��Yt�8���3�4 i�h#|�cmJ�͞%ڗ)/���K�MO����ۼ1q9�bc?G��D8xE��`��-�I�R���i������>��C���_ǆ
��NVH�����s�r��cb����%사KB�8�#�4X������D�I[��sw