��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\���V�fnvx��ÍG_;�ȅe�~�>���9�>��Y;�0G�CZ3��=�����#�?2��f=8�*k�n
h$��P�
g�&m�?��eAJ0UM��缟ٿy��7���x�:Ӡ���a��_%F��K9�'S-+=Y�<{���u�W���l�ɸRJ���g'�vj.>���,Շ ��Wd���v�P�`{��4�G&��`�}j���蟰#KP�M�-�ϲ��\��Vr]	�䄤Bt�� ^n�����06s`���w�������O����׃e2�\_D���V��ǲ,~�aE��(�q�A5В�}���e �I�����80�yU��y���2��9���⫊x��$U���ė���b�Ƙ�9WSA3~|pf��Wf�8���М����(F�����ϡ*>h��</��r��Pz\dK!�Ѹ�ː��[C�{����tu�z����:�������Y��`�������lf���g�XX?[T����آĂ���GG�pʆ�B�*�WρP�w��W7a,'��P����qܙ�/�QIC�πΓW[�������>!)����uP$�A��q ��NF���l7���X�~_�U�F+���\���:�fu���
�.��m��0��
M�k���{Md;j��s����=�y��O N-�^13�
,W�6�;������H�����i�O�i��G���.5Ո��]���m������!�����H�߫�N[xr)s2p�Qi�iEC�V��*�>���0٬����ur4�)����x!�ZKk�v�#�АV��k4/��5�
?�:(�C�}�!�Xcu	�\�y��0��Jy��1'�0��i�w���Ԣ:>r��E���̟<vm�oJ�(B��~�\���2�a�Z�J\���&�|8������N�u�l�w4¼�+�|睎$�1~�4��1�*w����d�w�o:o��?@{��;�ߐv[Y��l�Nu�ذ�=���\|��X��n�#D'De,*I|�W[$|�^u9���S��I�тP0�4�2�� 1�P��w<b���ğk-�~�"��+��`(�E�Mfr�1�E�)��T��ǎHD
�?��e'�j�*Kd琟 �Shi�W@$�w�qя���qN�Y��t��愯qO�T���u��z�N���8=�TG1�#ُ���S+�8��x���N�|Y�XL�簪�K_��2��EmG� �dނ٘��(q�Yb�NQ�LcT}�Q��,�
���R��Soŉ]eS�0�U2�9K
y�Ȑ$zS/;��]J��J���	��������8�Qsڕ�3e�?+T{J[��WlU\��_�b���1������٨��6�l�!�Dg��/����P�Pi͊�v��冶��B���������}�i}�R�m����`VZ�D��ي��>6��V| a���!��?�d�xP�!��R������e9�:�ک,���j�k���f>�F�l���k��*R�|����yJ{�h|?bZ���!�hH�� �� E��l쟐T$�g������ȉ�B�k����o�^œ =���
�mC%����CH��Qq ��|�po���ۻ�m��>b�y=|�u�5>��Q���)��O�������x�j�w�A�,���M�B}�����������lTc��<�I.��A�a�S���d�kO�x���Β �z��c<T��û֛�rI�rH=/��6eI�� D�C�uh�Ç����>B8���=����CB.`#V�hٺD�YO��ZwiX���,���e�0(�	�f1���g�����/�N�� ��W�Kt�mTz�e��r.[�HA��^M�ZH���y��B��� �F���PMe6j%�Ӷ��
z7���}p4����ث���%�Wa�j�vX��@���nW�B<sE��hGP��+\���s��oB"�2
2�
<��}���7�Ur�Q�G�۵��|@E��B�
�t~����ZuR��o:�ˆ������`�Oɕn���T��%�Su��J�'�e{M�R�N�t���y23gF��z�'1"�Y�,tMN��a��x�1��J�6��[�t�썃��HV<�>|܌�K9_a��|�W^|�D&a�����U���W��1��*o'�"��I��
���Ie��`ͺ)b����Ϟ��>u�WJ�h�.� �\9�ɼ��Ł]z���q�Lvl�TU~�+ �<��Sz�AhE!6vB� 4����x�������7]�*S�OH%�èf?M���1���߇�g��C}wKYȴ�f�Cg�zrzb����\���u�ݧ��|H�qY���u�����]Rn�����f���'��R
�b'I����f�8�^�#t��#o?Ԍ[��&Ξ�o�[@�
a,��-����/W�3��|k��8��U�ӻ�7�RVf�f������\���h��ê�~ə[��.LG�f���n��3��|b{�E~��PI��8��x�5����h/�`�.餳\�nd� ˸"f,�dy�"���WYe�S��ׅ^y��>�1���'j0N�B9M�=�/C)��X7.�}d[5|06��~V;���6w3��wM$��X��J(�E��g `�4Kd-�
<�ɒ��M�F�ir֡c}���B�������h��t���=�޸��sK�������sE!Z�Yǟ�J�W�?�@��_k8/r.�H�o�|T�ۧ4^�OW����z���nr�)��S(2���^����1,��`�A�J��c�ʕ�O��9�&`����Jz�m�m�F=��gM��!J��NAp�e�' i���~Y����%!�fd^�c>f�o�f���������87C��rO�����;��2p>���)g*V���v@�9�q�W5�G�>^�m)����K�W�u���Yh��)�����kUZL�`9�5�-	c���CsAL��9���Yϑ{��U*���L�F��������+A)64�""G���R���(�c��|J�����)�����u},H�ut�f C�5��)�,���|^=>��˵ա)UPǪ��h?�p,�r���U
;]Cp�R��ta'�M��D|�NI��(���6�CJ����})��c՚a��RI�����|��yb�`��f�/�%��)�>��7��B!
�bV5Ӹ=����;�	S���v�A�.��)Kg�3SD�@���j:b�<Ӯ Pd�k� ۬h�*�����FN1�S�+��(�M�O���J!��vL)U��@�%�OI/�^w��lg���7歏� ��Fʳ05�,�)a��m�rR�FO��,R����pb�7ٰZ��S�z��su!^�9 `�d��P�dè6��P��
"�݃��cM�d�R��5�����l�@�(o6�UQ��]4�̜ޘ'�����<J����H���9t����p�0>����B����B�&Ùc�Ͼ�
��X���ץY��-N��-�K3t՛^��K�ި���7	a����yJ�vf�][���>�4g�Ď,�6��+���ѫ�f�Df�V�m��v��q#�N �^����[�!��A�ߍ�&�o!s��TZ�����:��E�,�g���-�����*�8����$�.��	<`��Ƃ���û����o�φ��,8�v�)�[�,��+<�Y|���~�S���0�A�jz�+I2�+(�m��� ׻t[g�p=}���!&S �)��PW��L_��s�i.1��"zNG��<D���:p�����;a�g�F��m� l�N왭��4-;�h��n�)��4��Ӵ߻R�JJ�S7�h1&>&8} sp��P��ގ���ZbǬ���f_D��;1Q]�����Ş�9*�ږ�5�X문J��$(��� � ^ċ����4��:�,�Y��4m8��u���M��R��D-@���и�A��p���O��#�|7�ڧ/N�elQ�B/�p9Rɮ���*
F����`	���""��[�b��½%De.��>��T�Z�ĸ|�z{D�����1�f���ŭ4|Q�+!t7�#��p��:��'��4�ZM�3H=bq�B��4}��Tp?�	�^_���s2���ר `�v��4B&	_^�T��~<�^̊�S
������K:�%���/��p�@����T�fT�"�>(v*&���X�6�_�ʚD]�� ���S3�+�ەqW.Y	�kf'���Ƹ~el0�Q�\&�c��1s� 8����"�e[�W����+0��A�n&���=�:ɹ����0n�˨�*4 F-���J�XD���^��C�Y�u;0���L��^l�@v�p����},~�z��Cϡ#l��3�B�����M��țz���޹0���l���J��^��-�G�C����I�_�����T�v��%2Τ8Z6��nŞI��*�����c�M��D0_J~����Oy�W���W�ޒaL|�4�_a�OH�d�@0�4古����&������z�uNB��'(����3Sjlc��,g���N_�D�T��!��`��S9�ie�P�m]��Y)NQeE����ٱ<�h,k��yi���<�b�<�ǹ�&�F{��h�r���ܶ�i[�g�(2�9_��X�UfC>��HϗA�
�=L�]�4١���e��N�ڝ@�(�����W�Dp'��p��4�/��85����)��ȝ���1�Ɔ�l�����Ă{1�oW���{N�0��}�g��u�7b��˔u=^4������~����O)��.=z�+�ۙ��O��.�|�ł0c��6'���(�U%�����o�{�9Z�ۨ��Ì�_���wK��I�M>� �W�T�P؄��J��?<O���@#�Y��I$~ �	&:�!#	R	A� V�jԞ�Y��?G��<��>;"b�Z��?1?O����cl%�E� ��eb ��������v��t4�ڌ��>����Ot���;�����_Ǭ֏�	l��-kK�9�T��G�J�O��M�]U�h5��Ts㑘�TQ�o�_i�}J��7e;#<F:�m�I'*�ix�ֲ�mx�\ƣ�?������T���b����L�jpf�y��u�	�;�>���~�<у�pd�O�8��F<Q�L��q��o|ԄO�1���o��'��u�2{i7涷��>�f�9���o=��a�#վ��Q��T:q��$F�؋.
��*��a����L;3�Zp+�| �MV��c@�f|�B�/��r5[���9�]V9z�Qk�K ��?E��C�������k���`�jo�7��w���O$�Ȁ�)��'�"�$�%�C�V��t%�S���	�0���M��q�r���i���͊���8��w��@I7�FA����K����A�ka0��+�(�1R㞵�L1�~Ӌ[}]ȫ�A]_��-�\n���޽/_jI���:J_�;�1����D�(\��^<����)t���D�V�	��5���>B$�J��͜FJ�ޅCСzAl��e;p̧�w��Z���,oc2��6�G��5ڇ�����(�^����jB\�BFb���������rkޥv�y�X��(�.�3r��p���0��h�͡�k��F����[4��z���vg��豍C�(��Y��1k��>%��h�4������'��8�H9�ZR�Sf~���3Ӥ��*;�8£Kj���ڔp7���1��rn!�i���e L�r�ꌈ�����*�~�p�Y3�¾�.�����#a�zςi*�u��#]x�hnTa��:��9�7_����G����2j2HY��ae���z�����S<PS��ש�
ʭ��J͘^l�w�3&o���+�_6q\�Z�̈��m�I������5h/7�Oؐ=�+	��cV��%�8�ŧ�Oū�1]��b���P��'K�G��X����v��6�@��əu�!D$+{�7����|��gW�����s�M��x��Q��m)�
��'?K\�9���>�EU��lBj)lo�s�+��X��TMetm���͉��\��
~zr-�1����k�ʻ���G��I:T�0H���܆
����B�$<����1���o��!�*˸�	'E�cf�ʡ������ψE��x��RX�lT���8F��Zf�)���`|�bP����'���llj��{��օRU[��Ԙw6�=���}=5��ڥ���D��F�ό�^��lM���բ�4˵��2S\1�op�Ya��^b����$�5t1g;������=N_d_��_/i���k<0��� �*b��tS��^�>W�C q#��w���-�0��=�%t�Y,��x1W��)$�;�W�5�����_h��[ QP־�0���È"
�؋4 ��ݢE�lVb��@�0M�tSP�xK��ss�Di-��5�c1��IG��X�� -$���-%v�:�7����=���o�1?囑�0x���W��C�+4�J�1MNEcp��?'�g��֎ګ(,N{f_�B�`��TӐ�C�4/�Z������4��Q��P���gc���-!E�fD:��&ע=��᭕��Ǜ�0M�7�e�Xs�4��N�\�����a�H�?9B���?� �N19T��R󺘄��&�����E�h�F`�"�@���D�~9J��l5��ΥJm`�����&���5���ƽ��k%���������seg/=�\0ہ�� ��L��Q��bRfG�Ǖ{�kBC�ꛏ�� ^�Ah�X֍�T��g���� �|��t��>o�~�~`"
�C��f������ ����Ԇ>�
��W�ޞ�@�3��:UJ��GN���e�k�_F�Gw�*i��^v](�$%��1��cV�`�8qT�(���b�~X�9�̖T��N9I�H�-޵ ��i4� b�sd���?�пav�=���tf�E�^	S��~2�&�yC����n�m5��6��­S�E�;66��ɵ'�T��7瀡�	�r|{��ˁ�!+���R,>VP��L�Vt �3@��qw%#|��F�sVc f��.�*	�T,J���e��Iz�ALܬ^��4����<l��"T��Uʴq��奐�,��!�2n^]�?�\l�\����y�L1��l�g����?Ԣ��4؂]ŗK�$�*Ksei�|���1!�H`2��Ka��uV
? 6����)�ĕ�&�L��h��H֖�A(�fxM�Ϥ,=G۽��3�f��*'s�r��
ɱ®R�T�(Z E	�a����������>�@��[f���K�L��
�q����`���r��<�t��@�������e�@��~X��[� !~�,w�HP�4q���:�$��K��T:M��;?�Sҝ�����;�*�hS�'���N��}��tM��K�GB�fpݽ�R���e�8�7�'����&S�V��A����+'Ϸ�W�U(,ay���|/"��'.�4&U@=�b��yw�Y��T%h���h
� �x�T��\^���'�F5�:0sQȬ?OO$�zq���s�����or`&z}���-�ێo��!C˒�)��
Q`_�ו]��I.K	���$�O$�Q���]^���uJp˖�s�ꠡ���4���P��B x�Q�ߢ���M�X$!sz�
5��_���4��t��d%����b��-,�~��:T�����	�{#m��}�h�$6T&��b��8|͇hz`�(����G��O�M��%���b��:�X��~Cha�M�ל��c�o%z�E<�bʆrg�[���izE�A�	�>B�9����0�А�<�hǐWSD�����r?��j�|�##l��'IVb�6/�O �z�����}��_ůVv���i�?=/J��,T��s;�iF#@�6v����*@uz�E��Y�V���q~nh:�Xk���W^�8?2a9�w+ZǊ"PK��(?Y(�(�����c$�	��ק�Bܒz@�g� �۝@��� ���&�e���1�ܙ��`�7���_?-M�@���qp0s<��$0?�Hɓ<��Ez��%߫�^���.�J�'$9��[��g��'�Yx����>�v�W�q�g1�uC;�:����
2�3��/���J��av�u����~��"��ܵk���� �L�ۆg',j6�4�[�u[ئg"��`�ZΕ>r�O��PM>�Dw���mR��G�>��M
繑oI)�.���
��E(H��o>�L�!ֳ�Vʊ(H�O<`K|�q��p0��p��J�ڿ�m9�I�jK4)�gUR�s�v�'�����S�hXބq�|��Gm�?�!Q拣;�S�xm������Fqw޲)������������w����T'm}Nyu|VрQ�nb�&������r�̈�3��O�6{1\8C���ɥ�iM�f�e^vu�J�!��&�?/v�m|��Gi������y�N��bxE״��Щ��A�����nI6�r���#e�]��wi���=l�ǻ띮�掌�X�6�u�҉Ēz,�ټ�W���F��e���fzWY��s�B��jY �Q�tG��u>vt�}��m_C��wE�=
 �4��7�W��c�T�O���/��_�"E���s�� ��q�x���Ӯ��(ٓ�T��En���[޷�`旧��
d�d�+ ��r��?��=Ht_�b��u5��Q��[0�Qv	�N1JZ�'i���#{F��r�n�����U�4��|ۯ�^�&�B��:�oM{EflK�4]o�����Z�g�F^��V��[߲��а��7�M��� �_��iqS�@q��5��Q���6��������@I8�ҐV��'g<�vȤ{�@z	�Q�CrN��x�;��'eV�\:g\��ʙ�iclf�Z�ӻ߿�u�%c}٨^@��'��"�O�+
o��Z�!������Si��m|�4B�ʺ��
���f�Il����J���<�'˝���q�bg���K���N�
/>�*�-ܐ����<����RI�?\���bzb�(��XWo����M
����g�&�j�!%3#m��,9Z����<�h�w@(%��d�ё�1���cE��[N5i���d�`rZ�:��33Y$�$��B�f*�ݬI��9\AӰE�*�X%W�D�/H�ٌ�����	�< (�\�Iu?޻o
<����'8s�[��;R?�>*��am�p!��6���C��\��O�����l;��]H/��7'_�ɥ��%���41���ry�/�;z��D��m(����Ui*Roj��G%$R&�=�F��
��by�5K?�y?p���" )\�sm��Lm�M*�4*UT����o}�xsB���\N�m� 
|fh����0le�/'"~Jڞ-'�z:in��>��88P��\W�n6l���,�� ��Ҟ�����Q���	��
f#����48��S�-&gY���m�>�7w7{��0pS�S������#�
f
wJI�ױ~#� ���P��DFȯ�~ZmM�.�<ⶻ4��2���ۉ�ݝ�`�
{a, T�}oJ��*f��9!u2Z8��P�x~��)��f]�?��ȍ֢ܲ����cbO٬�Ǔ9��G'J-~!W;�a����3�'K��"����.���+��)(�"ׄw��ذ������P���Ydi&ǟ��f�.�,Z@g�d6]8/C-Y')�Xk�^>���#}��s�>�66�O�(�sVI�iro�幸��Z������T7|;���vV���UXk��k�}�W��ʧ��J͚1���m��;Qk��.�n��G�C!�S�񧭾Z"OˌYab7>�<�>�����3��J����2�}�4�+�Y��N�Q@4�Z�b*��
;�FV���+ޝ�~
��ǽ9��Øs��Q}`4�/U�Љ@�Z䲐H_W�~����Ftm5os_]��䢒l��-'F�)�Yo��k�Gd��9�A��㌧����� �c������X5rX�Iu��C>����XT\��)�f��%���M�nKI����I�琫�a-�
�C���W8P �D@�~�f�Fi�kڡ����\E�"\�!a�1���d�~v���� �o�L֩3�������u���q	�E�K���b��������G�	�����޵޶E_E��{�S��Q�gO��1\�o�Y�(ux*����DL�hm��	}��������>��1z=�1P��@�z��J�|�=�^����k�<K�K˽��jq��}��1�e��B�
䝢�T���x�P�s5H���.?�WY�J�ѕ�L�%�-�.T���Z֐E]<�t�q>�2w��̠#Հ�����&%�YO���)�P�Y�EO�/����R�T6Ch��z[��������������~ڤaʀ3ulK��Z�Yឧ=iWs?X+����B)�;J����gS,�dɰ��Z�B7�W�%S'��ŏt�H瀳Ӹ���A��Ә�km��Y�.w0�-X+�,o{�T�
���3�����8Q���GlPU�K�L�)١�J�o&���@ue��a�G�m��1�	�>G7�/�Q�HЋoI���<�Vn����.�-���U*r�;���Ո|Ҍ��$�����c=qDk�bn�3�*o� �]-vl�Q�#`�@�MR��Tx��ǧ;1K&�	Z�'�8�����7�_	h�(NY4�4���[ٹ5���K����0\��emW뒬%���S��5��6��pv=.:�M������(�ƊĹ%\xCzz�Ȏ���jo�{	����W�����B]JE(�x�G��r24(y����y�,T���c���s��W��}�[�?�S��m�K��vf{�8����*�	 �]O���6*�0&iK���1 �5�B�>��d�K�8�Z���#a������ ��p��6��#(c[=��B7��7��Τ�9�a|i(�2K�4�E��R꜄�4������'U�z�2K?�|e��_D�,�؆/o��	=}|=^�J�w�-�]�A!�|-M�%���M ����YD�d�����|���E��7��h��&P|2�;=v�k^O��L谾�nYF�<�x�y Z��o�M��v�!0�\��p�B~�B�v&{�������/�<ElURA��$Ǹa�84Aڢ�~�!*���.@,�\hW�������iH�#����q�X�G;���N_�`�4?w��@����_��1#�	|�/ OP��@�f��X���X��>��G�WB]�����*=���ldT��Xz�uccw�1 5��i��";��hu�ͪQ��x�`���yſF��/���f�c����q�Hr�v��U'��')׻��0���Η3孉;�����X���G�w��C�D�����k{ǭ�5Y�D#���2����ih��Y���J��k��O��	�UǦz�L-��� �2�F��E��cM^ ��y~��>��X����XT�/��a����������N���g��|�݆4����N-5%9�����+�NrL�a�o�1���4������? E�6
�WjE?��?����0����(G�p��H��FL՟���;R+�0#|f�ʊ��y�q4�P��c4�>E2��Ufl��D�]�����+AN*5f���Q����]�姶�`��DD�SRX�c���雑/\h��Z���pqLz]|�iCTn���<;׭�B�l�#:�p��Ɖ ��y��+%� �PN:���?1��&2��������沔�+��nTp˯ٙW�H����.�p22y����Qw}�x���V۝UR����):O�#�������Q�{�F�9T���^�3O����_�J���L�	\e�Rlu�#�m�J]��m��op�X yk�J|NI�_ڰ[�_j5 ��Pai���>Ł��l���zCۅi�wx��;������Ϊ^��HHvr`_4��}:. Jd֪��n$�x�.MUG]�VQ!�.�`�$}ծ�'�DV��s���}R2�!6:�kĭ���<�{W�� ����M��`���f�5qV$��l�O`y����S?�������f�a�3���T�z�H�s*��\��o�g����\�aNZ{�ި�B{U�	¯4�)�Q�'N��Te���!�⹵��l�4���c�wUN�r�����x��Ē�t^��]}���?�g���� �w�{�o���CJ��n�P/%�������Mݘ���]Φ^1"Z�nqpk�0rw�5�!Kv��w� �J�|�Yg�'K)[�@X�[U�៲�w
�yQI�96m�ou���v�Y�I�BO���ÄTs�2�̫s �����V��k.DP���1=5y������'޻]�*,�H��Ol�*Vk��k��@DXg�45�PR:"�1#c�gOžg����r�p8��m��J�3��>
�<�g|N�!��z�A[\�[���$Y��A�<h��e"R��O��8'3z��`���j�ֶ�#>�=
<܋$��\B\_/�v����t��� (���!�/9��
�3H(�5�;�P/�B��$�����i���
~��6�xߩ6^t��z�\�
��0{�~<(���$T ��?뺩L�?xz�dcsF�W��H���k�þ�]�� H14*I̬�XV���e��3Q�\K깓@���̈`�%����X�6�Fu�A��<�eO���jI����P�}�9{s���/��H�đ^��:}��&h���>h&��h��pn=�#޲���r������Z=�/W�M��`}<(�U��F`��uC�������4��/�vE&��񍥊�"���6]���V%�kv�kM���^��OEl��{d/�O�3��S���7��C��{��g^ l��ƶU�jl�d���Эr�w{�k��h[��Jǫ+�����uU��DfT�6���BK��3��|@8��6T�X]��W�@9��������&p�Z�M�W;G
��iN��tU\#*2�c�ϑHj` �J��ǎ4:�S<J��UEi���V�!J]rcl�TRL`d��|D#GO�\~!�������zh�R�V���k��!
q���yD^�3�h�Gp���a|c]�q�i���vT<�3���Xl`-Z?�"��&��(�Y���%UGQ~�(���m�ʼ2/�W�(�1}8�ܱ�fї`��B�x�/�����,{���k��'!� hPk��Y��N�c_;/��-*�]�T��?���2Q�|b9	�ѣ9�	��Q9A	!���v~T��w�X-UT����V�fܟ��Й�*>l�|��`���+a6�ag���3��LS)���.O?���y�qFo��Q���+���(�6p+��zJ-�L5ؑs����'���\�Q��(Q�3��1��{I���Ps��@󧛊��9��I�C�}���n�!��O��j͢Ϳ��[	]