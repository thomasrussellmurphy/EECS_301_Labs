��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|̪��q[�dswؔi޷l��0��`�K��,��6����i��Z����FՁ8u%�S�9oټW�Q�C`-G��h�Z$R(t��u��
K��Y�l�uG;��g$�,5�<V��۲ ���{����s�y�q�!Wf�$�z�.�
,`9�;���s͈u�t�(�����дR��9�K��s�q�*����$�\� o�����N��W�h��q�\m�͔�u��fz���T��O�h#��q�"��'$o�:|�!u�z�f���C�L��V���/[b�;���5ϣF�g������L�!]7�~�rB.����??��i���z/��˧�ό��g��Or�Y3�Ng�Ӂ�s2���ö���1�G��~��ʧd"��:��|6RӘ3F0�n|��q�eALf�˸zu*���)x�,��So��؂��.�,Uٙ>���Y�9���\N�,��� �)On�5m&�b��=.�>�Ő
��O8�
�1�z�+v�N�/�F2�k)�A�d�Wb�\4fE<6���#�X�{� ��Т�#�ɯ�n/N�
���[�&���Wyfyˠ��Y}����rg���GJ���@\�Ejp���	 �����@Y�c8�-�y`.S#9,Q�}Ǣ���5[��#�2�����n��^��UbY�"�[/n�4��Y��Z@� �<6787�7������6?m�6툂��\]4�x���3�hn&I���7�ߺmފ�/�y�jFF��C(|�{G�����{�s��G�_�1gVH_}�ٗ!��X����r��B�ԡnW�O�Re즓�A�t�{��f��HѦ�Vb�փ�
t��&��QB��Ē��ẑ�;2� 8�%%!fIK"��� �hQ�k~,��˲��0?�m�9�%Tp
��X�P���"��"� ���2�a�f�7&#�������JڹO��'�iւ2|1�>Iin-s�Q��p���鎦�˻B���\��ŐX�/ە�8��b.���	a�VD�]={�^�y@��=��ܓ�&�#h[jΩ%�´�aoH��7h������\��-�n��X�	v�����+M)�P�`h��ꔒ�ؗ�Դf�zmiݸ���=a �gHiy�f���iH�EW0�r��~r��֭ކE7��}0y�rc2}KD�m���.'�ԯc��D�$\{\�d֌̸A�3@kw�-����b���,������k�S�Ũ��t�TX���{�H 3R�����.N��xA��������+/��+#�C��!��Tw[¥��@��)9V�gr��I��8p�ˤ�'v⚼)�Y�q��vo���J�L�5?R4��g�R��d��Zs�H]��+_�ڱ�S�lc��mFi�OG~�!N���1[�X�o�V'8�;���~bK���N�|�j��M�����!QG˓����Y������8��G$�i���-�4"+q���ڔl�F�ϪH����W��O&S�'4���pIΛÉz(�r��|3w�w>��\��{�v�s2�i)D�59VTy���������,^��OW����!nF{j��ڪ��Bu��{}�+����&'���g^U��4���m�*�38�B�U35 ��p8�!Q�>9��&t��A�%���@QO���R�7M�jk�U"7*^��詿��9i�:8Fk��H�H�OTH���=d��)۟���A�s/7�LW����/78�_f�b��ţ�̾`�ʮ��%Z}ph�b�;��mQI�ׅ<ͣ��	W<�nsO9RL�|CT'%�����s�����QFYn`f�~��N�`����!5}���ڊADU���]2�'���q�r��ޞ.z�J�%�/��m1��ˋ��du�����/4�iqI�A��+>�H!�@O�da�4B�e?�Bc�h<J�$n���0�
����A`��E�Z:�� �F����-0�R#��FE�#\�����|Y��V5NMl�+��)��&km��7'�
vJ��sk��_	8X���˪ըXY	گ08�������V�@R�[��,�����r�Cr���tnRWnj����
�Fb�~;1LWN��/��Ϯ}pһ\���;�D@�`̊�X�y�s@�_�f��E��_'+4p�ȌY���Cv��8�8�b\ƅ.qic(��Q���ĮF_��?RC�p=�Z�rֈBU�(���S؂����rXe��"&_�MGGt=�~��j骹��8̎�j����s�  ��.^Q�����Xp�O��=��4��-���<��5�0��DW��/{x]!��^H�_���G��MT�+�rv-�N�ϲ�XKJ��փR�PXg'��B5��>�+W�����q��6YV��i����=9U�OF6��A������1)�	�E݅����I�C��;�ܳѻ�	yq�w�����xr�n�9�y�^Lڤ�1�~�%��������4o�T�h�eT�~��|!k��wa�c9���y�#M���sE����P�3<�W���!�~eHG�� �f�+:'���2��	sP�|�ŕ�$w�>`�붲q���Ib�і=�pۭ *�� �p1��
Dd�\e^�b7�����9�Y�lJvb�p�;���!��l@�����;L�N�X+PZ�T�*+��Ԁ�Ю�uɧ��άY�S(�.`aSi,k��J��ӟ.m/Z�Ў�3���m��5�ibjv�u	8�~�L`�������m���:p�;����*Mƌ�/�(Tf|"t~E�m��Yҕ��^� M��!�kE�J��P�^#��V�ړ���a��y|����F��vO��4��%��^��U�����w
����?�������Ʉ>u��/�HVQ��(��r�;*��UK$e}v�S�L��x�r]Y}�|��O���.;n�&##�����G[��){�FGTRO]�j�nY]�.��>�B�T5�X�Cz6y*�3�|��E����J�����̇'�\��8��:���w���?�д��h��k�9��+����r���K�1P��،�������$ߑ��i��]�Y������G�S|l�����b#~Idk�`���:�8]�y�5�7��fX��ݴRU��T|������p.�v��;�?���jZ�\�J��7�?�M�>�o�C���,����,lX�+�y���L;���L���]��c�o<z�Q*S�<�꼈g��h����=�㡰�ۉ��جz�^�C��k돴0�br�PGJ��Ly7Y3w��K��v���t�8ZY�\eG�{!�ؓ�8`�oں=�d�nQ����C���5b儴ɉ����NW�d1m�>�3�jP�g����^=���7k�1���`{z��n7^�jGF��=D);��X'��#ȳ��,�<��n�%�j/e}�� ��
{����K���{j��Ȫ�^ȏ��D��j��,��^�*�v��FtD���Bkz�I�£��?�|�����2��������E0�$!�1��<M�wi/��ߝ�s�a`i��oD`
�o���`�����QBB-#�G��ۺA�\�bW�+�N/�������z����I0�N����U�`�gʯ��Ai��7[^��z���5��h�_ĀK{�'(�����II��B��H�~�eNh1��.��	���V��i���e
6a�Y�f�S5d�q�rl��y��`�J�ʉ!�������)NX��ޚ�w���y �P0|S����"���/2�UoOGz��_"��E==�0���y����vTr6p߇9�6BV�+�Fm6L��%芠�ׇ���$�1x�u��H~V�J�%��#58�tY�Mֹ������_~	�L� ���A�T��Ж }O�v| 8�/�:�{��>��-�mv���+���:��K�D�z�t�7A{�gs)��W�M�9$���d�1;�N��`�)���D�k0or��x�]�i>���$r*��f,�������B�����u��c��E�OcPn$�@���c���S)�~�������0W5�
T�g�!B���kGf��%�<��*l�(�@�/p�F���bUS+Q`x\_n���Y��覮hVo��$?e0��q?V�V!p��"���o�X���Z*r�V?�W�����6�C�s�+�Tm,V�-�H-,�:+����VY�%�ƩNg�o����>�%5�
�'(O�ӡ-�'�y	2��#�X�����se�,T�t
���S\c�ө�#r�c*���A��(�OkeL��p3h���!���os��*s���g�]o2���ԝ�jQ�d�Ni�L40M�)L��>��3��@'�2Ư�k��(!\��!}:�u[y��JgT�w�7O�G��n����r��,Ǝ�I;��vC�f����Zǥ\����!�*��8���H�ߓ`U���pGD��P;v��M佦��Rig7�F+�\�9ti����~�u@`֬g\=а7;� ��N�N$��b�Ê�����Я�I��L�םXzBC��b�aUH6���p��浲�01�"
�CvB��a4bQ����L�\���|�w2-�ސ4�Z��"�
\g�u�X,)"�3�����}���c;y��B(���=k,��%�vb�s�n`L��0p���g�Y��E-'ٶ�
Y�2��t�4��i�դ_|�>�{��" ���J�3<�i�W�"s;/[R��|�h�g,_~k��Q��ʺc5�]BT��d��b��VDI?�N�{M�$�
i!#�M�kZ�����ה��\r��fW��Ya�J����.��S!Ժ8�a�9P�W��Kxn	�E9U�7�|��MA�P������R�z��(2tX~,��wZ����扥t��5f$Ƥ�y�b!0ɏg�$�0�'І-uU���a�|�9�M��R_�^�]�`΅�.�������5ȹ�<����g�+ �amǰ=kZ�jسgw�n��$��/�E�^�mAi_���L�D`ΏV��׫=�/��[BԨ�
zu;)�-��I�uT�[��ԍТ�.cu�˴H���$���24�!T��j��� �Yш�(�[�����t�C�.�G�g�D#˫Rȶ��ngE�ST�`�z��CD:�8��"FF�+i�A
l���--%w�?�M,�~ܥ��/��d���/b����]u����<�RL������!��3 
	�MLg�[�l=f?f|WQ�5�-A�xH�P|�%Y��â�nӻ�}�ˍlm���uI%��3=\�65��j�Ǐӓqj��J��J�[��(a�q/��l<^�