��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\���V�fnvx��ÍG_;�ȅe�~�>���9�>��Y;�0Ga�%m郵�W�N_k�)�����N|���ԛD5�9h����rv�\��pk�M�_�|qƉ�EӔ�6�wDiEmcd��2m��5��dE��/Ӳ>L���s;O�_��<R'2Õu������cڜ��h�R�lo��[�T�gjy"�*�:�J���j�k=�?��!-��N�Dev'�LHu�v���!y��_�$�TV)�j���t��4���x)�<%Нd�b�/�|�Ɯ�Λ�'�eV��xyK�pb���+w_��
n%#��ް�ʵ���#P�T���EMG`�˪�Hc��<�r�>%���aiK[{5R�W���Y=>�E�� �+$�V:��Q��� ��D�{�~�S��L��*,��{!�x�ǼB��ʃ�h`�OU#E��π`�q�Q��2���Uc�uY1F��Bw��XLL��'�TF��,8Uo׈��E���Dg��`}�s+L/���i&��Ҋ��A�!v�vN��!���Îv_���J�f����/��\��Yb�ԝ_/�T@��0��Q2		�H��!�Ĉg{Y2�-"�����������za��=�Qg�/��A�#q��M��Z5{�*�W�-g�C=���ĵ<wu0�H.�9�
q~";�@eU�t?����WqRI.|	�~�[��q�ke��OY������\����6���wR.�WA���&(�m�Ȝ%��q� �ߡ�U�IFc���fD�&Ԣ��@�:#~E(TG$��D�vy)�P�����vA�gOj,����(���!�z���Hm@k�y16[�of;�{T%\QN�*)o��Y��g����9�f���-'J�/��|p6�{���X$�P��#�Ybx�9�⫳�W�c�i�A�h��k��J��"�����3�W�Q�����Ap�|�R:�z�Đ��~T]�K��a�ҝ��D�.��M��WDN�2���U���.vS �H� O�X�E�n��2�7����	��"�'�RU�ܴ�bM��˼�xCk�S@ti���s�d:c���Ɨ����b'"6�ѷ1���F�����O�����GV�j_��'�ʿ��e��z���Ի	�'�(i%�2���\ǀ�;��h�\����� 4�N.�!�b�VuU����.5G��}�Cn>��ȭ�i��9ɑ?4�)3���9��b����Ȏ���_��9;\:�/�C��D���}ys<6�H ��+	��m,����~�4c���������y�M����уN3~��G��|�F�:�G�[ѷ��gK�%NJ)��V���Hn�3la��	��2���5�.%������z��!�ʮΜuxl�.>��`�z�Yn�Z�1P��6�T�ы	��.�A8��`�5�S�ŕ�'s3�{� �Ԟ��RE��]!����?���vkcr��j��ʎ=���˨$�9"�u�&���j�2�~Q�P��n;s 7�`��ǚ�<�rBˎZ�Q~*�.���֧��4�I;uFO��*?	��*��;.߉jKs<G�O�A�<�L���.�U[P	�Q�V6�cН^�EDF�DܻS���J-r3B(��?���/��
�J&0��B������Ήy�y2�+�5�?SGZf���[�d!���,]�+�R�>�r1}��z0I���^�G����.-_�'�`��[L�4?^��p
i0+�w[����a���'���U��Q�q+Х���~S\�!�k%�L��{Q)kӼ�7�iV����ahvQ�N]I��4-f����;�쫾�3��N���]�wPDV����`�� =����)~��n;"d<�_��-I0�{��G[�i����`-�16����2��#�W��;.���9\����_��X7���1o�^S�䈟CR�֚(�@��l�g4��@�E�n�i��~J�p'�#r:�`
�L�#}��l$�-q��a��+}d��Ab3��)����Itt.̦Vb���T�K��޿q�88C�.r~j�1A�"n҈��@�0�`�5�ݪu���5��o��v��rϦ�Aݬpvі�=GXZ&�q�e!F��&���ȝ��[n���� ��N���~2�������)����bI�8-���,(1�x�m�kn�6P5as��T���6���oz�#�1;ZC"B$��b0K��B�mL�
��sy��_G�_M읂/��ܴl�p`e\�k\�� G��;L�²����� ���|M��f\� B�7M�j`ɧ`3���}�*������^�ץ1��FE8W'�'�� U3>���jo-��;�w����7{�'��
�`��ک�Plb�p�F�GY#�.1th�O�����я�?)d0'�h)p����_C�����e$V�A��tD�e��r�V��o���÷{]��{2�B2�ػق�(����Le6O�k����:����!I̅Ni)n��T�ݕvHX�?fźS�W��'��sn1����v��5��%rAvOyv*�`���~ʤ/���$�y�O3��������fgE![��+�F�aVtڛ#Ĭ�R=tU�|�>S��g����n
���~+Qv���F<�F�(�m�:9��7(X7VųmnZ�\�/�&�؁��u�ЎO;��"�,�1G7��U.�w����]E�r݌�]�Twq�gBv$�"��D6���y�����x��AqW�y�_�C��^q�\��q���t�q��C_�e��!�G#C)�עXB�W�,r���	�VҾn�D����H������r]z�rV]��z�]!?|��A�g/�5�_x6�M̹/m�gP��{���DJ�j�M�Gk�n�(�%��g;4#c�1��h�<��m Y.$ �i�:�>��~,���SfM��r�hVc��R�XJ��
om@�� v.½꠯�x�m��C�RxEf���O��fN"��g���=`k�6vrW����a<�;7��[ot�р�̻�:�h#�:d9mEw~�F���k����e��QJ�j�Y:
���EI�&N��D隼�
T¤u�sp��.�E��yN}U>�A��<W3�l��i6�1����(R>�!�`�<��}ԝ��m��ئmy���w蠵��Ge����h|P�I7ʹ����϶��l�dO?m��~x��hK.*q퉶�;�<P���PL�l�߂8��n�d�H��q.*�4P˘?���"F����������b�=�ơAK�&��1�^���9.z��h�q���ܣw3p�Esȋ^
_����.E�&.wv����+���UP��Gr�;�g2�G����J+������S��#��[`��YZ�,!&���iT�^�o�4�iq�vX������I3�Fp=*1���E�zM�|�9�����f܈��]�m ���d׭/}��#�A���d��6J��
&d�~Q  1�.���aHh�ޱ9,�v���.�&�� ��C�Y7Gq�����b��I��A=�$+��7��Z��H�=��<���G;�K��,M�e���L�CTϨ(�N�]4� A^���-�Hr*G��%as�?���]a4�4������$����0��6��F�;`���\���S�F�C��[�)*�^��Qqy�Ws;�bx��n\g�� �H�����5x]Kh���C*��ԼL=-9ƻg* h�{:��3��$ss}��j>�P=���-��K_M�G�A��WfԳ�`]�k�s>꘯ښ��#{2�6�6�TC�Y&bA��md[�َQM�h��ȿ���N���Ih���L}y�� ������ׇ"��Oʝ" `�H�wcY�Ry%/���M�W��Zu�@U�\��Zt����4�%�çK���
+�Iq�oV�}����~�g��F���*^h{����L��jj�4뙀!����8�K�T� o"nz�����O�-����ų{��X	Oas��C�G�s��jG�|�r:N���

���gQ�u�l0���fXϯTw�m���k��(p�4�<wwϻu6e�g�)��H��)%{_/I@Aj�,87��>�����;N37�I��*��e<���]���^I�'5��r���@`���Z6O&Cy��j�}l�Qb�[����)%�����_Vqt2�a�O��/��r�Hp����L�\���LƏK��� W%��ԥ,~���+�?u�fL�]VOfY��C���U"����	HO�&#��wp�����UY��A�arCT�h��:��
�����F��N+��Ӵ�!��`[� z���)}#ADɹ�3_鰱[�������������i������TqP��R�D��,�����I����<ؤ�߭�)�m�+-F�f��]�2ΰ��|��>]��k)�l����:ys�>}z�,@���ۃM
ĵ7���*���ς����-�����vefT�nO��_�9"`���{'�]k?�a�mx��iگ��1�<{!�o߸���`.���|�*5=�s�(�"?C0���wG�pW/6^�I8M�N{}ݯ-�oa�k7����!^���qB�K��m=3�����~���тb!IcM��)�r��H-C!��T�ϱX'E�k���w0�l\�� "%�dS���$�@$fO�D��������|m�"Y��ԗ����|����<���������'�A����P��Q��1XC��
�^��Y���ԡ�
�4\��<Y�^�����{|U��
6��b��ǭ��*=�:��"��lak(�X��%6���lꓞw�G���� G�%lMc�������|(����/���W�l�#���Tۡ��l���Ł�`Ɋ���/]n��c$wR�	� @��E��<�����3dci@�R'թ+n��K�M]g˫��^?N	!q�Pa�	;ç'B��F�C>�l񭕻����qĘ[���v��ob�0�uL��3�
�,�Nw��G�t�Yc&��$��Q�W��3�_�l�u�Tf�0MVe k�;b�`����WByt�����"��P�B�t_~� �ߐ���m�j>"},0z��;�]�����-uR������̭����|4��o�����~�>�}�&�Q������z��"���:/��I�Ƌ�c�B2G�h�`:p�e�=0:.~���ˤ�q4R��X:�Ʌ��c������sP��[�Kn��5|�Q��4侢&+��[إA;���ɽ9��E�Qw����Z�qѐ/^�}%�%�|���T<�D��@�-ٓ� �g�X�mi~s�].i��P�8P?�k ��Q��w@�?�աL���v[%[u�~M;�S�%�ޯ������P�US�E�78fQ3�5�?w2QN�ş� �@{�c�#1�?���(�#�h���3�S7�ϯ�;�)�rRFB���y�%�Qi�R٘�j��m�9O����aP�~�������aL�q�SҜ'��{����rƚ�~"���ҢB��U�Y��}+u�1��L�d�6�j^��6]���� qH\E>�h��Ki�sP��pMR�FL$� r�DU���wh���.�m�S��l�Zirˌ:yo]�~�kB&�O��kQ(?z�/`�L��"�q�dC��'*qm�o9	�ek��1��kZz`�.[����C ��̍��au&<Zj�{�M9��^����ͥW�*�ᢞ���0��"�:vX@��g�@������}���]��٠� ���<8eGkB&.���S���) 2Ih���K�q��0H��G�����R4n'f�pG�I���{�j�b��<�OLc��	cb��6 ��2����f	�O���P�_r�lM�(lR�G�FW�z(����3Y��Y���*��i��(@෎���bۣȦ�\I��\��z?p+<��o��gk���Ҁ:qZ8ݕ��]��EЧ�,#X4ɪm݈L#�R�-��雏�ڷ��m��*wW4g��<���t��90��DYi��٪����zC�e���vg
�8_w��C#���ڗ���h��m1�8��|�.����Z8�bR	`$��{Hb�3� ��ZxP�ܰ*�(T�M�:���tU�w����ϝ��� ����&Mj���m&�\�Fc������̏�ji����liQ\<�l@(��6�>�d��DPo��S�mC�D�
���z|<,��A/:$|�8>�5�QFJM�4�\�\�<6%�x	�R��\�a�����!=��۽��4��u?h�%�
�o��KHک�F`ՠ���f��x��YE��J��)�"w�)��0c6��'0/�JP����ƨ�����ո�HN�݁KJ��ju�rJ�\�!�G<����d���'O]�g6��K]��T��&X��ns�3!ˡ�f��,�c�͚��.�1S�:��ߝ��E�E�u��6��q���dx�a�A%���iք�`o9�k�rԨ�Yl/�<Ӻ�k
:Ƅ�I��V�7���^Џ~���&�(�:��2 ��ט*�r�h�YJ��$���v5U �y\�������(� _Ij絾�%�����O�r��!�]J������	o`�:�T���@-�of�s%�CE��ޚ����%M�e��� ��~�0^ZR����t���;�U�θČ6���D�����$��t�����Ny�ͨ��w����Q��<�ТX�o"�
,�:$`
D+>��"�Չ�����yu$��~U�����.�~������=�0Y��1� %\}�����c������.'�ˆ��k��C�f�7��婊Ѽ��`C�0�ׇ�Xp`��1xӰ����2-��-��cN�l|S���A6) U�JZ��Z��w����y���@�lf]ChM^&����5��`��?��ozBB�G-�?Dh��� n�J��P)�s���B���Ԯ �!
n��� �A�p�h����6\�����M�eN/�ʉv�'�*�v�eT��Y��Z�����^u:��?f����ֵ�^PK�[�I4*�7_G���[Yz�����I����a"!���9I����En>�������x�X���@�(RF=�^'�VL��Q�6��V� ��W��8�.3W��?M��at�h�wq�=u��P�T��#[)yx�|q�i��텮�o`�s�rKk&�y帏���O?W�	t~��a�	�9�j�&��`��SL�����_����.c�*|�Y+��^+�~?�y����
.u��o�-�;ܒ���K>Ո�W��$ 9�M����(�.|Ӎ������$����ȳ�Ex�8BFM,�%_�^��}l�RI>��\����+��I��^�-e�SvC ��#����P�� ���W>`�ߡ�a����Jz�yv|4)m�s��-'�}\j���9�e��ܼFY�
@�X�p[�"j�M������}S�z͢�֜P5|هg(�a���lH�A�J*��c˼�Rw�J�<+����+�)8�fME�
K���CN���T{d�36ZlثJG�'�eknՇ!���X_��;�IIо�];5�Pa-�{5195��k"����	ή2?�G��Or'jB/]x~`���_�����;|JX~QW/��f#���f&�w�5�^�R��@�z���Ef����bv���Kz�m����zC{P\�aFL\��@�=[+�u����e�]�\n��<����Y;GK���7tak��/5K�F��� ���c�������3�B�訋VE���� �[�L�������ԫ�$���ƾ�ü��4�H*%�HyZ/��+�V��T26r�ىS��:�����d!�a�i�,�۲wp<)GˊF$���k��&J�/�`�E/��R\��#*��Ԥw遇�c8�^�EÕ�Q��IW.���?�jY ?��)��\\�+ �r�wb4����W.ɘj8���=ըi�����G�6�m$>
�ޛ~�L�B��+�7N}�3��� .w�6�����]��!�����n��8h|��i�ac�,D�{�!%��r�.�>��C��e'>��tT2���	��f�,����j�'���5(���г�U�O����I��}E�����I���/os�T�R�- �p�.n	����<����@��dp���ѻ���[���Do�/۟��k�HdQ��q�3o��+������ňY�a�p���+Ǖ08�����o9��3,��:\NV�ܪ�+U��IP[nʾ�}$�+�!�v �����$pFQ�8`��>K��0��Y,��_��<�6��N� ����=�j=���P���!O��e�
6�e8����Nk��i�.^�ZmG��TcuE��rv����_��]��Qj�bt���B����co97�ng�^ږ^D-�C~����GU1�>��mV:x��dA�i��ᔺ���1�=j�t�,V��Ȏ�n�?N;�}�e��_��}<�>���'Ӿ�V?Z�������A���� XKmO�p~���wAr�M��|�����s�6��t��ۉ�5:̩2�I���{�b��g٥�mݩA����U��sr ��.�m�>�QfxT��|OpAY=�U��m����hO������J�?r���SY�
�߅S�S�Ų�^Cޕ�/op��fǢ��"�Р���g3�bV�;����o>Ŕ
��}����縤9=�Y�W�J����-�=�7XiM?/�� YF�,�Q<����\����ZCO�
��j"���/�W���s�� �Pm�F�D���T���	\��)6J!g�y�:� �Z;�*���8H�A�{ؠ�d?-|}��f����./{���e��cSR���#�-zKN�y��B|���$靜�?�Cl�֣�b��+� U�
,����]Tp)�;k�^�;�z�u�1����� %q4��̀4[G>�X�0ݱ��,CI� ��kr��ѯ�"�P����|�����:<`"T�P*Y��G�G~��i��:�i(���<�e�n�������R��$A�!8H5��r��oDߩ-�J���uy�����5ß���N���c	����W���^;�i�-�H�+�+�0!�]���oj]t��4��č��q+�,��"K��(6��Y_�sEq�	��oy�䋳�
y�������*ev�����|D���	��W�ѻk��:91?��>2a��JL]M(�"�8���=��<@�G��ZDqӾVPk;M������FU$����M�0�f�x̄��|	4�t���$�>=$Yn|�7|"��=!U���Y�7���+r\5R$�f+��P�р�NUw�0M;�8Qaz�]~D�L�tyo�"�'RxL B�R� ��e�T��)5�$���se9�+�N#l<=���,eH�s[uN�m��E���Ԑ��6$�����>�_�)��В=��2	g� �?�.�T���^3��J�O���G-��|L��w[s��l[PF�1pt��2fv1Z}����P�T�J�x6���1���߇.k/�W��/��1Ō��h:�
�f*R'��>Յރ��%�^�)��G�Z~����"6g"9\"( ���0;G�6KaJ����eF��o�K�Hq�r�_�:g1�I�r�gv>-,�`9R�n�� ����s�L��${z��n� ��V�X��KWݺrl˯N�H�B�f�j֤�M��c����^�����1�/d����s9���I�&	�!YY%�1��ofFzc�E�
Ѩ�{/�� ��8���KF�9A���8��퀘���=2[o�w&�<��9��ߡg#@����|�SI�O���,��1��;n�ڹ(��Vȏ�����ut;;>�\3�N��>�{��.��ZX��+ v"�k!��������p���.��*Yԙ��uI�y^����B�t�Mt�L��D8�ƴа�z��EM̲���1��\����<er� 5j�R\�?��gd@���g��qDK���w��\�$6|�w��{-�ӛ�QӴ�ZiĭV��2۝Ul�a7 #�������{M5
7�B��M�(c!U���t��t[C�D"]�vw|�\�{��<��r��{ R�Ξbs����Z��K�� �+�x���D'}l���<
���O�Jn���,�$vJ���%^G�iJ�@X�|)Q���e�	$��O?ܠN��:7 Dg;��>Bq1�����m�6JwdΙpSs!z�\[����6XK{�X'�Sd<;�b�'�� �
�䞇����¢�B8�}�n'�q�I��5�4h�|Z+iw��V(^4�H$���`=g����"�8�ӞP+o�D=M����<3�N���vB���Q'�&�9�����
@�/+�8�n��KK$n�0�s�1R��cn%]a�}Q���V2�Ҏ�<7�^`!C�=��e��v��IhG6vd��-��n8�t%{��P�fD��HZ�Wn����nw[�?iv��;����xr��M"�HXk(��'�f���N�����>�n�&8��ʒb$fu�ѫ+�^g�{�l���b�b���V��1Ԍ�{�u�2�+N�Il��X��8[�-��  B46�"_l�h�7t����5 ��+Xr��O�א��jҡ��*�2�i��H�<�����
H�%X�(>���g�x��SEDP�L�Djn�^��e:�L�!@7��Bn�M�
E�Rc����I�nv:m�9攜ϑ�����ܮ�$:\E�/,�>ȫ8�o*m�jP0��7Bz��Y�A��~A���O���*�;��W�_7ܨq��@o�;\lR�&�[�TfQb�V
��wx��	U/���M=MV���H�r���M��
Q'��<�A2����R�x
�q��j�E��ϐ>��zf�sD���'�+�kM�d\aO��,��5&��(�>=�q��ߛ>H�����d2/��9*@Q�gq����,�]��g�?w:��E������mQ��	t`�&��U��3�s�H`*1�|�������쭇��Au�$�h��JDe�?�#<+��w�խ:4��n�I^��B�<p�<Z�����yh]���
~��x��|?�f�#�@��q�j�ڍ��;1�����m������x��i�������ßJoax ��)2MKk������0'ׁ��y>�쌞!�z��8��p��R, ���"�郮�p��m� �{�������jd�7�6s���^+k�$�=�.�`���]�`����-'�eb�.�]�U����W,��7�ᰰ��B};�/�	��3�9DԲP�&�=�������%GV�c��K3:t�F�tL,��V�o_�F�;��4��}��T,	�n����S���)�(٭V���[��	�K�,\=	C���J���pv��b��7<7��v~�=����5��t���O��_d(���߯��g*���F1��
��n��+,�����s�%�?�9��8vS	����1�*��ҹie_�\i~.`��ɮ��E�Md���������ܱ��(�b��7���^�M<����J��ug�j�x���+T�<GH�I��7�!�D4���{�"����먆�~R*�R��S�t�LTm2/n��yk��Db�p@���CCJK���ChT��F,Rۈ��揢'��[��	��`��ܓ�]�bPj�?~e�s�8T��g��/x�5~��B���#�tR#�H��Dp��Z�/��D$Q~\�Ndz�����)c�j���Ep'����ƌ	's/�#I[���H!�H�[��t
s��BrSG�})���yh��i�";%��5���ZQ�b�ܝnw�1��,'!.��HH�J�(��qqMI|�8a����ht�-r��$�4۠`Q\j���b�F �1A�d!�ҥ�6�{���_姞���OA>W%�����\��]�ʭ�ep�*L<\4$�<����0�"?��T��]�8+U�p�~����Ͼ���\�ޭ�X]B�	J�}e2��	��~/���)ೠ D�ꆤ0�k�I�{�M�����YMW�{�I�NR}��Xɦ %|�?�pWX�/ ��m5Й�S\EY���XYd|�x���8�z�O�c4�����J�
�<҅�,�u�g3H���gه�U%}c����o�i���
ݟ�LTJ9�<8�5�H�K�(B`�P|+U��r"������JtfİG/�n�.0-	h�L��Gŵ���od���3�|3��4�*D&qo�9B�2���l@j�mK�
W����"p���ц����,e0P��'Pk0��S�^���*���x��g����@��F ����tz��N$�U������pzf�J�ӶT��w^saa�@��;f�X)*�î�NhOT��H�Et��κ$�U\{љUg�������C���"ر��D�c�GF�=P�ž=V��wM;r�؏O�$H�P:RL��ye5�ݠ*�� a���m9��S1q��pvwߠ}��}�L�@f	�|X�Ly{U$h�	Қ���+��"Hff� T�������ە�̷���Z�K�1-�`~�c!�������m����s��Κ��Ց�%��^��d��N0)�r��!PS`�f�O��
�.��0ޔPWz���^Ͱk<�B�>��%�'�p�T�7"�U	N��X���0�w��+D&dO�,�M��Ό�h���?�m���;�4*"�H[�r�<0�㴠a/J�̆�N;~�X��7���ԃ��3��-��'���B�,��_(����p���V����\���I�J5��v����v��׹�$����Rʌ�&<cO�� ���=Y�/�Y$��1_(L�&���lx�����0��ݰ#K_�s��`w�c���&1r�[ %��4҇-f��T,h�U!�Ӱ8j��	��I]��40�5��=��~���~��5�4�Ø��_f����D7�i˗u_��1��w��"f�I�Qsr��C�4�
�*6��.��]�4˗�:�A�	��X���;�B��%4����Kh�p$1��a5�T5�ǖY���;G=�f~�LqY��
:�무����'�~�^��N��JI�ml%m�Q
�*��BhLA�Ҕ]����=m�b�xS�h��u���u��)| h������ve������H�)��.������$މT�m�X�X��Ҿá8:���.�q�.��O�T��]lo�����6�/��*�:�hz��z�{����
HՔ�<�܊�=
�&��V��{�ButA�:2s�φ22r����:�[�q?	������!A~E]�|Q��U�}�>����?+�y0�$+xA��Z��
��Z'�fv�Y)�X.p�.j��h�bo9T[6���U��}��g�,e���f���θ�53d��6,A[x�H;s7m�d8ת�d��{�q�-P��3��x��΂�AJ�m����F���ݰrd M j�D�H�p9PFqC�w*V�����zׇQ���cg��;�Fgf����-Y���8�ݕ�:��ѩ��1'� ��wN4?:�p����}gؾ�V��I��0�*�,�}�� $�=��٢~o�M1�ɴ�vҜ:�_�n5���w:\�!{k?\�s:D�}�%렡/��.x^Q����܌!��p���M}�P�B�A!��+�<A6���E�`6�(ߨ��5k�o�@�t��j�h�?�\j�0
z8Q�x�d�7�KG�-�;�����P����p."��;��ʤ�74h�w[�����k�>�v�N��<��t���z4Q�mc��3]N�zq��>%�#~;��,S�O]
�x�ߟ�N(y��v·t��������f�6��ĵ�-O�[e�J��1�#�ݴ�mc�88���h�����.)���F�'��
���]����
�#���[.u��e՞x�	�8���ѳ�Ƿ�+[���;^y�*�6w{rZ�l8%�;�~�p^�24"Ry���������:p3B��|J�*gvU����E�[��Ŏ��oj������X�P�&�� ;�k��%:�/ֺ��ӂ'l@\��&{��d+�h�焊j ��*��k��RE�[6yA;*!B �^��QHS�M�WP X�Fܙd���Z&!�����yB��w������{f9�kk����槥�(�����]0��W4�sh������{ [óр��Ei9�@�V�U�� Ղ!���Ô���ƪZl�n�U+]�Ǧ�v47�z��V(vO��:|o���}1X����.`􆃯U�q��v�5±)��D`�Ż����<3�����o�D�}誢V����O̬|ZHmOk�唉�Ic�8-/o`�y���M����J2y$O�5��&��锜ŢS�u��4Y�]�t9^66�6�)�k;��0�Y�F�ȸ�A�8�8�lzgǬ��Y�[�����C��O#VJ�,$x��A~�᪰t��S��~��G:�jK��ɒ�����%��,)῔ɾ���o-�<U�k{+K�$W���[닢�|������!�͂YU�]�EN �T��l��+����%T�ghc��VV���T"�_�,}IvP���� �f���Í6�U��ۄ�~����I�!�p;��l���2����!�p(k#�$�EK6.���ia�vhhc�v�!�:�j
j8GI7Vx����ك������U�hA%9�i��)�BBjKX�w.nf>��o�+��<�n�`ĜA�|�B��-Om'ƕ����H�ۼ�/\���'�	5��N�M~��îW Ԑ\i4������ϥ�`1�{�)��e�4S-��e�t����7�|�����9,ɼ�7��&v{�0D����4�gK�v�b��뒳��3Y�\�cV���rR��[D��e����P(m`��n�f����٤�Vw��wCq�=�y�iU��Z�}����K���@���*�%\�{��x�3~�9}!��`�?\���/A�x �VhcQ+��[`4j�|?v���iݻu��p29-��·��$�5��c!�9F�W���A�:����Ɓ��6�|j"ۨ��=�ޣ�]�=���˝1�AJ5)'M�(��s'���iZ._o>c�K�vh�{��r�x�'w����|7����ya! N��gx�i<�����?[)z�yw�mY���K�N7���@��#�8�E���m~� Á+G\�T�$��y�T���wN��K^�/�E*9ȹ����
�8t񛤂%��D-�r?GwTP���]6�/~���\�D����9��D�7��c`��`C�I]�2J�~���\`�&�h�鯩�1�U��|���W����B���V�J�]�,	J���#� x?�+��i4��D�b�3OW���TE�&A��@NG"���尙y_��6���:���i�D�m`�پ�G�t{@�/��ýWߓ�<"ku ���-���hu�4-��a+c�-�)��`��~fβ*e�,�w���y^�*Qy�Vw�>TB+��w`ap����\U�읐��r�=�B�w��-�D�?N:;OK�������
�jٔÞ�����z9��0�� Jd+pu�D O�)e���6]b�$�0ԙK���b���V���i�pԬ��k�@�B�v�2�sp��6���kXw�	��n~����`"x-�Ӛ0�&���~����!���(7e�H�Pb��i2��ml� ŐOQ�Zi�7�fa����n5Is�8�,F��tb���fD�e�=&�ln@����
�����~c� ��vR�?�7.�̖E_T�$K�p|��c��e�����Ϸ�H!.�N���6~�(��&(�bʕ:b�iO�~�Sw|I�������~�7�Ie�g�f�L�*g:Z�Ɗ�����Z�-�0��2�l��r�l��xk�X=�����-��#��D?��ߺz�-}�j��9�}-�J4���l�>{'�������:C�R�3��[&�1�{���3�=H�i#���i��<�{��~2�����+`k����I^��2H��a J����,�I݌�J�B#WW��z���/��a��I`Pa^@�)�M�sl78�n)إ9�T�[��Q5i��z�U�c�>b?2~|̘��'�q� =���6łŢ��f����A����XW4
���V�Ч���ֿ7�3�Uf��e�F3����*+jEӉ�B���f��W'���-#��׋|40f��y��O�:�&�!��Jh�	�2$Q�`{a�P����U�	A�q�wX&ڏ�J��y>�ǎ�'Y��AH#ʊ�x߮�:�JX�m6�?�n�,���\�+Bl����^W�3��'<�V�}0�������Y/O�Pn�"�7�F(��j1��-ƎyU#�"A�Ȟ���{����J���xȹs�6�al�����)`F��à[h}+����ڪ�3�Ks��,9PB���Fg��k��'��b�K+$}��
�Uk&	4�	TCݡ~F&�p���w��R6��.��:�J�@vAM��65���4VaZSF�������
�Do���9�%@��4+���RL�ƙ B�F f b��sװ�Y@?f"�Z�N��[s�uj�\!3w��s�F}Rbz��^�<��#�G���+~aq)���G1>���w�U��a�"&x
��!�"A��ό!��$�(0�/��3/᭣�'I%�%r��g�x�D���\<�p������WJY�3Mޕ��\����Or���U�P��i���y�����|��}Y�hTX���g��F���7�Z��*~���Q����������>�:��W�o���Y2�a�h��UZ�������]��v�?	ӿ��A��jEnb���ۀ��MP�����ʃ�����ӑ�LoNθ��|h3�@�:�& �r%z	�5�����#kf��3�yE905[$����5Y���)ցt�f����������Ԋa���Br��]�'�����.UG��4��<OӶE̓���'�`���iۗ�|�T,9s�?� 6"���e_���}�=mܔ��^�jj=�.�xP;,��v4�&�q��)�Cx���I��)�_K�����+}]/�/��G�'��
~r���8�e�>�j���xW��d�F �
?n��[ߒ�ro�W)ED0⺭S�.�-9j�HqM��Ӣ�|�z����5��֗�kϸ6B��|	�D��ү�����N9'�8�|گ���g�ay����7
�"w�B�E���[x�n��iM�r��-��WL�\~>��B���`�]cRn���r�F�{W[�?~�hi7ٺ�)O���X�W=�I��q���M̮���3�?A��^'�� �@v$!Ʃ$�ͤ�즘��)���ҍ�zh�PHwp���~�����-��:k�Ou���!��V�Ɗ=��/l  ��t�Z̽i`DЍ��r+�R*�?@��ea��1��O7�;F�dgSV�@�d���9�L���/�!����g��%C��N�^��<�e���дd'���+��;�|���쉷�1��m"���M/�r�NT�F
���5;����4�r�m�l,pV:pIO��mňÃסY����){�����~��t�m��P�z��A���*զOv��<km�&���lS�hu�o����q�I������<q�6�}��d1%�~�MA��q*���O0J~Xf�<��	ԼBJ
�h�iSQ<��mhugC�����o_&H5q
`��]�(j�9���W?�wZ3�ݵ��ꠌM1_=Έ`��,V���Y��xrs��f�5N���"�D�}�x�������X�� j-�+�?�S��c.=��]J�͗����i��K���(
J��|�"q��mϚgD+���=�M��d�5
 $�p�8@��E�K�=��N�#??!�o�eP��w,�(��/׬�~��VUٝ��{���;�En� o��bx����k3*���&ވ=��J#!='d�Ey|o~E�aN��M�4.r<��7]3W�[Lu��x�w	�yV@:g5�U���Pu&�O5F���Y��x�_���Z�����˧Y?�.�B�%&F��
�/5�|����"����ㅍ�N"��3�V�B�N��0�<Q)�#����G# ��e���f�Jy�!zFM�	ށ�/] �U����S�;�56�����	1,2���t�4eH#��|�`Y�f	�nQ�L,۔�e�%G�B��������ˑ�֌	�����Sb�!@���zy��8��sV��	Ʌ�����J��,���7� "ecJ�CG׳�XL���'6��|r���Du�Uv�A���Pu"�.�&�'�smA�2���s��M�
�U�#O�J_����;> �/t`Cz���2ù%v*�ǳ5�u��/<D��`���w�0�|{�?�HBi`����џ=��#��1�+��$�=sG-�`⿘@)nn�ǲ���4�$�k`���d���n0�K΋��/Ol�~�!��|1Hg-=���E�צ��UO:7`�I���s��C#f�!D�2�O�z%�`�}t�*��s%���3�u����_C��(�W�?�>g�w� MC���,�l1P\�l���E��Z�j֣P��J�{���H��)`C��eø�]Z�����(�^d_ N;�����4�G�fm����\Q�䲹�sqtf_��t!�4ķSd��S\�e@�^ʶ#O*h�(-�|��=VX	�g�wl�����AE��ފR9���L�7�L�ׯ�6�S��*�-�ņ�;����(�jw|[�5�X�M��5���~��SF�i�O5YwtW%D�E��_���k}�<K}a#8 �s-����hjňu��:'�	@�j[`=�D��9�������OI���t��L�"�����Wx	��sJw��9ף�L�r���yp�N�Y�.W���T����}���>�(-�\�_�t��j���d��zJb<\v~^�<�߶�!�7��b���'�=A�0�����&�&Y��7l�:ŇPQ՟f�*PiԚ�G�%@/���4(I"Nuzv
���1�Ѧ�\4�!aZ�W��7��p��ͻy��L��CM����f��#��e���L�Щo������ń1�Xx���+K�����D�ˎ�Z{U0�T���C��u?)��.�4�Z!�Ɇx��i�}R�Q�ݹs^C���Q�La�z�n����~�F���~���~���ϩ�62��V�X���׫����#,c+���j@�؎�)��I�hK��y낸*Gk��,��䈦a*��/���2��HA�ĉ���%4���z�u����7�]@��9��(/���\����6A�������������'W�Sai J�v�h���|�����Z' ag�aZJ��Q�hX��B5v��tz�D��;�� =U�=�6�[�y]q�������Rd�~�F�KA]-\��yMy��6���^
�F^7��������
�Yߥ�z^�)�&��(��D�d�pW��%�8�/ȟ8g��j"T�n�T�x�&�˴ 
t��^�rKI���S�'RIn�pڏYb���f�6%p�G�8�w���u/oZ��o�IRXz��8�>Rprٳ�����tU�٘8��`U�Ֆ�C��Ĳ�?����/E�$���_��=�	t�/Bt� ӭ��.,��2�� > �2�c�ØF� �9-�G8ծ���w���QA>ө�:��X{-�D���ٱ��S�<�sA�!u�H��-�)�b{!f�~�{oI�R/�[�����y���o�g"��</�̴�9���7yv)��X��!y�Fz?�i�֨��!���d�`��<.�A�����EP�SB���t�����[�?���@l�ְ�RaZh����9&�ס؛�������'φf�/�x��|^�p�rU1����7�>��E���3�K�_��U�����&�J�����E��������E�s�=sѡE�꿑�~��2�/�o��FB��i���N��oq��E�u���)B� Зv������X�b�㻋�����^pX��RVޮ��a�s��f��7��"'�ѳ:skv��1�����!wD(w�1Cд��㼺b\X����\�|�����o�ȋ�s	{ �"�6�-�)u���C4��c��S����g�o�@(����f��g�%e��Gn}j���L5�8��Y�ۍf�k6Y��#_��o�WV��ZX5�F�w��Kp�U3l��>��g!m^���7_�MoΕ���1QC�� ���u���b�'RB=ҹk�T�j�}Rţ��a��!�_.���`%�ɰV���b�����Y�~;��T?�w0SHvr8%��<����߼e�J���@ �6��P�EU�&��0��K�����$5�ct�
�r�_�[5���ļPJ)s�*�Ǿ҇� {��j��#�i�{��)h�7`J���+v2��2#��K�N)�8�6E�� ��7q�<�P��,4VT������:B	XI���z���3�3�\V���YҘj�n(_E�^��7Q���i\�qx�Dw,w�M���ˎ&K�G�����������H��`����k�Q�~�Z��GR�0^DwQ̯^���
�����fIۭ����[!^G���ΖG�B7�|
(H*�E�a��H�^�O�eK(̮6�Z�%F��;Tߨp��۽^��Dz/E��)�����������V��\���Tl�ظP!��3݌�����+^+�=���[�c!x� ٌ58ð^�=*w'u܈j���"A�vz�;�i���]G�2�_�dQ֜ۋ��:W�n�l�MI�n
,�f�Ǔ��7�@���+q�i�:��j>�>��)�v�_��;M���
��������]Ώ��r��;0��	*v��6�1��XD^��M����vn�^�����3��>b���|�}+��KZ8�ZN���N�!��B�,����1�8Z��
P�I*x^��>��ї����ҧ���|b��s��(���4�DӃ�P���8]Q2 Q+a"��d���C���E��-� �W�P�p5\9be]ª��$�� a��*���~���H��5v�ȥrN:��՘��uY`����M��-:pt'�B��F"���w���#=P��ތ�_`�����o�y��)~O������N\�*M��>޾�d�>�}i��h:��U�M��_*ڐ��Uv7��}�~0&8b�`Ik����=ҳ��k����U���#M����'�.HU��j �]��ë{<��^�o\��J�����`-�Τ��&(<�v?�� �5Ձ���f�_�C�۔��B+�ff���V���u{�(�X���H�m��eo�Ԅ52Q?�����PnK�6�H"]��#���y�p�y��Q�x�����~�h����˳7��7 �^f�^J"J�0Q�t���H��������6�)�Я�����H��M�jPfK%�i{���7��2�`HL�t�o�<������b�\v=I!WFj	!8�n�1���\�%��Q(f�� �i{�2j����@uJڰo5�-߷fR	sw���%Q!*F�Z��4�&Ǽ;!b���}vJv\�a�E$�R5�����*8�"״�A\�Ǵk*Sh�M{c�C!�� U5Z�e��eA���9מ��Q��c��,ya~�/˥=���~�cuQ�=������e����.���L��e�V�~� ���r��:�b�������������?�?F��\_���Wz	��).*ύ��vx��I�
��R�r�d�+�."�nޒqi${�c��ݡ���]�����LMCk ,��'� ��yA���o%(m��%HC�I�W��ɯ��2���ۑ� (鴒�re��?q�K�OP���6>�Ot�v��X����>m\Yе��Å���� ɉ�`��@�+��-� �Ձ��Q��c��XnD��Q�K�!�%��ˮ<�hʓÛ��D4z�ؙ,�h�ن��S$�����3�I��5��H~e3KƢڶ�`ءMt�{ٖ���Da�ED5od}GX?,�n@{]��
J	l����5��մ8D!t��Ȟ��w>�B:6!)7'��D�B���SK�Z�:���+��kaꃉ���C#�l����@-s�o�|<񙰨	6�jT����w*��}X�%=hM��S��� p��k!ȴz���qP�:�sr:A�$�r�̣n������G˲�;26,��E�j0c�bo
,u>�����H3I��A��)6y�Y�ao<Љ����]��z�� P)�V*83Q-jY�!�����Ҝ��ͅo�K����Q��X-ǆ<@,6P��J�|jM�=Y�Ȱv,@��Y�����S�VU��`{��%��7i\)�0��g�Ep7
���BΠ�5�4{�8,~��y�Qz�!�l��qGt8�5�^*����W� ~�T蝊�/��Ȟ����)V8��48�d��#Z��M1v� -Y���~�,� #����߶��]��iy=;��ױ�C��:�J�)}=!WoQ�7,��	[�l�ͨR��V��q3>�y�sC�,�c�2�1'����AVP��g���Jk��6����%~<
ɭQ^�];�8�$u��M�L�g�}�Vu�O7��U�{�����r����&����8�����V��
O��gL�@���Bg�6�+Jd �ʥ*���?��ipl}M�ffD�����m������@Է/�!��,�٥0 j�����e�����@m�L4��0�^ ���m�DJ��P#��]R4=Tݑx��S�2�Y�/�&��e�l���%{�	��nN���ߦ1\��|$�c3��"�7g=GB��k��������a���Su������Ɯ�3»�+��}��$��E@�1e+��wz����(g��.�4l�e�$7��.%,29��ř�pE�6'
Z� r�4�*x�q�� �!(w#h�$�A���a ������F@q��+�Mxa���V�e�	c�	�Y�qO������n�c�e��0i0(hs�~�ڗD�[�!���[%�Z���eY�Ņ��^9�Q�aګD��WwrF�v�8�R���^���iS0�?Բyi���g?����W'���u�vB8��g�!R�H��`g*���d�yņ����Rq���,��!�m����Hf���2���<�����;����� �;��eV�y)/8	�"����w �	1�Hx���ؗ�ƨ���t�=�8�`-��vo�ģ�m6�(����*[�G/�r�Pz�����T�>�¡��hMt���;k��Q��3����P'��>��D[��CU�uW�|�<*�Ge�BaG��9�,&��K1�=A�(�E1hpf
��k^C�� ���I���H32�b?Ր�<��b�=���z�ӄR����٠��Hnϭ����:	���1L\��X���)r���a]�wR���[�lc@BJ��~����X�Rb��NgP�9�a4�Bu���;�v�pm�N)i��>'1A�i�v���S�ǽ���귭4��Q���m�NQ�ax(��-���y����4�/�+�!���K�ӌ!'
�����yk�[��꿎�� �v�8X=�P�q.��p��}��N�K�@�]�Gs�FE?ҹFt�`K�2�u�{(����F@џr`���Vs(�M��}D�8-pS4\gm;�&&���}�M������f�MO�S�;k������V����p�|؟���;|���;U���!����=�*d)�%�'��j�l��f$����\� A6�$(������O)X�Y)�e�æRYj����e'3�\��8�d�	���3�Di�a>�=y�2{��b '׾�1����bb���
�2���=+�!��-d�����k���1.\I�?Fja��k�3�u7l7/�@�1]��I5;	�}/�h'"� �!4	�k��\�O�U�ds_�qsճ+���4=(`r��'ڛ���by߳P���S��`�RN�\S�� 9ѷzB=Ů�8���������Ʊ@<M��Zw���Z��NCj߆me�+ϷAxZ+�����4.oTʅɪ�%W���-��vv���<��x`Z8s.�)����pG�H��~��iAXmBI3f����z?>�#�MPSF��T��OXw�Z?)-��RQf!�o9���X=��(z�����|X1�5�t~�/�@��|2Lħ��*�3�����76$L-�γF�����_`�NPc:FLi+��cϙMO>q���rM��Ɓ��&�4�+�8��1�wO�6�	�VvQY/�X���7��4��f�$|����g����&��y��5��=lY�J�HFGP�{EV9F�HUY[OH����pr����;!PzjMS�������K���}�kR��)�w6m���������IV`����@�T�� a`j0�"Ĝ��E۵�B�ѩ�J��PX�?�f�r.m�*��rI&�տ�\xK���EJ�Ei�����wj�+�k_��C�����ă�@��?���6b����p��{:��oHۉ�9T���C�e��$5`f��d�®:VkB$1���
����`D]�elj������,�P�+�Nq}��l��Aϔ@��cʬ_�(70��A�mR٠wP��4X