��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|e����M`p���}wi����l׻�ti-�ou!��mڊ](�����G)`�o@s�lt��M�x���@�8f�Ki-ku�����:ru��p�Gs�n���:�y�3�(sQC��J/�.,�v�0.*3l[�Rs��U�y�_�G���Q� v�^"���"�Z���Lpۋ���!b��I�rV���)"���	t*�d+0q.�zǾ&�ƹD��	��4ŖS��j[�&�XguJ
���4���#<=H�f��
�L�%����DM4Y��s�/�m�\Ʃ[n�~�;|T���;����l�P
�Lށ5,��D!R�
�g��ݿ�ň�n~C��wu��\x�-�$�y�ߟ�f�ĵ6��`�s���Y���w[+t�8�L��ک0�����0T������<�^���J��̊�����rF����MQ|� � ��>�[����@�Z}���D�	��Q�[�vޛ����C���|��������ga��}L2��ס���n0YR:Ε�:k����9��Ht ���Y���
j������B��X�r��^C�K"��A�v#m���v״Bի�aJ��i�+�p����r����NpM�]���&HF��ڵK� 2�#����x���"�!xo@4�kAb��y���&o}���R1�$K����e�>Q�}���8�c��=�,�����P�6��g'�V��K�6˖�K����$��,��K���v���?%�&�<͖M�ῤ�/��e���Ap���D����g��RNՐ�Wݛ���5Dw�2(�%"Q�u`��Nv�
[^O�����%�NJ�iGX��bm�+%���F��m��A����x��ϡ�GQ�T�5�'��:s�az��9�~})wQ��H@D8��uU+}��\���W��ʞ;������
�x8�%��}�Q�䢠�DW�㍍��T�&�9�XT|�K^�'o�y\���6��'�A^�麋��x{t�Z�}�3&�W��#�o ��(b���V�5�iF�; ���ɷ	�[ݣ44.��M���:KoiWG9)�.E����C��׎2νM}}��>
�?�|���Ta�7�)k0hc��T�K�)/���D�]֘����r����n�D�s2s
���-Kb��S�ˆ1U�r8��6�v@N�H����"<�]��a��`F�Eq[Ix�6�( ��'���}`����%�qh�Ô䈼;y�@���׌_
�T��Q*��jT7�E���HZI�5�H!���@��S�u�Lቫ��T���A�����az({�8%`��?�/��N|�u�h�������{?v,�ƿ��<�O�$9Ƹ�TDK�p�i��N��B�I̪Җ�j&�YÑ�<o�t�
95����
��9�����=̖ &d�)��~�G�$��P��a8��aM��}6W�T �,q����H��H��7�Y�R�{����ƙ���Q��TQuDE�BsG���U&��C�/�ԑ�$	i��&1�k������#���G���{�Y�/�#�ڀ�O�Cm�u���^5s��PJxM����8����o ���'��@5p��T�\���q��nF�ʫ
w���tހ�%y��o�mæ����]���8�q�r�2"rVx21�N�b���P[��KfG*�aI<ޟ��A3%�������t�����_��%��F�W}���%��QG�x�(�H:��m���KG���a���9�K�8Jtpx��8���G8ƻ*��F���ܳ'��m
�XeV:�-0�s�љ��w��l�o}0� ��&��n�_G.{�O���T]�L���/�5�;�Rć8eej���@��*6	�sG#����L�i#�(ų�^�l;�L�
CH˅�A��٬�f�cP��;�0B7���O�3 �˯�����)#LXU5�f�aI^��0E�Q~�"�}��⋻���.���p�NϾ�;�d�����>_$<:��� ��Ew�Qg~% �_�5��}$��i�9@���pV;�?
yE�E~i�Jp���ed؅�|W��<?�b͒C�cPz)���l� �M�5����� /h#d�26�!�Ƨ�r�N��ڵ�L��𦁣���y��v�ظ����\�ku^�;����s�6$؅o����!����"�gb�u��U�y��*#�B��$WF�{��{m��gh6f�܈6!��O)_4��9�&;g�5&��f��2�۪�U�kJ���YAawpK��Lc0f��IF��'���>coY2"����
Ǒp@�U�nğ��֑�`�mժ;r.ϸ`���e�3'P�*���c�����[A������L���0�E�l�c%�ɚw6��$���1�ߙ"ni��ʕG9��	\�Z5a[�Ot�(�����N��U|���5�`%fV�U��<	��g�!̶�Ǫ���7!���
A=�u*�v������b�4A9�蚉m0t��_�CA#����XB��e���'T�#*E?%���i�v̅����̦��F�G��/A�=n|L,������l�$>�<(�- ��>��x��"nU� ���[�@�Yv���M� ���Y�ۡ�P�I����t��0%��'�3�sV�Eź5�&幬�	�v �j�������Шk�$`���?{�a�������ѳ8��_o����RKP��׶�,T�H�]N���̄_[o��F�V��i��a�����p�S�z���h��rs��+ \u�4�Ȭ����5$V'�}9|�֫ϣ�-)C\};oGd_>�K!}4�pe�J�d�}�o���9�)B~�]ޫ~�K��KD�@'šf��Jk�0�0�f��b�<��"Ln���=����ԣ�����aA��uy��Jz<q[�I�?��.�4Zy\;1!�X��y�blߵ\��_2�D��^��qȵʣ/���&	8'��<)�%�����{6����y�iw�$��v�
(kDn�"����"�{���Jn=O���B>a����&��8����>LƇ�ZB¢����y���m�h��ΑHT���.#�~z��`(z��;2��5�	����%���nb���YL>A��h*6�q���B�+�{R���}uD�����Z%,�/�����+:Z�49���>�>�a		G�6�����2!f���=�R�Mu�*���~������NE8`�Մݻ�:���1���`>�ĳGXm�!�y�e����*OP�}�*�_�oq��n���
2�?碽`��K�;6(qGA*�	�]��\r�>�q�;�z�*ԛg=!�Κ��_P���~m�)6��8��n���F�^o����E�l�e�q��X&��%�Q�-Kr_G�/�ޯ'@Z�J%�E~���)I�_k�[3K��Y�oXx��p��gIO�21h�Ư%Vs����Yr�6����-X�f�u�O8Z�C�΂M�]W{��M��	�%Z���ZW�i{��ʜV!��&U�ۻ�C��z���+���y9�⌫��2�j��Rg����r{v ݅�obu��&�S5:�eK�8���I�f�^��@����K�Mx�K���l9�֘?Y�j5���}����)U�4&)EB�0�����{�XUT�W:-��s�"[AN��	h���)<��w��T������@���E�����~��s=�k�T�G���̖4T�j@����n��A��<}%��m�Z��8}��$U	h�p��5[N���р���P�}��pAsL��N7M�P�K��?��%�<L;����'?�+�D0gSA
�[���(&y���4X"�>�+�C���a���J�b3�,�K%�8���r�FZ��A��"$7T����S�����|T{?-���N	��"&G�o:��f_t�#��9,5ޢq�5/�Tf��]���~�, x��ؚ�P<�Ή���h�������a6jD������Λj�q��6�h߃Saf�ݏ=�/r�.n�!d��@��6�|)�րO���rt�"���-�(ʧ��(�x�
�� ӯ�E�Bv\�G���^e�MNj��3���_p���9��xK��>�ύ0��rۉ�N�x�(=���nYd�̛�3*-�Ϸ�H9&��g�a:H�\��Y���?�-9���Ƨw)4>��2���)�-��\P���c��YOtȯK�E�X	��U��'zLG+ӊ�<���V} .y�Apu}���l�{�B����j�dzoIMU�'����E-�bɚ7��9��k��F�c���-b�����`�i��Dz���I�ҹY��d1(��h\���K��<DBi�]/�L�V�ȶ�1h)FG�At͊�(�[�ͻ�C9040|~"qۋ��^�?'��9���|
)�깺�����H(-Q�n�px^Χ���;�y�w$��{7eK��od\Gnz���No��Uo�h{v79���<3����ωbⴭ�:�����Ն~��c)��C��e_E|��O�[O� �ݙ�VK%�W��`͍r6*Q*d�����{@��J��w����� 
�.�P@0�@X_P����G#c�T_����؍\�!�pd��
�M�$�N�/�w
��5k#Q�8�T��m���?%A���<ٿ-b#�T�x*����C1~��)���O����[H�k�"��޸!�Ұ��N�����:xϳ���/�#j�7Z�+'Xw��H��W�pYC��;�@�k���G�W/�_��9��F�T��h���`� 	sY�P��ټZ��k�7�ll	W/�7�0ApоE�Z�#��]#T�`��RL .�YޗN�6��%�|��0Gdr��<F������Y.nI�@s�E֊VZ\�J�Օ¦�<�����Q([L�[�F�� ��=�Fg�(r<����<
��� =�;��)n4�$�$tZ��Uā]���sYo�(Z�cp�GsL���`آߏq�?����	��ūƜ{�j��C �PN+c"�����B������P
��Xݐo}o�KnwX4�#��f̶�+��PN����a�D�99��X|�o�U�sJ��-��[�{��F&��C�۱c��]�I�W^��t��#�*}k2��ܓ��:���-OT���7n����U�
������R����g|��iԴ���Y�)�'[�zs%��3��p��'�q���g%�K�XL����/���
�[���K}W��/��k"n�R�O��F���t�n��\1�����=L�4��H�-�Z�ݩ��.]�����pD��ֳ��x$�g��}��&{�K���!M�{t����ǀ��T�(�h�+�>�7�E��3RB� p
��nu?����G$X��M�
w^Ŧ�bN����5��%���Q����Ƴc���ɜ{':�Oh$���%K!�2�ɜ�oR�paА���<^	��}4�����yf1���!v��N��H/�������J��Ab����|%ܲ���1�w�+�1�R�I���Iw�og�]�6�F���ԉe;�^tcZ�o�W�.��z&�F:"2h����pG�5�|�'ܢ�N����_Y~p9����$�&'��pQ���-�E��侌�\G2����ή��|�6� �ߦ��||Mj�ջ�F���W�z��%\.N��@��h.��Ġ��>Vx�k����dRUw�]�a�!��8��`��!O��q��}�G`e�,̏-�BѤ�[�GxޚeFW�J9��Pԣ4|�kr�"����y~��EH�t@L`��H5 �1O�$P��_��ٗ�Lb%l��̈́�ᠨk`8W��a#��Ɣ��/T8�qV�⯎��� �w�����!i5����s�-l<'�B�8s4{��ܫ�ov<	� <���B�b(������uaت�����p.9�ۃ��Y:W=�i��Rއ���%2��I��pXGT�P�0y��}�u�򏢌I�@|庵�ֿ#��cc�l�"�7:����N�jь�C߁Y��칏��S���}�UR�^/� ��l:,j��K:�x��9v)+h�I� t������0���xP����=�� �l"^�2��-k91����X����K�	[|*"�W�{�z����-��X�W�n���L>�nk��(���P�ԁ=��!��/򹫍��)&����D8ʊ�M��Q`�V��7)� �t���i҆)&�Y^�����&\쫙Gn"�c�XTd�m'7\�zt��z�r[=Bs#�ho�}�i[��M�y;�y΂3Vq�q�(�^�b�i�;}�H��M�=��_ �A;S�u����c��yr@i$��7�����Es*����jpD�p���r����m��H��(��^��{|0���S�4���`Y��c�v� �]��aMN>����8��f#^U:4�n��Q�}����������&�F	7�T;F����h�Ed8R$?��! �iq)�OJq�����9��ڕ����H]�U��GzGģw���i_q�ȋ[��Y#A�Ǳ�N��ߴ9:wi�����f�'1�*@��p�O������i�f������b�}����՗���JR�R���U!�� �б��XR8����mձ[�q�Z<�M��+ie���ŉ��!Oʑ����l.��7@	,o/�Q��x�	~c�X6�[OJbV���ƐP)Ȇd(�#zu�yy�t��f��ToX ��p'(6܋��W�N+�M��E�m_ۓ"�e��ƭ	I��P2t&C����?��QG�o�Z'��R#�OD	H_<'wy� �%譗���R�lP��u{,�J~V&��C�LwE<�Ҧ*�/bP���2� t��I=~;W)�I�~�c�8c��'q��Q"�(A?��.	�	;Պʬfo��]&}��>}������
�u ��&i�?�����&���E�ݾc�v�w��U�d��3l�l��~0pɶ�3Ws�5C�)^�P,*	,:�K��;&n�8#{ãW�
���*>��`�ԘͶ��qz�jq�0	)I�C����RJ���<�~uXx_��^s	�7rP_Mq�}��1���`x9���J�Ρ�O��*]R����pE��\�'����K\�h�ȿ��@���?�p�!�'$È	�5���I�Ç�j�K��G4�2~�\�k���P$i��1���C�Z �ڐ,:����iup���+^�#��h�t����F���U	�����q3��>��� E=��A'l��@��$1�*a���j���6��9ȭ����a��5 �� �T���"�y�U�ƣ9Q�c���ׄ�c�ϳ:GeMC��"����I`��Dg�̑9��OB�i&��ҟ��A;l�8(#��Qe�C�w�~�tg����Hh��R�=�ENjZ!�k��qU�����_7��a�^�ևi���YE�}�$n���N�俤�A6YA�Ө��������f�2bePC8 ��鳯>^��H�4�M�#{a��<�.�`,M��hۡ�'�٭��u�L�m��e�2*,���RX#�e��F�|���x��\}_l�&��V��]�j:A�Љ�GvV@݌+��U?V��v���%��M�a�3Y ]�ӌ�FK���.H�,P*������R{'"'�
�\;?�|�O��דĞ�9I�Ͻ��������
I��ӆBE�6dW������ڮ^T�+�Ԓ=�(�g����|i���h��h�b���9��8Ie�~R��t���: ;(O��ֶm1�$�oY�|H��7�oK���u��'�i�XA�1�Xp��m5<�vK*S�7�ߵ�a�n��\-?eO��[̵`���H'�������$[����BS�`�x=��A4���������3qVX�9��ճ]8�JZ�5�	1�c3E��|SE,xS8P���u.7k*�O���Gӥ#��N���n����@�O�����`�jW8��*�A5�֕�����wW,Wk���:��h�W��=�具�l�?F�����m�������֪���Gi"�,�3P�I�S���7������w0�@�qb�bF�S��P��_��?�t�3��Y0N[��|�2�-;+쟔Q��3�k�"@��~l���� ����T�"fDv�KZ������<\�f�u�#��ql2���ťrx�&�[��1�<9K�랛(K�{(�	�V�#yɽ�J��4��N��8?Ǆ`Ny�2$*0Q�rV�Ѽ�+�:�M��a/�;5)P�ėG�Z��Ч�q� �'X���T�p���v@Vps�����Rrބ�D�����,{��o%�|��k�2A�P�:��+|��Y]6��8n�vV�oWf;�Z�>�.Lphs)���N�L��d���!�"�pYj����n������cl��� Nڛ���͌f &#	'��}\�X��Ӷ��f�p=E��E3rkCt�^ߺm���Db�7�[�t��������#pX4,HbK�L+�&켎Iz(�M<�Ф�]iǅ���w�m�q_P�?�k�Z�BH[�}��ٽ��P�E���0�!I�ޜ��T�O�	�F�n���@\����<g0'l�����B�S֣��C|�a�Ή�B��^����I|jv�r��`�|(��+���y�_/t��%6 �g? �$.���s�����W-��61����'4O����e�<5Cî�/��5f{c��$Ͱ�����F1D��*"����l�)���,V�6�u"�~cWA�]�j��4T<R�%	�<�4N��rE�>�͸ !w�ሳ�k���(e�\��V�6�Q�Pd�܌�*̌�<r,:�]_x1qbf�'��?$% ��]5��F���(r������4�~�����vx�ι>��}դ�u����ƕ)���Adԏ�u�H/N�50i���]�Ŷ���	&?��5��&�3E�]��nЀ��Б;�AX���Oe���0
Cݱ{�7)~�"͍U�;��������#{ܑ�K
��a�fs�a[	/u�N��}�W���>�$�HU���X�/��3b�=
��ї��� ����4tvz�!���m��2�ɤ�N������J�{&��R��x۠|%ⱾF�r�(���[SV�y&�	��q��Et��L|��_�M�t��I���u�r��Zd�[$��+���a�A+���
�����=|� ��
F`�+_��m607��>j!���@e����	1Wmz��D�&݁\~�E��"ɉ��(�,�������b�ek��EI����P����2���E��������Z�!� H��;���ۿi$}�ev���i�j�9c1gl����Z4:&��q�s��4h+'i�?�t`�>�%[c X-{���'����k�˶�fS�z7��������_�<�k���H=��J�x0�+h#|?-�yW�O�3���+u�q7�>yȊ�a�^�;8ӕQ���0�r�, G���>�$|�[���\oO������r��i?��%[ �y�����;�wγX��-�]�5�^��unG�Ǎ�/
��E����v�HGbXF�4�`�S�����y:���N��to�p��ZU/v*���@\��D�?ʀ��F(߇:���E��5��i����Q���ַ'���g�*�-a��e�Y�cw�^|}�8  ��,���5����Z=��l� �A�Bi���G�o����B0�ah�'C�D/��>��m�fw���[��W2a�(/��Ll��/������;�.V�i�wd��_���'��t��%Ú�>n�'m���&G��+�lϝa����&lm�(�/TN�`�����p��d!�Җ�����Y��S���������((Fp�멿��ۉJ	&�{A�f.��J�X�iZ��E���:��w��S7�
���oҦ 7@r�UI8\n�'���\&#�Y���q�S��~�>����:�y{#ye(�-����s�?�כ�����+�������+7q�B�Sb�3����p�<i-7���c�S�J�=�d��=�})MD���R��7�݉=�|MCqH�' m�Ik���t	mD� :��T�X�?)�iG_ �l�R!�%�0��{�*���;��yr�%��M��!Z"G�u�/̒U�.@�2mU�v\���5�+;��zx�L
��D6�if�9����KtYH��2���
�f�v!ީ���?��J���K�Õ-ϼ�up��Y��Ϝ��<ţ,����K����d) ��$E�]���p�.ū�j�"�Ő���=�!���l��1p���l��8���Y6"�lwV�%\�
�����]�X8�O�㙑����t�{� ��-@$��0W�G�6q�dr4�p�WT]���E �L|�$���r�#s����&���3{l�3/e�T��T|~#T��X�F�u�������2}>ޢb�	!�� cD��J����� 1��]�/�.&���N�e_-u4�st�0�q �N�m�e;�[X_`������Ш'+H�yUQ�g�zF%����Ug�qR�xX���]O��j�9���Kxv�v�N��ō�@ڛ�	���u�8�X�P�Cm�_� EI�Qm�xxoX,��Z�� @a3F���"dNd6���^��/Ϯ��o�����c�F�UhUj"%�{l��u���N�rx�#��� �,oA|dz�;Y���5��dED���r����;4�MEYs���*��gi
_,G���L�h�O�W�5��!Π���ӹ��I.�Q��#��lq��pk�x��gb
.`a�ﴙ��hg�cG�ô�"�����?"W���+��挝/��P�!v�؄�[[����AV���V�z��[�:�x񗥐��0�9� N`I�@�0x�4KZ)�����0E�>2�<㗹087Z�NgHkc�'�њz6Om��ң���!0���t�+�Q;�J��������}�
<#�UGx�N�$�Q%���;C�;K�z�DY6���
d�����+��G�����&e`����W�����	p�q1��&�[�ٟ�U�RS(��jF&.4�^�������Ԡ�	Ϙs�������-}+4n�Lִ�*�rp�z�����k�ҩ��Y!�hpB��@�!�UA.�0�8�0<lb���Ť����Ut2���룵�_�7 ��A`�<���RUD�Ǒl�O��y��d0"C�T�H�/;S�)�sJ3p����ͥД؛��D|C+-L�~��E>�`��/ŝ50�E����tNL�/��M�-`/m�2eqAy5��d�
�4oH���[����# �Nl�}�.���5 rP��AF�[�}�T��2�gw\�<�6�!Z�����_�4��r@���X��k	��4��%t^Wt���˾z�7[��[G�����ut?��V	e�肃w�X�O��S�IVb�_�4�f�&���>�K�r�����Z�8n�K�6�܂� f�:h�$
�zp��,B N#Q�pR	�3(� ;ӗ�?gw�3���OV�s��	 �n�--�܈Q����rD0�m���Ԡ�8]z�� ��ђz$W�o`����$��|GN#�K10�Bn͑]���y-����H�ƭe/a�ay���j��XK(��+M[W^ٱ_|4���z%f�����`�6��@f'O���.E�z6�SkX�J�2�V���������V�?�>-��+�3���|a�g�3�E"�a�Q��v���7ᚋ �F=��U�`	U٤�6G���N�.��ۅ�XC�8S��`��&N@̫���r} ��z�k4��3aMw�IFb�d�`c��C7�ۢK]}�ҾpS��{���(�/����Vئ8y�Ѭ�\:�W�(k)i����U����9��G��À�
zb�dw^��W�|�����-���`�L5�t�W��W�����i o̹=.q�͂��&�Yp��9I<�a��G�V��*�A�\�RfUI����1�7���[^~~��X[T�l�[� �6?�3]B�T��ڄ�/�=5�J������!\�pU���1��~��_G�ƻ�M���m��?�4��p�ѻ�yŀH��o/vr�u�/�wT՛+���]��锺�S싙�/�u�*���V�B+�q��Y��J�V�*'�w�W����ò���k,���6�a[cr��i�����H,�hO @�i�P�K<�}��ls�ގ1��gb�W�%�'�]8EC�-�@9#��ƞ7�mo|G����� ᐴ'g��q��Ƞs���I���3�!��#� ����P�>�#"@'Y�� �<��I&�zf�-�`h*�<H�S�1�J��Z�N�2�� 4�`SpP�Ͽ� Q�^��-/���g!�E#�ZdN�n7�)^%�4��^:q���@�k�EI�s�Ъ��C�(%;�W�C�Z����Z./��A�:��+��X&�2�`�AI`;����3ꬣŷ�B���R��=�H6�qy�D:���D�D�F�&Z����9��������n��LmAb��%"���P]��[���Z�}�ǒ�J�M���x��P"�<�#�AÙ�p�d�V�0�>xu��V���Ƈ���M���y��6�	<Fᘍ̈��p�	(�y���v�*YG�c��wT�F� '�e�+����.dfx�~V��F�4�\�zU��]�1����y�xJd�T�o�j=m�&�$�s�:���7q�,�`��M�j��v��M�n���4I.��`�X�]��D��.'����a��ΣR�`�\�_��m Z$'�ْt�79�oq�(^@N�"U%YX�x�¶Qs����sL���Fm}��vb~Տ���d ���� |�=�Ũ�f2<a�+�G���s�r�q�Jt��\���UO���iP���Y��k1C7�hݻ�K��,��?b�cn[����O-4�.�����0�X��g���6��WS3�\SMY����~D^�Q6�X�J���Т�U0Jv��[�6���CYl�n���S�Jԏ��ɱ+� SdnA�7��� ��3���EC�0k8����>�����=+�>%ڥQ�15��)]��*�]�+ڠs:�Q���'����H��FcϲǮ;@a��d��˕1&b�Xܵ���}5�X��2.v�d���@n��7�n 3>F룄�<\̦��h>����HUtب8��Pi�#~]��;ñ�Y�ޛU0BM�� ��f ���PzJ1% ����6�O�
8��{�y�E"�'�:��1BEͭ|��k�f�M+���L�=e`C���|�l3� �q�D�4FC!w�FΪ�voY�˨���ķ�}6S�(D}E�H�����<b��N���w�����Fi]�͵��挚�ؕC��K�o�ٜ��<9�h`�B�������xG\87X1E�H�'��|!�NH��_�����\�s*>~X}U�{Ƴ7�跅����ߙ>�)�F%1X��/�\���_�D��aO�pRJC����2��Sɇ['{�N ���1w>z�n��g��\�d�?Sa��^
쮄�q�T��a�/=��_���E��aʊ��s��E4�%�,��'�p=�2�Ӏ�wa�o��g@��+�L?��x��%iZg�8ou�K��+-��@��>I�{~�u����,��Sۺ4Y��.��im	��ޫ�.E]��E�~ܠ)EG��7��H��l��(���7% �;�%�k��&I&G�gO�g�6	��>�jR�A���F�
�-��>9:�3��2ag���u4Io[-U�$��sw̯�A5�Q~�x�ƃ�s	�����$[]����A+�݃�t!w-B���x��K�Eǀ	(	�Y0�R*։7�[0w�(y5�
ş �r '����rfԢ�C��a�ڜ�b|9��pq��CF@�b{ J0Gԍ��:ȍ��2��9UqA"��,Pz=��K���;��I�4������z�(�)���o?P}y��=[�s���2��%�����Q���%��۽0۽�hO<_$�"��K�d���a!�]:M�)7���nX!�C�mz��F���S�7�[c�a���g�؃QU�ք{�(ŕ�sv��e�K��mY��H�΀����X�bO����iL]�,<Um�l��q�M R�m��ó�Z�P^�]D��>`D��*��_����,D`�{Re��֕`�W�f�4m�\|%p�^v��SJ���� M����P�GV�;A��dy֠�]�!�ϱZ֒��D_&	h��," Ç��w�������]v�7 
� ��͗�ѫ�k��Fg:���D,�i(ZIܳ�

�o�������KbP[
1C"Ut��M�
��?l�>���tE��,�ٛ+0P}������܈;ذ��d��ɧ]i��%�W�+��a)9Q���S9�|6�=b����Ϯ�H�J���\���kB�k�����'|�}�<{��ǩ�>=Se>�޾;�8͖ة�9�����b[�c�Ī٦֪�IP����ΜҮ{��H�9����u�P��:�F8�ι���'c�`�YG6b�]7lq��/�c�5m��t�����JʕhÉ�'��̗1�:�Y`�}�6䐿�YЪpD#<��;9;��te3�%^���P�T���1W�XaVc{0ry�#D�rJ����1��8������Ɣk���8�w:������(S��s$d6�r��Ɔ�|�{�^j�]�'R��W1)z�n��Z��Jg��,��m�n�	U���K�>�ߖ��r�A,t���Ns�:�>{(Ji�DN_4B�����p��>��HIЌ�5��nJ�����p�uʤ*H�KtD,���+qf3QW�s�����xa�Z�ZB5:�l��2�/<+����/�_NU�/��L��1*��,�[�$V�܎�%O��,�d���`�����O=ق���IaU��9i]�� ������$��?�w��vY?יk��~:R�����O�v�|��gs EiGt5�(\L��=��*�Mo�P�e�������aט�cե�Ŝ=��i|��E^�B��cɭZ8����?h�Ѵ̪`P�w��*�\Lr4��E�((9!����mǺ���O~ש�퇼����'�\����2a�/N���k�� 3�kPV+��S�i��M��σ�ahZ��1]5L�����)��% ��(r�VP����������o�W'Y���(�����L߹�N��B{���j5���-s�E-U��#��T�F�q��T0-y�O��8��Б���IÏ�8r�m�0>�������4�H|#�Y�R�0�?��
R�]�2:��x�"rL�t"��`�������H?e���jf��R	4i��>oX���ζ�	,\<�4ԑ&<���q�����m�6N(� �o�������Y@8�y��IF�h�Bq�Ly�XI���+�[bq��W��Y,E�n�ņxHoF+M!�_���!�����»\���O�Fe���8eo)��eѴ���� ���f�����}O�S�B���Ӽ,m�2k:�7���C���2�6���ӹ��T�5��S�]�	��r+�sQ�-Ғ&#4��*�h#r�%޳��	md����o; K��m���W�������R[R�Df�6����q'�T�˿9��?��Y7)������d�?��\΁Aܗ�P���u��׫ZC�,x��Zp\�c� �-Dl%EH]fP��BY���x���qr�8O�A_�Ĉ�H+������r	��/�@��u@O�'�)��m���I�7�c�1w���x����"Ǔ_�1�Eb7���j&���[K�t�����M�3{��Vmog&���aV2Z�M7������R ��c��!~� ��lC�H5������e8.�M�mG�/~r��6{�F�#�K}�/�nn?�~�x��Fjpca�=�>�⌴��($�vF[u~(�yvFx��blI��E� �nIv죆�����9;����R���ؼ�?I�;$PITH	�v��}����#�^����,3P�U
݌u��	��\��u�������ksԣu��l��D ���w��YKK�AW��x�tK7P2`;��3��~��LL8W�N�2%W�<�-9�k��&�%+;��n	��i�nQu����ΧC�
����ط �2�?���1�"�u���y<��E@!ُz��W\6���#/-� ��'2��<ls�-o0�K\�����SI������Sd����Vq�����43\�2�8�[޳d�?��i�����h��M�D�����'��xil9�����z$�M������Buevژ�@�0�����{P[3/;�+m1�e��t�9z"�M��O
�GN�k�ֱ"�����$���|r��ߐ�������d|�ekX\䳩�PQA�(w�~��� "{���F<�Y��x{}�{�a��f�?�=⊹H��|J��@<G�Xu�'��х��� ��o��w�/�A���o(��b��1�BZJG�v^'��a�M�k�S��	.�u�w���=��2͚���x`k-B�i6��2|Y@{1����7��{�1�Q�	C�t�&�D���t� �'��%ɿ��R�����(�$���ЌEcGYpE�Vb��,ç�"0ΰ �JV��/���gyB�ƕ����
{���N��mf�e����v�uE�e�w�>X�\�?^F��	��޷L�m��S�ყ&�)<�� ���K=N|Ǭ"5�+����3	����2;��R�?��&-�"�r��!���R)c�?s��H�l"��v��\�M�Z���'0U���yR0��ۧ��U�/�v^+}��M̥�nQ��
iw���(4)�WT���i��^ȥZ�������R�K9���`�%�#�Ͱa�$T�r��d�∥4Ru�I�D[�������x���W�[�{�
�e�Y�7�ҟ�{�lh��4�i�p*Ms\g8u
؁U|J��lB�Z�XI��Nq�N_qxQ�n	\h�0n՗��5�&�T�oK����Rjx)"i��M�c�9�nb(!�}�j��,�<���Kl�r��cu���XsV��Al�-�IdpR��|�w���E����	�����7�#R͎�L�O?�V�V�i�~�B54��S�0ت9�;~��k��n�m6��*(����,["mb�!�Z}��h�[%CaT��#�}=���0P�b�|kV�ގ��氓�(�JԾ(*-�k݁ �N�Z�*T�:�4v���U���t4���>!nH�U���ʝ�����`Cfh��}�?��4G}�.IԹk������ӓU��+y�X�ˌ��WS���<��6.�4�-F����kgtxe��5O�����1í����r0v#.&"�	��,�O�2b�_��B�lkQH�t�Ϊ��0�O��ru�Ǩ����ߡ8
�߉���`���GR2�G\��E8�9L_bM�Џ��o��a̥���'�щ�Jf�B�b{�5HQ@m�#W�<���DE汒bo�������=��`��1��7?���*d^���h���!q�85����u�dh� Lc�^J�ec�#gw֜���N�c��l�\�'�
8'�;��NT��l� j�u�&���WQv��tjJ	3Bf'�@<�ܼ�e�	�:�V��1�*�:�=�:��J�y~���l#������ڞ/V[����튠0�Y�T�
+��%br1ԓ��ǝQ0i^{���ąB��@��gy�����4 ��].5#���A���oF=�l�0�t��=BD�%* '�=�2z����Ѷ���*�k#X�>�:i}߬��� 7z��B���)�t+�	Q����\)R雽�8�S7?
��D�O��������@ONܻ��'b���������5�<2��>?H"P\Cu�FY�<Nl�>��v,K���m� M��S�#��L�Z��9r{W�q'�v�m`46g$���b�5s[���'wv��bm)��ICz��̌�0��8˴­,UP��n���{'���`I[��zX|"����E:�3ˢz�����Fx�s�y�+Z@"��G�4ޥ��=>��ʸ���g�\�%�:�-܃oj�\���t�Gj~/s�u��N�W�h����T�+M���z�=�7��/�P����б��k� f�P�:�Z��bۼ�-��ԟ��(��O(�/=Ua�F�a�D^}����,=��j Z�����_�}Rt.ɣ�໫�y/k�G���ꂠ���m��n�ЦB���2�^��ށF�Ը��{�T4�T�Mt�蓉J$ �o`L�|�O%�u�>�r[NF�}i�_�����'�Bp%�.k�9���$]}�~�A��D�+X�����L�8kYL�ي�S�}���3�*�c��0���2�U[-�����o����H�f"��|O(��3�sQH#fF�#�J@'�BPV<캸�GS�m/#g��^Bb5��U��䱴5 Fv���z4T��n��Q`"	��F�+�ֲ1�l���?�o;L˚����S�a��;��i߉��U�W��/a�w�oL/�{�a�\��?�ݭp/��yg�� �B��xm`�%�qs2�d�^�͙�������~:�#�]�.p���T�C��?��c<N��
�PO�ʏ�K+����v²���2p^;q2w��8����ncj�<�A�&#�b�φ�d*�����a�BD�
_��­�;�|����5��&���ˁ@��LE�6`�A}E���4k��ҋ�#�
�S�*^��۸,��7�zfb��5���ޗ�B�'�k���=N`t�٘� ����������O��_"UG��8�( U=l8����$��h��j�Ǻ��eY!|�Ҥ��}�ۜc.'dj��Ε�õMs��F�?\�Q�4qL|�������s},ոx�](NY6��+�@o�DsW_z\�?H�!��ϣ�"�FÔ��_/]�ʉ����+�b��֖�>)���x�x�<)mmM�C;�@#c )��RK�<��rn�񊍤�s�/��;TA�"M�9�>_B��BP4�:R�8�5�&�j`�mLB�%`��\���eF$���ۮ3��ø�~!��@k؋�'{�g�uC�
`IG��e�#�*�J�r%�y�x�����38oT>��B%%m#���CN�<X�[���$͜5�M�m1��ך(��;�Z�o���:���T���2,xd>��Oаbo����OQh����^U�F�o�˦��k��񪨛����Rǯ��EU\t�i��%�G��Q�y��aY%0�f���5��n�]<L���x��Lg}@Y�f�Ԇ�H����*H���Y����̦f�R���zĵ���e��q�5�![ 9A��( |���B`�T�UI)8�p0D|�-���Up������oI,�h��V�g��ZlKF��A�;%d��� �75@��c��4�� V��'	��T�,'e���� W +���W�֦p�x]��XqQ�6[��,�h�� &'ߜ��A�=����nm�HR�����i��5���d �keZ�.-���8S����'�5��c��e@�]<�
�?��!�@��	k6b>�������if��r���	����7{�Ѳ�)e��BpY�6�P�BӲ���^�!}�C�	���y�%�����{D�����0�JD�R�L��\0-q�L�t�;'����뎰��~���Z3�	 ��|��av��R m�$��eI����sEO�N�5�ң�\L;r��>j���s#�vbG��ZIO���!�'��hGSU��@����-���Hߍqk�)��ν��$)��~���I�V��Wh I�!'�F��2�N���$h>�b���O���_2e�������2M��UON�d�7;�i�H��'����z����t��12Q���YX�O@v)�w>^��]��S;�9�.�\������׫c*|�۾�v� Y	T��\v�k��k$eؙ��	M�ie�^�&?����v���?�������k���9�Şg>��w!k��q3'[#�{93�(������E1�\��aG����c�j�J ��Ӛ�����`:��~�^�Wu�Ί˾F��@�r�(7�n<&������c�`7�F6cT�7��~��DvUu�Q�s&	#�,44>�S{��u��1R�� tE�g1�b�f>'�Z}h)�Q�+�V��t�i����"���
/���qg֮"���qx��t֞�2����\_�5-ͼ>KtSB^��+r�H�FM�G�T�t��t�.�CN���3
<�:�c�f ��s���TF�d���ep��J��4OhN~�jh����<�y�)=E�+�o� |v��s��>��v�)����a�v�o�'*������Mg��
�Ҷ�Ρ�A���F���r��Ch�-
�93�����)Ѣ1���fv2�sϵz����/z�|W�U���#��N#��0��I�W�Ju�c�x��i�L<A���㋷��X�W9r��T��u��c* cyb�98��l,��\z;^�;�8oh򍻐+C[��Z&l^�׿4`��:���j����9���i~���>T����}��\���m- ������@�^v�g���VH�6��;I�X�o��~߈i��V9/��'�@��{%�2�8 �,��/Qsl;�i�Y�*���+���c��$|4yK	��o(��&�a^b�ٚ1���|�_���W� C�nb����
q�Ļ�t��I�+ =��F�`k��w�" 0��m�"@��{�e�J3��!�G	r�&��Mh�ث��]�x�u�G�>��3�R嫭�0���H�AQ^����;����s��?�')��]ތ���E��,� �n�����2��Ɣ�MF$�ӿ}�o����
(G��R֊�)%{B�ұ�ɉ�rrT�Wp����z���˥ ʶI��ϐP��z"�٦�O� ��+��~��h=��p|��K��3Na�p-��)mHn����=(}2dI{��ω�Ò�]�*B��4l =�kYΜiZ��3H���\��$�P~k\02�!�.(�_�Ο��kh���8��zt���n��#��.ܹ���o���P0%�t�3��T���dYoWR0`�.5j=8�@b�z/.=io,��G�G}�����N��#F<���są�����;�w�2!zO�S%[�N�瑱�G�K�{;�m�jw�wɚuC��r��q5 �_3fkε��Ӷ5�)��O����P�Рc��*���i�_^��Tb�B H�2��|@$sr:�y,Ió�ѿ��R�t/ �g���]��<H��e�~��ۏ.�P���?������Yl�r�4�P1�'Rcn� �۝��My�d�5<�i�Z��d�� Y��d�$Um��x�|��M�Pu��
��R��^�~0aj:�Fɇ�]W2���H�?�C�&�./�OorA��R��Xŝ��}I����z%�4]k�'a�㕀;&Ԭ TW�l���%򴻽��]�R����(T�)J]���/�j��M��@�P��A�!�
��G�ӗ�!�D��0
"�=Tz{��e9��2���k�;�e�&W5v��	z):C�*��<�5���'��v�V�1iBxL�f�M�a8;#Ա�~x���5�����)ɻ;e�"�'?PK+n"K���?o'fE
�O_�h����,T��²����c�`O2��r��W\�H��t0좍=�����m��1�M"��d� h�ez&�b�>#�
%;1���������ʆ��~��5Bof}S�^%tЈ�
�}��بJ�d@�6S1���qh:mgF�`�k@��E�?�ûw���.��\s�PJ� Rp��M��[i�l���pƁ��b�!G�Y�"T�n��&�U�}��Z�J��#^�Y���@Yų�C2r�[��%��L�ix}]2�-�\�5��㡁�w�X%V��1�̞�>R��E��\e�c-ԩs�i�*��d�w�}��o�'/ �;_]:*3��)���C¿;��$��0E*r�K��@#�,��&F;l��\�("�0[@Hn�v���m2U.T�B��x���,!HO�`���C|�w\YWy��B��:$�^�h��֙�s��
��u	�.��n�]���a�{ȴ��p7n}q��Ť�%4�A����8�iEK0�a�����%�3���7&��@��F�)i��R��) ��bז������K���SO�OCW��4�V�7��J>�O7���Ҩ�
��&���|����Jo������bk�l�t��
y/�|�[��F�V/$����l}�w��B��y�,���b��&N�[��IV�i�f �G�f�,f�&R�`�(|�uX����4˽Z�����������n[+����DH���HR��tN��{yx�uH��;3��m��Z��Y�zGT�.�o������%q;��<����}����dX��m��xQ/��|85
�r_Iy�Ė�o�,	�C(ػ�0���n��Cs���%�o09�䶄������b�*��/=��������_�65���x��@+����?�+0�m]�&ϗ)��Ic"�r�!2P��O� �����!�uN�݈2��j;��ihR�}�vcncR��^��J�ح��m�C�S.��;�(c�N�-��~�zl �J��~u~�_~L	7e\���-e��� ˋG����=�ah��� ��D!�%�D���^=�)v���%��3�I9B�BVSS�O�{��^����y�;��=�⢯���D8i�����=�f���E����%H/y!��q�;>,�%�(�4��&���ɥ,�	����g��J΃Oy��8`KV)l�aD��3$���Y�/0J8�MX}�h�l,ϼJ��tMP�-v0*!���W�8.-0��)$�@��@�6W�=H��9�%�����5%�SAM�zJ1*4��
	/sd���v_�4��ۇ3�+q��J���9ϊz�1���Q���D>L�4,� |�9,��nmٯ^���IJ�Φ:Cm���K
]�ck0�*J��yY�`��V��=���g�I�䟫RW�G�����`]�����0�QG���TU�,)�H���JPE�b@�7�t������N.�c/�2|6:~4(#�	hi��\���(w��L!�1C���/Q���NEJ\Ҳ�"b���D8֨���������~��E�
4�}�Bɠ�bY��}�u�����$V-�&[�	�p�X��<h=YJ�+;���X7�?�������+
z{2#���V8Ô#�f��sz۝��6��P�ŏT�Yy�����;gd��:	�9�T\<3=:6��ߪ�� �+���]G�6��7l�*���!��f���uςk��H�s�C;k���S^fܲ쏭p�� V�%nŝ�a�SJy��8ܢP+�$�aM	���	�]�_�{�v��BD�D�!`����g�=�M�N��ã1��_���R�!�9}�&\ݿ��z5�R��.lVX�
(t?���
����4-@ḻ��ft2��|%3�����l)l�ޚ�N_�g�$���A���sљ�G�T!�e��+jS��mͧf.�֢ci�0��k"��:#@��	˒I� qRb�,���?njڤvn��C}���=Q��7z��Pݡ�-U����\P�:K����@�ؠ���o�7�@�:�c�̻�y�)��Z��=�"�Q�E��.��g1�Z"Ǻ�R�.�-��um�Fk9`֢ٕD�\����m�Z�\g�s��<�J����R�k$)��1�3�����}��G��D��2�s����]6��ř\z3'}�W�K�r\��Bb�lsVRM�1C�3,?^�_8���}t))?;�`WK� �J?�a�|��
� 6�(&�������~eɡJe���/����A4�{;�7(��QD�E��w�/�������izV�Fm~�y˗u�7�N�e�� �eg��oU	<���Q���ܿP�%�֗̂�ǘ�5��%��@Yu���c�����#�5��u��%V�(^�*��;���Ή�� ��gS��o��͢L�8����;$[���/���U`d�4
���'�]����T�3tMARU��T��@0e	��x�-��2֐'�?5�S�b���\�3[�g��tůd�?wL���DjR*C���>Ղ��m�W���ԡC�l��O�8}ޮ�i����_�V��n�\V	ݫ�M)��ƻG�rC{��׾s���D�j�UոH FM��p����8A����Ʒ��G���.�����R�K�:��7�ʄ��K^�=�1ol���9�B�]��s,i�%ݯd�A�2�g�g�F��a�Y��kt5�ޅ�3��p���@�:��)���\���p����:[�+~H��I�� �]�ӏ ��]��-�kEv׺C�`��9���?�)W�k�ʘ 2�zLڜ�.�TV\��M��p��HFnuJmO� 6��D�?�eMט�K�aá��G���q!�4�_��)ؿꦯ��|��6S v괕����m{��B�T�R��Q�Ӗ���HB?\�~� �L4���!���B�v3��0��P޷$4KO9�����~�v=\Yd��S�L�p���<.0V�1u��m�͉w�l�3c�шKt�P������~��/�Tja��L����w]�;k)A~P$����T��l�t�vْS�Y��2��?���4����zf�
�nsH���g�j7�� ��X������^]"H�$���u��x˔�7-��
�YT1�0���Mv�KǦ��Ȕ�S2p�ꡰ/(�v&����%j6u�"�B����I1[�'T6OG�F���8��R�A�������c!����.!c�_�{	hS�.+��+"�g�˛��p�7�GHm���]g�����7X�"{���!ٔ5u-��IN>H?����_~���4׀�n}��n��:"���E�L���V�!9[�
��^��F�,���s֋��U�h�(I������&K$�g�8�']̓�<j��X�p3t��l�j7�<�����\n�f(�^d7��F��.	@[}M
�+�0yER&<��T���B�R{�����m��p��~�2N^�n]�M]�b!7"��k�M;��ӣ��
���1D6��\�Tlai��C�@�%�+�W.��YV�kB5��t�b��"�ޤs�9��ޔ�M�<��zu	c p�D&�i�$X/�����N��%�r���.e}�|S�@ߝ;�H<�/xZI�A�c������	�5>ܘ�:.�L�2��1����w�,
fW�����_����/T��<��uH(zˌ2e��{ 2B��o�C��N����y�c�"��r&���󰋚o@c��!U�����&=1��w����?\"�5M�1�qZ�Md��1"SᠻNڡLF�G�HT�����n��,�����>�g�S�k_&,�j�Y�k�\��Ÿ�Nc~�`gz'@�W�+k�hk���jfv�}��gV=�[��s���}4b�
AMR�6>�FV�@���0�]-����1�s�g9������dZ���W�z����������l9,�vN}���ƅ�z���JW�N0� c���u�(�nTL��؟e)bk��"��漋��,�R 3�J����G5�s��̞��!Mq,�*�b�3��ϏWd������}���n����[1�� ��%�J��#TQ��`Kvq��73�i�ղ���蒗��|�{�� ��?���*HO	�][b�s�P6kf.|�>t4��/�Ŷ��!Փ�ԣ��:�>�W\��!����C_�r�B���u��GU�4�N�A��:��'&���M���廗C�ʐWx�� Yl�ۙ��=���iRZ�$�N�/ҫ����+!��X���um����?ͥ���O�g�YU�ѡ����!�a�w.Wm/$��`ڮw����]�[wh([�'n����8�Qx�� �:��� �5<�}��Q�Ǟ�J�~WăW�7l��x�����Dʕ1%rQ��F�������W�z�E��c��