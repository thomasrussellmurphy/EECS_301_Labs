��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\���V�fnvx��ÍG_;�ȅe�~�>���9�>��Y;�0G8є]]�d����k�B�Rc(�4wKK�,a��$�T]���R+��(9?��D���t�v��g.>`���� �����1kK�A�ô#A�vz��q1R�(ӈ$T4���c���T5����8���&�U�����8���n���N�����f=���ph����T�U�{���W	b�^*Ӻ%���;ʅ�:�D ώ��=�0���=ܝ�e6����Y.��񰼗�a!3J�����_o@�����h~Y�v9���秣�G��@�r�A�w�)KpwJ�=����[Q�����^4�W
��d�}��BX3`����#������o�c�}��|�t�p�������ףm���N.'�6<ɑ'J~��29�J�զ��k"2�:�n�W����Pc	����xHR��)�c?ɫ959��*�w��y�L(n���Lpn�H�Y����N���������KpA�p��"(�d_� 4�JxM�`��ߋA*��`����-h8b���a����i�W��iݖ���z3�8�n�{����J ���)�PPV+�яf��Os�{�!	Z�\��󙩙ʞ���wJ�1?����%�rD}uѿ25�O3�DKU���>�29�����K�P{"ݚ�;cZ,���ǖ�2�-�-7�˶P~���nhsv�o��L�x��+���"������-v7�)@��b������lp�ć�L����T�SݼI�(��(��f,���+2Q��6��6�pc��Zv�w�}�:Ԛ�� �N�p��䌩�o�
/,��h晝���˯��p��U�h�HUs��[:�����Vig]�DѢ����������о���2�����~^պn:�PZ�'�v��&��䎶����u������G�A��i�:��+�_�I���7-0`���,�42�'�m�9I�J�b(��P�s;�b���E�P��@�R�IKO@.C+	Z�"�&�>[J�Ҷ.) �ك靖��z�`��f��MP$W���L�߻ɃmR�'�螴)TO^�5'�;�G�[���m�g���j�?��i��c7�jэ6�Q�	]��;��DF�}����k$O�-�������0�:��8a�7�Nh(wa�x9�B�f�U��5�Z�y�	\>͎��Nç���]t<z�~������L��Lc@�-J�$�|�y�o��Ǣ: k�ޱ:���v�^�����#BTk�݆7�8��b�PXR���6:L0yrX�}#*<̑�ކb�D��]��K��H3z� 6����
eQ�3{
mcv�9� ld3�P�c��������i��Hv��v��M��_:y�=m�M*�jTsW�4nDƬ��X;�_��a7�B r�Ų�$kaʝ��W7�YQ+��솪!��D��]�3+mШ���S����a/uq�Q���Lf��v��t�P���,'���F��~�g@5����G��vBbpЭ�L��fd��NN����coO�z�aٞ1^h`նx�A�
�S���a���٥sĦX4�r�&�_�!W�TxIu�()o(~��}j3S߾{"�C������Uj���v/�����߰�0(v�/\n]��[�-Ⱨ����|I�5����OPõ�Z���NT�P�;����U��i�T�_T�Fg�~�ؓ�4�;�x�����x�YNmj��o����cQ�00��:d[��L���:e���%��������"���m3?V]a?�=Y*���Ԯ.��W)��<F"Mlk�5[Z���� E� �}_���$Y�q{M=le^���<	3B�9�� ��ɩ׷jڨ�by���oJ�d��W�?����Φ l��[�tD�u�TW�;��`�����������faV�b
�6UjF����z&]_��P"S�O�(n#Ƚ>\7�{��C��x�C(�����^1J���l~�2����jo|3=��E~����i�6s�?2Z�ZY�T���:�W�Eg9I[�.��9u#��*�@������k�C�be�wƔ���2��,���yوsp�0B���"����)�U.k	�sd�����~o��mDzȘ���O�A�#���Hh���.����Fi婘!�>sȧS����Z���~̜n�=�2�F��Can��Zk?�Zџ`��%�SeNʀƪ�BU�C{D<Ӄ{�3ЍUvGۈi.������؅�t�	�I�aƨ�/�f�n���h�L��ߩ��ze"��U�Z� հ�$̨�ؒz1*��S����Tjd2�����T�A�(w`���Q_���V�)>N2���@��g�0��!�ey^�C��"���?���4#4��DL�|P�i�ʖA`��m�"t�By���e
&)u��͝#��W핡hr�1����5�{�����r"�X�V�sk`�>࢒7���||�����;$[�g|e�}��X����3~7�Ԛb�5%����;�_�'+�T�L�I����)P�HOŌa�Û<tX9`��Ӓ��oP��,�'��LNpf6�Rҁ��|p�Mv�#F�2.7�e�9��9�6P�h�*U��L}%)^As޲g�3f�4:k�sf�hc"R���)���=1*�ؼ�Λ-����93�e����'�=�uF.�_F�Ǥ��rD���1��&��qg�>������i��vAl5%Jx�������a�	�'^�`��5�w[IH�,-�W��I�2����^���%<�+5Q�(3p���6RՄ��7q�����@fDV�w�r�#A L�7x�؎��<�CȬ?!�s�r�	�tc��<��Y��.����l��?����z�[���ec�,�0"o�h����zf#y1?��c�[��^��0[Z��w�A�L٠>0�ٛ_�esxw2���=��9���H�x�|-q�M����;{��l��� 5�qϺ��-Ƈ6Q;�$�C�y����U'�}�s�[Ĝ��q�?q��ˌ��{'��-Ы]z��z:]M!�dv�[{�D�]���u7+N9��KI����S��%�@@0�Po��Bx(A#]�WU�Y���KbF�m���M��0�q�"D�7yt��%�x��'���q/��f��N����r�9m�$���W��u���[i��J� |���;����\�fS�����gEA�IT�m��#ۛR:��N~c��*'� V�B	�؎��_i�V�4�({�eӽe�/͇�4H&��rf"��t��˨�m8(L��y,���ݮ}I�k�ŬF@��4���}��$n��Cr���+�e��qg�ւ��~x^e'��&g��pJvYBR&�f���^���c���jI$
q�Gp>+���2������s��bO�w���l�v ѾA(Y���ŋ!W�2��ya��}�72|7i�ꫜ|l0�&f]�M�VCBgw{l��W���i���ֆ��uٝ��������(�pU��+qM�T��m��_���B<��A�}A[B�T�#�ck��3��� �CT�R=X�i���(baȂ�v��Ċ�},=�1߲)����܊|u^u8f�YM`�D�P�В��0$��BF��c^;[�׸�p��1����:T��ib��WnM���$��?�˒�������9�����B��1I��E׾!j�ׁ<\CQ�k	
�a�(6�`�M�5nJ��%�Kj�3b�n�,~��r��t)%�`m�!p��)��ȗ=:�bh���aQ�M� M���oj-�Sܪ�+�@"�����y�IO!����β�OC��{�֭tv����2��ѿ��\W�[��f�l�����J���;J������\ܥ^,Q��mN�q�����
Z`B/~����V'i�f�J�8�UD1��L��ΰ�o�
A�C�v�ϭu�"-/��匒0�D}^-Q�k]�����8����[R�
ؕ`�w這��oB�j��?g��#�?�e@a����i���[od6����!�NK��砎
���}?r!�(���Dp'X/����.���5��!���8/���k���Ɓ~��;�q���R.o�bE�~�vh��u��H��T[��zR`f}��5��i����p�:�Ҁ�M�,MV�X��Z��b%�핯am���!��V[���ˤ�7����Zfh��;:�ʣǓS ��.S:8��2�oY�?$���2I�w��_̱��v�Z�`!�{B{�@��Y࿴Y�?E�*����ߢ�oU<c� FqYG�(O3�E�m�o2�"����;+�l�h�s;_��|�1�� ��u�*]`�{	6_`66Ep>^�Ks�b�}(�[{�/*�N�0�cڭ�:}�P%�\մD'v<(U_��&��I=��Ixd�042��A&!�I��ߵޯ�S�D�A��[)��}8���|+����c�G���R�C��D�<9˵ɽ7��ZQb�6:(�F���d���[������f���y��[6��t��2M�7y��a㒾j�|���>��:�D���
(W�+�F8�j �rtf��y.��C\����)A�jj�ڞ�.=��Y\��4�<.�j��;D\��3c|������I/�A�7����;N"-�-����U��1�i�.��K�<������0��%݉)�x�=l�%T��7�J/��}juZ?;��dȶ_%э@����8�c���z1���)���1س��-a��]�(L�➗�*c�M���E.�E�|~h �y�r����yG	�|T�D8m2O�
���������k��z�ƈ��m5QL�qd�F�K���[��bBX1�&ʉ,�\�y�Ė��R��1�;d��!b�.�����U��th6r��4�Q�@8�6	m���+�vf�&�q���݌���-q7�r�ì���Y����ix� Ի[V�U`���A��:q�~oꃏ��yoWK�� ��\���_a������>�F���"���J��'\M����2�AjM�!}`T��vu�:���A�x�q���z�,U����-��r�X�*GUZ1,���b�Ru��y=O%]�K��cj�E����Z%s��p:�k7���F�>�?ϑZ8gD�;��<f�7��b�4Y�T��ꈼ����v{�����Ă��b���b,C�0;��U����}N�9�X
9� �=�򢄪�3%��wλ�e���RG[L� �Ԫ�����ſ0���(>/���SV�Q�XRpLT
���������~�D�F�W�i�Nܯ�9�C��=?O*c�|N\^��3wN��W��Y<a]U��e�=$Ү�|J�a<���	U�l� ht/�}�ߊ�Uނ��T`u�4�3ι�"�����Է��r��">G�_Nҗ�3�G���\��n4��̿����/
NE�Њ�=��u	uޘ�\u�2D�C88 �k�������4l
Be���.���r���FVk{\'s�b"��(P�� ���9�im=��9�=�\I�$
͈��w��٦�8��t<*�=�0CV�˥�}T�-�J;����e�0P	/.�ú/���ᴣ+��Z��$�#�$�P���1fl#ӑA�V���.3�A���ЯEVٙsa�{\�}��d��<�p��Ɩ3����*^����RD�͙c��,5B��ٕ�+���"aalؙ��j����9h�����!ԴW�a˼�j�a	�Yw8��M���+|_ڞs�B<�^�q�;49<��D��& �>�����-��L��ܸ���u��˅��G��y����?=ƭo�g�P2wa�+���޻���a�R�*�O����ߎ;&I�u������V�y5�2��g�d�<@�����EP�w�7gNsr�ݟ���9T�iy�("=R�m��O���e��4�8B�}&�3%i"���K�eρ6,v�fkw7,A�,?���E�ʽ��@�٫R("i����K_\�v���eu��-����2�O�ċk��Q�!�v��5��t�r�z�6&K��o�SO3%fqY0��Ұ��K��aA�Q$���Z�ɷH��� !���S�	w{���f�8	Ue�z�,/�ߔyrȈ\���c��p�^�zQ��h4���k���-��QL�(���bvVb�a3��L�;;'Ձ�h�Cz��I#|�� ���ur�-c6�d�1�0@��0��n�� x��&�F���盰�x*�~�{�{R?)�
'׭w#; Ed=�'q�{ļ֌fR/���z
�g/�k	4�Th;KU�Du���.`#baLi_�/��Xu(��7+3�0 �5��4}�v$�XűBX��d�j.܈��Gz	n����Z�PV�_�'RxN�@#u���3��D���~��T�������*�ؽv|D_�kЍ�4D12�Zp	�+��e5/q%kW��������_b$,w�����bF� Ҥ~Tꐓ�
[B� �v[h�F��쏰��a>��X3!�U7�/d���8m���Y�<�ҫ4���`�
�,�"���H�{I�����D"���Ӯԙ�A�� �Z~� ~��}��Kl7%���]	��߭��m_9]�)�����m�}@�E!�6=Kψ���w'钖<z����Hy����IjX^*7 '�>ş�T���3Al�,%$�4��bP\L��sY�6������\е��|Gy��=�"���^[�h�ۛ�6�>t�!������1��w/��������v4{���*�掗�P����i�@��3)E �/�d6:��8�ٓkgFj�j�c��,3E"�ׯ2,ё���;h&u���x�?�\Ʌx[�e�CW6W���q��G�>a���R���S�Įע�?eOY�mX	f�ynI�Z>�L�h��I�Be�E)��Qӂ.�M:G�)�$_��"���'&a1�`�'����@�d*�#���oQ��(jC����\�1��YD /�%c	ӑ^N�63�.�j�!d�:g("6Ai�L�o�uJ&�U����t�a% �׉�g�f�p�4����<�N�A�����񘙻#2���7���aϴ x�<�����k�xa��	�W��ϴ� l��wX���	M��Z�U�1��*4���Bj���rN+��!L)�t��:"��y�}�����Whf��m�������O�Z�b�G.P�m4�y���V5���]׫ q�T7k��DÑTo\�ѹ������	.sS�_�<�ȩ!}�T�%�Bc�� �i$#����A�ǈ�f��S� �y1�MDNp��*Z�F���0�asT�Q�]Sm����:��j��)�2����J�XG8��x`������-(F<�BJ�ލƇv� AiuEmR8�� :�h1hy�$̬�
����I�h䧍ga�+�y'$�{���E�qݫRukA7�h˄���{��hC�{9�q���ӬH�?��l���;W�V;k	F��d�$G|��_p��Gr����5XT4�*��3`��g��<�ui���;�� � ��e�pt�^Ja]N�bJ ��ŏ�=Y���9�	;�����aZ�T�K��ˋ��U,jn]_L���y�Rċ�N��ֹ?��`F��	-Y���k�LУu�F�O�<ڰ��yIv�29����_jWW2Ko�Gʳ�6�i�+8D�����9��.�bGŵ�m>�i\�E�}$tB�
�q2R��w*~��'�YӼ>Z@!4��LD�p��V5��ӄ���Ƭ��aF�V�^+�Bޚ��LL��;�i�1]*�=�R����úM�nd���W7��]Tz{:�О����n!Pw�����+������j'���M��	��U�L.G
~�mq�D+P(���k�Ff;��Ψ��a��@�����	GW��+����z~s1N�Ӫ�v�p;�g�9+(#Cfp !d`��yE��9�R��tjS�p����4~l\�O�8�j6��xy�[�d7�f�b�VЋ���[�'9�Jt�2e�(�EC�@f� r` �1
�;lO�~t��l5
�0/q�7�i��_�:T���|��5�g�4�����ؿDY9;[3>�c�������������6�f�rH@�	�m<�{��{CL�g��-�� �$4`�@j�u��jF��v�XF���t�N�ɋ�]�ڸFy\���/��)
�7�� �#ٝqD���ҋ�����` uC��
[$�,�7���)��ʢ��!pOLE2S `��O������#s�͊���*n��{��Q���BW��DPrEւ�e���i�2J>������,�MX� ?<3ף͂������bS=�ډPQ�N�11�26*x>M��^An�|>F�B�� { K�)�ǫ���n)�o�8V�$`<͕�����@��� ���顥� �7X&Qb"c�Ǒ����`E��U@a�ޛ���Y�);e ��]REO�-�I��P4}~�%Z��-M|�z��'L�>�A�M�^��!�%�?1	^&�4[t��9�ͫ���T��q ���(�s��h�0�)�{1B.`�`B��|�ý� ��\f�-ͦ�
��[��<�_���|ӧbUM@|�L���IF���j�Wx�oS�mQ���䇀 ����.��qi
��Y�&[ǲU���T팣�řv�
�Ĉ:c���Pﭿg�7�<�R���e��yk�� �2Ǒ���lX`�*�2ʑ�LgE2���#Dc'�E4TF-��S-,�s���?�d�jLF�|�L�Jst�!�u`I��k#����{*5I,�$Z���C������;d4�QM]y҄ޮ������W ��^���*�5H�>78�D{m�=�N��mf�%~��H��y$V�;�����!�lYq7�u�K��s�i�4�?�5�9(�Y�i�m��k.n)9��ާd)��H٠����K ������Da�����,S���/iY�z��a���\j�s`b����v�f�)����d�}7�R�
5f��w���PD���P!'|�?���� �_�q��_>�6`GF�2s�Hdx�*<)X��v֥>�&�$P0���|�D�Lk f8�љ��u羥^�����ַ��Z�+�e��<Й�wU�<&?�
���sSCW���p��O��Ƽ����Auχ���[V���s�Q��21����π��.�:�m������,��&�i�����e�q?�������`��|�ӛ���}�O!	�Cb�э��"��ɑ����к��F�)�D�s;��N��H-��/��	�����#����Ǝs��#H�� e&$>�ݛ崙rQ�)��ͬ7l����g;ab9��Wu�d6�?�	IW�2ٴ1s���D�t�U+o+K�8� ��2��	��;��C�=M�'4em�z.�oP!X<;�#OUO���_|���*s^R�D���!\q?�*�j+ݹc
���<o-�:9l���<�K�0PvF����bL_����:�C�.����A��耰��d�a3�B�8���	<D
Q
{"'$	z�
y�}��>˱Z�b��B�X��|'��E�dt��>ȣ���� J�𣯮���w�#�u��-�!kU��7;sǧ\����=!�j��4�CW�TZ��C�#����K<�o�����M�`��3���XZ��#bӻ��cU�|8�Pt�7o�?o�M����@xd�*��>�4h�.��m�5����8r|O~�헦��5X�Z;��o)6ǔ�;�{�qǵn�*��J�Y��,S7y��]��x��Y@����`��'&��J�nM�K	뗽z�1�����PD�2Xd��
����3,�a�7��	�g�����J��,����R#Ϲ�䙃�eQ�Dŉ���rCjef˃���Jc��?_�爁X`�w�?Y���F{i��J�=��J+�����C�!��2n�'Y�q4����A�Ɇ�9�����|�se�5�����V��!z�ٿ����O�����53c6����O��l��E+�7@���v���ힽ�!�k&�5�=	��j.l�������h������;���a� SA8뻗����1u�� �a��F	t���`����H���m���v�E�|lNw��H�ۀ�bd#kr?.y$��Wv�{FsN7�\�X���:;d��h�c���̥k�Q^w�-�|>�r����s�9���g�]T�ظm[���iv�OD��%��y�VW	�Ez�%�]�?�m�DƐ �7���€a�8�X.�``��Շb�ݵ	L�`("̬�f��n�$�����L�/ض��q�7���h�̈́�Xa"_��(��m��8��Zޠ��n����s�����*���
bnoW̯Y�'+���c�7Q�i�����*���K
JTW�ԡ  ��Nۅ5�S���o{)����l���xR'
,r�-R��h��\:��`,��at����Z��n�a�ʏ^"D�/c�5j ٧���ߞ�+�I��|�(����b����9��\��&l򨖜��75�o�0+�계�������-D�&��0�#C��f�C�X�s]���N���gL���E%����s_Ŭ���L�n��Xo�����،0��/M}d{�F0�� �$��e���2��Ua��p�e�Ks�`��( ����=/������֫d�.�2q?�Kd2#Y��_��ó���'Ɨ��p;��R%9y� T�(n�)�S B�A�M���QJ(DLZzr�IX�O(!�̔{#cѡ���1�v�s�EE��Oz5�
�v}[�i� �aom�`*3m��_;cW��T�tx^ǲ�<�Q1�A� ���	���b��S�UeO��ۨ\�lbޅm�TP�h�|u�Z@�@�(�}���'{x��vٓ�9,넇�{:�m��7��Y��t�e���N�<�A;���Gf�~Ѯ���?7e�Vt��r��/�k;t�	G�����r���Uf؛���-���,CZ�>��aLd�":BC�oc����  ����g�j-�D$HT�i�T���o���!��hb�>j�K?�k"