��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\���V�fnvx��ÍG_;�ȅe�~�>���9�>��Y;�0GP�5����	$��������6�3 �Gxx�Li/�(؁O�r���/����a�9\+!�gA�\GwO]����jR�@�Z�2�S����9]�~U�*R�
J����#5�퐂��(*�ٸ�?���4�^�l�g��o�����Id��)�`I��
@x-~(C��uY�[rr�s�jg�?*������^;������P���xT�u���Z=����75q�D9�g(�*,��^>r�� 1#��ڬ��l� x;.���9O�ߝ<����L:�8/��0T�>|��m��ݥ�kh��
�ҋ�!z�άH���r�tk�Q���z�٥��9^�4jW&���gTa����kVoX p�s��~�e�R�Y�����T/!���0���Ͻ��I챖�dC~WO:��}'��v��Z΃寖�}*g+*lCYg������wvkSiU}B����H|Q�X�s�qxp���=��o(~�cLS	(ֶ>n �����󽣠U뇓��<���.n�v��*S�-Ԏ�����l`p�T��9AuNx��>��|��7�rW`�͝�j�]�ޝwYRU+:/�q��T���9ZkG�pcU��X����?�Xȧ>� �w!�ߣGj�£�������i9�E�̌� -<��H�:'�b����VG�d)k���v}bR=�F�
Qd�Gp��AٽJF���Ls���{�ֳe3 
�َ��]llDJ����*�[�M���~ޱj���X�|1̲��K��x��h���
BF�t��[<BtdEjfU���@2H��R�=�(e'�oHg9��۶��
@���ӝ׼�avYn���|��1�Ŗ�Կ�lȇ+_�5h=�@7	�C���¼��k�X���3��K���e�1O�3vqZ��W8r1=~;bG{ԁ��64�ۭ��aA6�?]~�p*��qK�o.]ԄK�ed�[�ʮ$a��|U�ƛ�^���e� ���)~b�����a�s�Tsh䅹ٲ3�;Ɩ�y��@5��"Ο���v�����{Ԑy��R0�JI}d�5FpU9q�:�{� ��\e�J�ȹ
���Du��g�/[�&-c^��0��ٔ��|܇�I�|�7hƿ��mlF<�ςւuWAՐ�[����)��;���t�#�����w�oP�����&��n;�]������.�c�V��l�4(��A�)�-Y�5i~�V܏9��?���&�U�;e�n�O^��c���aɗmY"}�l�oQf�KQ�}-Y��Uy��ٝ?� �G ���s�g$>*�Oq\��v��5��v@LCzt�^'e���[O��ͦK�"�<f��:2�^)~Dnk�?�ʏgfn4�i�����ڪ�L�J���(���j�:����.*���R��%?I*��Khz���������K^��5�&��4v'K���f;������v��v�I�x1����>�}�וUcv �:wHE}��Hs�^�+F�9z��/N
	!�_�W��~16�nXA,t��|:,ht��5�e"�2��c�p�Iq>�9
�5��0;Z���F�eĄs�o۴�:ΝE|;���{��F��Uޙ��a4A�SnE�X'@H�5�b�3���)�|k ����O~~%4�7�)�Tʌ�ޢ�4��!Gb����Z>"/$�D���m��ۣ�*�BD�7���8�:�*S�$���q�%x8��/v�oQU�1�2S�(�uoo��3֥*��Ew��M�=��N�D�%дVN���J�HW�2�^���P�}ʅ�ӄ���eoc���Ӷ�k,�:lr|�G+�>�~��Mr�kX%��vh��_��H9���Pi���8���2�o���ٜk���X�z���9�� f��\OHh|�6F��7�{�i_�eaڅ�� ����v��ep�zI}֕��0��Y�~,L&�a�a6����#n%��O>������)���O��� X�	qXM^:�@��Z	���2�Z�� o?�0�+p�P����=�G���gU�b<�u�m8(f_�Y�)�a$Sx~�=�'��0XC� ����(^-��4�t;Z�"Gn�Z�4��vւ�j�%hb\u?��xrű��8����R�� ~�	�gx�Zi5�$��N�x	��6_)6W���"��y����� ���!��)J����J#s͈2�3H^`�3��w	[�>yX��Ӗ���5���呚�Ǉ���F��u뫿ylcgV���9�	���\�$��x["}��Z�aEC|(c��>�L�?��vD�$9���J�]R?"pý�	�r�%	���x���X-L�G�c���wQ ݎ尹�Dv�2�#�6^j�ev��j���M�������σ���:|؇��技-�Z����/v|tA����zD	;�7{��ml�1�\�,�o�2�8�
�ghR�PL�J�X�(�z�����{#�^�~)6�: d�"8V��2���b�5�1� ��yLGk8���fYMU>H�1�q�х��Ѳ�UDر�ʔ�ފ$�8�x'k����)���!�����f^k�V�C�Π0n����j�;����)h�膁Z�5�����E.$Y�?������/�K�~��d���O��"?ƩJ�Q��<亱�|ڒ��������J�ͥ��a7�G�Ȑ�7����C�N�R�uz�,��O\��B���C®�U�dݐ��-�����K�^s���\爋[�5��S̐�;)G3��0�eg����S�C�n(�g�i�Qf���?�|o�]z�6ă�]�5���v�*xx�}yx*O9u������b)��	�}��hY�3�y�EN�>x��S1��{����w�6�C����K����&�Wd��Q�-�J�V➈'p��f�m)P*a��2���oT��m�4�Z�[�Jgod艭8���ܿHL^��~},�&�RT��mY���`�O����5G��S��b7Q��ոn����2z��!m��_�2���K9�S[*�����)$�ÑC����	���gF��l�L��*A�4�օUY.^�7ޠ� P[��� Ci1�����ּ�����k!���.3�P���O��6�C'�s��Xw��割����b8t>��+|��f�ws��9H��)*Vď�nףq^�&F��a��@j!.�B��/�Y��s?k���������@��[��tZ#��v�rY�A7�l�t�)�Q�g��ra�e�G�z2&n���}��=�fx�~
m��S�9�0L��ZQ��.~ĜUfx+p��ea�^�~a�K�i��\d����`1��f�L�����8@�u�����/��@(s��.�8 Z>��p/�DA������H��V�s4=�o��;��>wQ/�kǦ6n{v|<쏛���S��k�L��qDɀ�c���>���Y��� _�e�|S�v�j�ɼ�6�ȓc
�;�h7���0%^%��������5�׹���7-��S���Oi2h%_V> 	�5�!u|3���2�xs&l���ڈh�(�k҈x_�̃,!!c(��<X���E�"�If��k�cے��	�8�cG�:`ĉ���i�tnk�a�ܹ0�MtYȃmޜU���'�}��P��E)1 �1�f��l4O��._�Rx�v@$��v����N\�A�uv����R��N8�;�@�o�\.(�!�ء-Ł�>�j*�Td*WN����䨟�b�â���)��E���!.k�Vs�;�6�@Od}�L�K,� c&�{Oyˎ��N}�r`��������6��+_$��/����V��h"՞	��;���d����#��>��Y�i�I��Ĝn�%DQj�	F�g�Z��O_�K5UFXM#,:t��آ�b�:V2���|Ȅ��b�.Z}K$�3��B����Uz�f�<�H����c�ʍB��AL�1�1��rE@Ӄ�D���G�y)����2�]#������&��-��E�s��u�ēۃei� ܧ� ��I~����{a;a]C���l���E����u���2�ԓ�@���_���[X�yA'����n���� X�ə��E�?qU�"��uLr�@�۱�}�T�qa��_�S��	�J�E����L�#	�]"=�����`P*�Z�i�?9����������5^{M/���ޜ˙����K��2���'0�JM���D��\M,Hŧ��f������E~�ɲ��5ȟ%���${FxL.k��J��8"�Hf�����B%�d����X�✻2Ώ�b"�+<���(&�}ɠ�(p��ʀ~Dz�ߐ�u�������f����3�|\�r(�����)����Rp!Yj��J��⏨�hK7���`DO�����/��%�\��É\%�Mx��1��e��'QC��߀K�|����{���y+������D�
����/�^�y#�X��`WCxډ{/)$wz�Y�3����}�z�O�P��a��>j�	�cM��JjG�JH��kἄx
]	������m��"z�,՗�e0���OnnD��%�J
�r�i]��~nQ�W�ћ�;�i�2��p�p�t�Sb��i���7���zE� <���ߐ_;���n���<�7?�"�z� �������ԧά�ϡ/�vQ%��-�V�����c@�i{}�9N���q$
�~e�π�C��&�M!	
2,i��޴&��ؘB�J7I:���GaB��̯���S<�O�sl��R#Zv���HSrO�m��#��Aq�1w�Y�J����A��a���{�w ��)�^`���I����fXF�nr�8o$	��0�n�].�6��4�'�x0w)J�d��9iQ���;:� D`��+��K��nZ#M�!��d3��n��9��"g��X�]��qAH�M�}�-������2�HqS�殻�W⦳��X�P���)�����Q��q�U��h��B����E������Յ���K�����Hxs#�nW�G���*躹�Al�]�(H�r�W���<�	�ds��rPi�aK���&	%�!u.X�\�/�'L��ھ����V;,�ȡ�P��:����ۺkb�!�OLN^��e��G촶��ԧ-]Bd�^��9�J�?\ב��v �%�I�	�͹NNG�OpY�}y�sr��H��ߑH�n�&��Z��ȣ���5[�������8���5ռ���>	��dM��"����w��)�v�eh�^@�	T���cP�@����M����� 6��f����}�+�,$A�\�`�4�$uo,�!"�x��'I�����ς>���ܧ��MX�yO*O3�z��a�����G�`Y|4���_��V�[�"|d�THj����	�Ե'�T�۲j����*bS&�]�z��|����d��R��UD���M(CC�Lr�.O�g(�Y-��H X(}T�i�7��i�_�w�W���÷�N?�*�:�lc� j��Q \�޿�0c�X/������mE_$�4�JΛ3b� Ua��SJ�I
3���㉮�<T4�n�v��9Ƙn�TΘ�l�Õ
�	�gn�i��広���w�b���v������^����W�qi�������?c5�\�>=t��U{�.���ܵ���b�io����l�gs�(�*a�9k(��{y�=.��@h�v�Wkh\=~�l���ڿ�����^L�]�M���{��tW0~�(P(��� r����8�ZYR�p�QR~���z�M{N��gXBHu�z�W.����L�}���j���]�d"�b����/�E�Cy���/9#�_��t��0F��f�� *	�bi𐳄4������KY��dg�[P(����!	Q�rV�3��1M�C��z8q�^jm�rj�n]�MVW �%O �"�����x]Z|��f�V5�Q�0.8�{ �J���D�\����_y�&R���;�[`�{ǣ6��]���?�~HWdX̐��z'�ET��ν�ā�j�(P�.ʿo�
y�i����*�O؊a�Q�MSCA�Yec]��W�U�ehC�5P�ةL֟,c��5���W�"�)%l#��?+�f&�a���:�w�I:-F���"v/]݀	Q!Ͻ��dF�oƎZ:��e��[ݮwTyv�]���� B&7��Ɉo������ 6��L�����%~�qA�����K��Ի�����K��DA��ݡVϹUz�S�Ö��9B�L�|�,h�f\����̀�>˜��u2�M�����`@@r�*\��Zƈ:F�d���
S��aL�	��sI?To����H��������sF�=�i��')@.�=��'�������)S
($��w|v�����+oT��32��"�H�4�"b�eAT��&��(�z?�ɴ�dM���#��04�i����`��?��Q ���W�Y� �����ඤ���U���5 ���j}��־w5�����l�׀�qW���{7��Fk}���E� T�#N)����3�]m�8|͋_�)鱎�q���3���*B ��S���T��R�����D���"D=l��ѫ�'S4A�ݩR2v�,�7��l�[PX�A�.�JP�iĝ�"��W|=��q'K'�����5v?7��m����J蔒s��g�+Oe@N��ii��}�}ʸf��|��V�U�9�	����hk��W����b|�<^,���H]�	���q}eʋX �J�}�����x~8̩�o(�M��zE.����&��XJ_
���L�M΅,����׫��ѝ1�"W4���;V��Ni��p���K*�⎺"Ci/A.�?t���m�6�`�u���,�ڍ�J�F�g��I1�%�9=��	�b*����$B��԰���v�(����Y�����	�
z`akLl�d���le�j�M��Pi�J}���F��g�~�,�lGiV�*Q�T�	%%���g��u�8uc��E��ǵ�z�4O Q�,�:
����}�`S�2��WcK'Fn��=�Û#
��쏐��q�\6d��[1�[E��3��7P`���F�g� �!��;�^Ѩ�y3�g{��lο!3���*t��17<���L�[��Gh�(�+���e�"��s����b�r��M>?%��9I�r�42��| �B.*�KE���1f�q>�|��n2�<�Qx
K�5�w}�J�^�b��_��C�"f�=^DZIwtQ�.�98N�����M�i���H,P��?X��aV�8~lsD8�Дk�mP{68������i��11�f7F,�N��D{���==��%4�!r.�����'�U��
�R�X� ��{e���j����}CJe�[~Iὠ�-�E<u��~��2��Y�,Y�\NW-���X+L>�� /���Ue�T���z*wx�8�$�i����sզ�g�`�)�i- ��_d	g\ƿy���hp�}#2Gp�����L3�%��I��msG!*	W���$V��q���[�P����RhyU�Ơa>l�%��m��/��`��~���z]���Bj�q�jAh�����e�8�4�� �g-oI�ә���[?eO��n�-�`5q�|My�~擧�����Iɐ�I�vA0a���U�j�a���H�� P7P<�SD�,-Ue�a9��!��H�B�8�:�@���X3�#mt6��#�������\9�푨�T5�2g��Hc(?O��e�5�p$�kR������
�"����	�����3���=\`�=����\-UD�cb��.��S�Up��A�3�#L�`9.ŝ�
	gcZQ��*[��}ڗ�v7D����u3��E��i�.yWL�W�}K�:�fx M[����Ø,+���K�N�yuǠ ɮ`�<�Y��7�E���-���ٍ¾`[t<+F�5��Z��_U�t_�9���M��,�`vAڡLk�$9iT��W �M�R���>B����38s������B@xi4y��b��̈��c���s,��"��n�����n�A|���v�}8��Fz]��Rk'V�>�d�$ܞ�⍐�s =.NS5[��v�����՛��Go'{�2����e��6 �l�4�YxQ�&X�%�,���1�L1,i�,��r��@�Ӽ6Ļ�?D�0LY��Đ��"�Te�8I�4A�(D�^1�?e�ZP�gwױ��5C'}�y�P��$�@ߥ��c�������q����al�=������ZQ)�y�� g��Q/���5�k�&���D4�
��ˈP=��\�}G�_�7N%צ��^"=�e7Ӻ/z�E� �>�xh��Z�HWf��~��O� �9A�����/՜���\��V^�}K;�A�R�3�]��woa���)3�ُ;MF��4vp�ސ��Z�v�.3"���L���\ˠ�G��C��)� uk-2B�CT��*�m���!���D�*.�����w|��*�}[`j�!�d�P�'����s-��K(�<�����>��4�iR�_�e��n@=Hs��+���L�����ҷ��KH���5A$*�ı~��<���x��7/�Z+����v	ɱ[��m�,Q&F���y=����k{t�SƧ�����XjZ%�cQ�Z��U{e��{��d�d�!{J�d|����&5�?9�9N�/Qz�H�7�G Q�D���@��=��%W^�qw��~����j"��"n4�%P���z��E_FeM�d�;����������rLh2>{	�B�i	:k�oi��Pp��u�_*�'#�"U�q1���g����|6�<�{�O>47��b��g���R}{�LD��e��]$��<�D\(x���)�'.iF<����X���uDN	$Ry����a�&���6-0:���)VF����*�ܸ�Q7{�>���=��1!��d�s����R������?�!�T��׏�������R-V -3lٞ�hܠ���E�3>��'��y�}���ۀ�����)	���^��k��P����(I�73/��N����Q�M /��F��{�!_�Z�Yނ��]ru<rH���8?�z���3R��e�&���4�'G@��fS�M�mK8���%l�o(`=�S���q2R�<*�)c�:�5�D�z��aCw��[�s�lE��9ޑvO�`>�*e+��%`\�l�^"E�M齜�ڷ�J��#={q���) �OW�ȗ��8�7Y�C�v��2J=����e�J�X�D�++�A�E�X��`S&zGZD��Q}<�Rq���+9ԧg�AX�mRr�p,�5Z��oH��Z7��6�DL�t�eW�c�/��%*��q�c�L�^<��vH�7�v>3V�,�*ZҶb�&������Q�(������!-c@���{RL�'n����$g�&C��ͮQj��� Dl ��M�g����t-O�n$-G�\;�x�����+p;<�@E����&9��B\U���Y�`�����"}�]�2�� ��)�qQ���ǫ���O�?��&y|���l��"�HrɗQU	��y�9B^�V�`�N��|�p<�B���qVK��*���ч,b�t����?�s�?6`�E���9p�V:�h�
�0�=�D�v�0h���at�x)���ه[%�i3X�
���aҜC�ڰ��Ը	�b�k'ҳ��:��Q%�ë��64x���ZY:c�5�or�2������+{�m�8yd�)G�E�7�;^O@��*��0{ﴳx_��+I6B�+�_��p&�d�l'ъƨu��&{L<�lĽ�Hn�PAQ8�s�~a75�!�E�������x ��l�t��?��aI}��NW?�Rfj�$C�zC�Q��烞�I�V�BA]5/.+�e�ա��M�������92=m"�|�"�/nÉw�Z/�۩c�  �O���� �D4T�E����(Ԏ�r9�c�O���թF�뷶�V?�@�N/�v�V�tCz�@�k��;�:b^�[Ik6:�ig>��.@!��WA�g��D��7����xi�8�����a�j�+DIJ��3�c�IN�b|�#ԕK)�^�iLJ���pH�>p�"Sf:�z�ZbJ�oo����o��8ׄ��?�^����,���&*$e\�=p�&D�EG�ۊD2�6��I&�f����I�~�Za�rLB��4#MЫ]����:�R�0r�G��.�Ӕ�&����(<w�A������=�fϙ�I�8^�ȎMy#N��d>o"�_�f��c�h]�ۘ�;.�*+� ����N��r-�F6� �-y��Z�'3`�J2�Z�����-����ݚ$Bؘp\�Gk�Ȭo�e��0NJ�,gy�"Cl�@���⣲�ֻ	5�^Z��?Z�PH}�&�F�����UDlv�P ��U$j5ݹ=4�2|�`�e���'�<��Ma�Y5C�7nb#���nd
'`���T��ɥ�t�����%��1�h����9�8$ {����j��_�߽1S�W+�p�l��`Q�<aKa)�6۟�s��ky���	J�x�gv�\%#�pʐ�5򯣊�Z�_��DN�[|'A~"D
x���$��ț_ֆ�(�cU���R�����=	2�(T\Y
�pQ����0�3��j_�{a�2 UAq{�PF|%��� ('9L�B�*���q�j9^�������D��.4�r��k|=J����ׁ3��)%a(p�U����o����/���$&��R������R��T[��&�`��f��I,�[@t���d�Dec���(�Ϫrg���S�`ݔ���Tv�OI��<�~%�!��(P?@�W�U�&�(y��e3M�A��5B��w��l�ST%��Cǩ@:(�,6R6�Tsg`B���Z�~��죮�Y_w��9��csa���b��u�V���HW����m�����D�|0o�@͚��cK5sT+���lX1�t[R�vo��T=o���OrE/�*�ѹ�ˤ!�?�� NS� AD1�Z�ܑ�'��Ʒ�sUMQpw��o(?���
d�n;�L�;AL'P�UG��0ybx������%���E��Ϊ��Z�L�3���^�ZW�f��A�YYvƷ/az$�1>^�{��s�D��}%�I�~G��>,�.Q/��%�?i�-�]�c\aR*�-�<�?�9i<�7�D#�.茏��������됵�y�=����m�P��y֥ޯ�$���<Y��ɚ%�wT��kgk�TB!��p籜@��� �����k뼻���6:9&ޘ����Oq�#Ev:Q��L�IG(�ӔU�RcF��^H��h�ãg�C�;�6��x�՝�o].}�"����Z5a]δ�.���S(?�ob0��mi��*)���,Y����zlt{��ri�|�{��1U��(���VZ,x�
�w���+|�1��%}^�@���9��m�N ��,Lei�Ocl��-�ۤ{B����O�L�N��o�F��r��� z#�-�nHUc/�nR��b����_%���<O����RJ3��V\I6����]�� /��='�������@����(�^��?�Q�>;]�9 eX�nl��~�.?,��/DT�(�������;J���c�AMsΏ8d��ˊ�����s��W���� !��H�h�&-J7RDo�%ӳ0�`��{U�xͱiT��;M��=|��Re�n�D[;�Y/������M��Q)uVc.kGq@�O9A�����~�s�Z|d�D�2���BJ�� ��v"v��Ԇ�'d�G��R#��d�ڟ��n����7��`���X
��'�։b�jV@μC��č*e��'P���"k��sUG�"Г��_�VJK��:e�x�}D�����B;Є���1+8c�}x�f#w���d������V�3��	#(��:1�żĿɬY��T�]�NUv_fGG��ܾ��a7R�����Ӓ���-��D(f���J�H��&z_ J�:f�\�l鲾u��4�Uv�^��4�&A�jܬ��v���!��� R�#���d���&h�X��:�L*����)O|�ND��,���}齴P� ����֪jF�	%��@6T2�	H󜘷\��,�l���Y����\��F����X���V����mG�J\������^v�L�1vtB;���zC�ژ�+��j)�n~�-�E�,�w�?U�i�b���[���=���(t.���V���vW��tSn�AI[��
�t�g��^M�۱�����!Zݚ�}o4�:,�'�u��ۃ��h�4|��k�<m�o�n籄L���{�wg$��<�r>�VҖ��8��e6Ϋ�O����\1�9�XMf������M�/�26�~�ʎ�Gĥ��`�9�/����,"��M�WR*j�H�*�	��.�;I���WP��`o��9aؑ���Z��}�<T�r�d͔��?�c���M�bwq��
�R[��u�!�CZ�8rو���b�R��_����7�UP];�ʔ����}F{W%�Bo\�& �{\5ma��\����y�VI��{�� ��h�՚����Y*��4��H0����<�F1�����=9�6�>�u���G��0���ӈ�Vj6�c��JW�Z%��vn�}N�E;�^�ǹ"��_!�ԮR5�l�.��,�G�j�X�	�{�=����b�k1���~�*7�E���ݎ6�VKú�/%c�sk�����lc�/�YJ��k�å�_������*�VU�h9yދ	�'6C����T������S�7��uWXL��3��;�܂kb1=pRy���oB[$��@t�ҋk������}��Hā���u7�Ӫ��7k�9��nT�	�dJ� 4!#� �u�����|��fѽ��g��|�,i�Ը����EF��T�����Z��O;�Q�}����X�ָ�V���*y1��(����w�Zr�y��ТIxP�ԀB�6!��?9N�Q����Esi�j㏅����zQ�_k:-p����r�x�{5	'2e Ec3g�  ��Ir�G��/���-��.������I6kǕLݷ�5ϽÈј�$��r�(Ʀ8�WN��DZ�pfDt��U�B�>�s��VW=�0�Q�����i@�(�g���
�oy9����Y���+��&��� %��x⑽�?2�~C�Ūk=�.�tJ�^�U߅��*I�`F^��T/��D��}��%o����#.�{�����ʅ�v�z�m��띞��������d=�g�c�ښ��¤3��$v��A
.���Q�c����)�o��T<&��h-"���jϯ�z��F��6�D��"4
�dՅ���㋥y�G$��v��Z��Ȝ2�TrCR!��H����P��*bR�f0��*
�*�ϹTK�>Z�X��Z�|�&�]e_�%�$3���^��]:��^�2�e�n��"���E��(w?����Z�lp�	��I�ױ��m��]d�ժy����տ����˘����
�-i�V�S�5�Pծ�`q?u�T�r�O\������`6���M����kU��r��������M�w|����Z���b= f���gg�"�����M�z� ���k��;����>ԋ��X�0�x���a��5?ڠ3�#��%��>Vڤ�++�� ��/���Hf~��h��M��'�12_�͋�H"j���;�t�������+u���Q<ll���9�ؔ'��jA���@��o�c�gA@-�VL�I��(��`(��	��� �76�<s��ߜ�^�EN�Mո�1������2��>��Q����f�գ������m��#��_fO�\ɸ�ap,��Z�����j��-�sJ���F��|`�����hT[֒4��a�
(�4�Zg'I�B�%���ɶ�ؿs���{��,��H�Ƿ#��PIk�P��!e55|�#�i d��n?�L��4��z�87��]�����k	O�S��{�ұ�����vqb�Sh: ��6|P��F��ă��P-�b*!`E�L��96����xM����YW�:"��v���~�ˮn���G�%�z���Һ��v��8-?@�\}�M�p�W�Jx�t?'�Y��5t"��?Lf^r�U�\���.%V�?��M�ԣ��/��ǜ�S�S���W�'"cx�R!p�BWD�_�S5��s�~/ �g7��J]m0$��q���;���F��~�5x�[@��G���C�@�;,�[>+��e.�
U��t��/��ҹg8�6����4����x,� Q�t^�p<MQU]-Sdy�ŧp�.g��F3��'^�ޅ���\�bQ�ff\F���^���.��j��ֲ3U���~_�3��D�q�'�rl�MKs f�.��BV�	j�\�I���n��C�Z��db�褶�/�D�P\zVTv�c7���!��]1}̀F�E��	<!c��P�83N��������b�<E�$�W0�M�Y8X��M��j7��"�I'����ժ�R;i=g|yp4�B�[]���Z1��oX=P!dʌ�|��C�d���]�}��gLV�w�L�7[d���@�������5M��u���O,A��Җ%&4����^VẸM�ꚠ�?�a���v�Oɾq.o�ST4�"�w�#�~���EZ�e��P�	kԐWwc��T��7���sc8�!]'ׂ\�<�׈\�rJO�W���
_���U���i`������
΄`e�>�jz�Ņ쎰��k����v}w�a��U���`v7'3�o��,I` c�!�Ղ�R��;�\��������M���&����Br���La	9O���ݒ��E���D̠��;�[�`b��7����.\9ɻi�k9����glx�td�(��I��=q����2�κ4ؿ�j%�'X�z��>�H��P�A�b�"��ܡ8�ؕ1�����>�i;�q�FwPA``%��%о���X�̣��E{����P<�Im�i�|�=���n�s�XM�fE�8�ʒ�t���1;O�;G>ښ����/)P��I������DL��$HWq�YmD�'�}l�wʡ��1h\�~������18��/F{�������hmr�y=���l� �
F#�0�xm��H��i;
�Ȓ�5h:�B)�w@'���U?�B�=I�g���cӨ�k�rU���_t�G�x�6��w�˱1Jn'jq ^��, �������Z0qS·eÈI��r�0>�� ϬP?�;a2E���K3�<���-Jo�c�
;�jC�n�3��E�[��'$��SW;���y�J����Ɉ�qC�3��*!�1��׃���5��oEU���g�L_q��yH";�L~���%�$ӏw���F6��z5i��q:;,�RY	�F�I�2�h���'���s��� ({I �E؛+�Yomq~�,1+	B��[� ���>�$p.�@�@��X�D�me��Tg�<��d�
uq�9gm�%�,r���?8�Ҽ���^�rLV�:L���A��m�P����P(N�@�b���Z�GL3�~d��@9�� ��띨������Q�����]렒Fu1��'�@1z8׬PlL�Q���$(��������3��,��'�������*������Rć��V �>��:��3OqpOA��*�+�+k䚀�b�W |RE�[k�b�Mo�U%%ҼE�5��@�d���U>��|���Q�~P�����g�o��{u*[o�|����.T윰`�T���n˒;&��I_ځE�a�/��8�i�[�%��A��"���o�@���ģ��4ʝj���פF�U'��/Ě�x<��TU{�&wۂ��T./\n+�ac+M�kCP�3K�D;M�|�j�d����O����6$h'��@)�"�0Y�_:@?����ɣ�k�w	��#T�g�P��0L΋m%w�}��C LS���9q���kc1[mj �#��X=����KS�!S�pnY�|�J����o��9C�#��=����5p*�zw"^�oS���o�ϻʤ��0�*v/��zNg]A�p�f�hB�iv��Zdt�!�0O�7�.0(w�l�+���7T�A�>��bQ�ru
�v��a �c���	h�o��'V4�.B����X���eS�B%��t����tRW뇶�[9�*
p������5��4�U��FΪ�O��:#}��/l�hJ���%h�����)�]aw��g�"�����K"��/��JkG5��l$#�Vm'v������"Ȣ�Y!a1�'�+r�4�<D��&ZIzؚ�w|�+�5��9�DncDY��qV%�Ui�Y�[5�l&{F���Y��%|a���4�#4zkb�ĴS�m��ك_S�&�9.�=��v�������!�s����w
5-+�j�ކR�sLn]A\dU���2{kԊ5K�MT/_j���"���% ��~��k���oaM��#!Ɉ�K��_����-��$*�=#�v\$24(�V�TJ˱tR��8���w��L$f�q>��򺻯�푒�5�Fqň�-�c�?zWZF1M������R�������Rw�C�����M=�*4�t�����%'Q|9C0h����k	���:X���#�� �P�a��� fڮE^JW��#P�/��Ι�C?�x�ƿ�V���n�i#/琊@�CIV������o���uT�8����k��_M�o��З% bq����g?�8F�9��0�kz�6�L�ufz��f�[���#J���e��!���"'_�1�A^�˫:�lx�ΑG��]9�*w��6���t�=��e���'�]C�Hɇ�.�M\���Vɐx��*�۟�h��#��U+�x����k7������z�r��s{�Pހ�?bϚ��Y���N�e����{XUp�U�ex+%��;�0VXc��X��{q�5�bǵV2S��7�VBI},n��ke�����l���"<v�4} V X+o�T���r��<�EJ5B3b]�0�i	��z�Ӿz���@*�R�[�7� �'��&5��=E�������̚��Kҝg�Z�;��>�kˇ�>�Au�d������tɫ�Y�YEA䡁b@0~	?����^�b�k\+ӈ���\�ɐ{:�څ���e�C[�0�3�q����V���I���G��U�5/Z�Zs���_��=�s|ȍ9��q��� �2��8q��qL2*Ȑ�(�w�1f�q���r"�̌�w0�k�܎�ְ�H�8��B���m�>�&�׉܀����DV[+�5���\���JG���Sl�m�lةt�߹�7�A
i�@�Z�S:��1	�6u��	�e���*��V*/�4U��[ފ�6��ҟY4��Ү���r5�8�)��8�����J#�dkv~�G�M�ӨM��^��InC}�.���������b��{���Fo�Xی�漀v���~bYifL�.C[G&��zD7Ս�z�
�i�����F�@��P^�㲯���������A���	����@W�������+��e(O0�(���ҍ�"^J;�����5@��b�E\�4���7�y�U�N�����T���>��7YX .�!9�"$�sp����r�Y��:���j.�ַw�K��eR��7V��x�G�˘��1D�y����΀ߏ�z��O���$-�K$�h'Tj�&�,�p�rm��H�S��q>6���U�>�"�-�D��e���D�c��/ӂZq��b(+�hqOΐa�x�-u���A�I0�b�*������/]�E��1p��<��>���ur���4��Xb1�;.�l�NJ��Pnj�~)fK�0E��Ǒ�����rJ\�э [�<9O�Ĉf4��`0�4n��>��i�U4Ք ��Z$�o9��)Ts*��2����ۃ0`��������B���5�ì|Ы��@��`ɝ!�'C�(��:�J4����fؾ�L�������4���U��������-gp3�mU�M��Y�hE��iZ�Z~�&�%Ĵ��������)/�#:`k�|@�S��
�4�d}�'���(E1&�*|�F9=���R|U�#�N��#��+NS���$��n��aN��d_WB�:�JH�n�A�[e"��_Gp�8JP�"��s�|;z��*s�e�r�1�wX$�[�lY3)��� 	B����ES�6h�� e��A��g������\p�P�0������JZ�yS�pi��č�����mj������a�Fi�8-9c�����rb��j�y5�(b��_���;�R��l�ݶ"Դ��Z2���v��S[�ˈ�(�Ԑ\Gϭ/�;�l�$_�"8ǃ	{ݥ>+�K� <����6~���GpyZ������[�n,t��M�*pRei��iFݡu8��$ӳg0��>P�78^ze�hݘf����a?}�CZV�ϕ�Ù)}R6�=%��n�`!�'LZu��Ⱃ9|�?=��,*����K�bk�Ѡ@7�(;�SJP6���-�Y��v9�����|�Z�k]973���:���F#������y�s�
p��{\8�7���j�Ⱥ�@۽k|L��a�K%%v����g�k�JK�Y��v���Z㋗b$,.˥`��_����}8����Fk�y�nh؝��u?w�(/��p��j��h]j@�������%o+8ܧ9馄�	�u�y��j[?Ơ�}.�>м��'ĭ��ZJj��}=���j=�d^�	��4�B��  ��D���X]iRI���w�R�����4=F�7	�:��q���p�>����΅�a;�S�e+�4�ՙ��r
g�NH�B
]�;5��X �$ݟ9��|���W�L��s�X�o����=	�x"�b��7�&pm�&���a�"���Ɵs��w%Ą�^�O����qb����Ů���T�"��'��O>6�g�x�'p����o�ʤ��[8���S���M�j���
P-�xi(h�p�z���5�7F�_{�%à�X�VU���f���UXȮ{�h#K�����Z���̈Y�����Jl/�^c�Y�$87;����~t����q&39�M��Q��+I9��O�v�=���M����B4�Z0��aG�a�7\�����:��1������_���&��aX�Ai k�6�gNxs,L� ��ȑ�L�S�
�qS��$��2h����Q}y5<��<��0��B�8
񫕵��ա4P�v�R��B�'�lO#s�P7���n�\�T< ^�y:��?���j��U�Wq�P�.(��#w�Ȫ]6���3�&I���=�kG�tf8�h�^��{��9�)fa���Cn�<-s�3e�);����ub���=
湟z��7������jw⧒.䃅�­������:���0tF�2̓��YP(uz����%�M��(���,�{�-�ps����y{]��QW����L3�r�o��N����G�x��F�߳bq;����֚��L�I�N��!�)�g£��@E�K�AC���́QK!���?mL�yjJ�&��+8P�փWj��%�xr%X (q���s֭�I䂜�j��1�,K�@�H��cҍ�6o�?�v�/>�ӭ,q��G�d��4����D�Q�s�۲,n����/�(�t���=Z�B��;�7���m�HL���WD��eA����ݽe��-I��n{dH1�x��յku~&� ۴t��Z���7������=�g{�&YJ����w�=u	���Ȗ{u�ŨP�h�eV���Rq��4�"��^�̱����wK��<c�h�MeNo$$�<�Zn��aߞ�F���IX�/�7կUTv�H��8gR�L�%�/��A������B�����p��pV3���ѓ�=��C�,�E�Hb�t�<i}p�`hUU!$��7�^K��.���_��1�s���%x�RG�!�v��R{��Lt��lϱ��������
ִZ�����ݻ�6�;b�Ǻץ�"���J�9d�F����v!+r1{�|�Q\��-���T�8 ~����:W�|W|tvY�S�>�/<x�#Ak`�,�K <`�H���&H�U/E�)�]	��O��WƦE��
��b��X�-�~�Z�-��Ձ	���
��/d�ބh��:]�UkW�jfi-ݞyZ�5�iNM{�f`��"���Nɇ�'h�K����X�"^O8�!m�ɟ���9����E�˯��8��o�����NX�)�sE�0�>l�]�!ʾO�F��Yi�w>c�X��ح�7\آ}�$�+ <���&'Ox��pa��o���fd9 �_'͊	sa�����g�MS��3Z|b`�@6u8Tu���M� ��GC��� '+������KW�]/�eڛ"��7͂��������guS��%��Ps��k�l��O��1�J�=7ҝ�&��J6�zo��UOI��y�����~F�o�P7rF8��bNG��b�������LŠD.�,+��q�+Z�p�B������B���񗇱�?�N0�"��mb7ЅbLju��?r�Jy�8�����V���LV����8'q�"K�Ű�/xx�?���KSV'�M���u�#��"*[��2���7˭���t^.&t����o�*{��a��WY��,��`XZ�|x���	���N��6����t1��g��^T��q/%8�J����Z�H������%�ץ#5]ܣ���gx<��f�i����>�J��ߊ�<�o��;��h/*pfB������m\�K}�ߨ��
���+����o�]�v�wqqӛMI5/&1�e�Z|�tg V�&��ē,s�{�(�{�w�tWg�$��t-o=Rh�:��_��}�|�[US�Q���qΐ��J���b�_ͧ)�Z=��!�/��&B�# zRV�lN#�Q��;���:�����Ɓޞ�m��~�$�+[Ԍ+@�{atF�L0P�X�4Y������/թ9|o(w=�@�}7��[�[��N��&�6P=���Ym��7�U�FH^n%%�G\����ϣ)�&��e�t���WP'�5�J/tP��D��s�>�v.�kp3s�TJF<�<���|���k;����OBo�*pkA�\�S��lXN��֍;��A&܄4D�T#ʗ���[ܴ�w���ή���5j���^�z�����'��kBΗ.7�$˓�O�򉄢>�t��5�=��x(s��xx�v�-�e�75�ģ�1D������0�?M`���,㕛�;���%�i�
T�֭��s�'t�C�y����b���j9�*�O$����QG9UTS8�}/q�b������~F�r*�s���u�5EМ�!h�_*0HSy#�:pnDf���aW{6��W�E�j��b�	�8X��/�,�K|9��݄�Dw�ӺO�5xyK+d]�L��F%Sm�b;LхI�?�ȃ�^@&u�5��/��oV��_��d��+\����T狆 ��8d�4p@.����GN����}���9�I�<�C35H��G4�
��t�,��̖�L�����0��ⱿnI�R��Y�!�e�)l�o���~��.9i�-�`��B��J��_x�O�3:d9 ���LpUN
�b��cC��9>�{�.��qAA�V�ܧب�Hj/"�҃��#�tG����9�%l�9��ZKZ>�6��Q�� ��x���{jX�I�E���r�@�s	��?���f���
G8�(h,�)��?�q��0;b��y=�Vg"/e��}T��Fw������S���|�"��v�%�"�r��jꢵ�cC9��zh~t�ݤcbM]|^�{~�c�Rڤa��{�U�vS���,`X���@�`�]i8���hN��M�	N��'XG��u���t��$�X�].��Đ�-֞�o�a�<-�a:v��?��v���q$y8�rN:�+8�K7}q�	�G�(Oq�)l0}�}׿��*�s=�lsD�[��������Ʈ'�OC�2�`H~v�@Τ�5lm}�6�(=/apS��A���|p�Ir�5n�3ԮT؈�<vi+�9ܠ��ԓ�*���A+�}���M��\�NN<?z��Tu����o�JZ[~�L��A��{��0#�_���8����%S�S���V���	��rP��}��ƽ��C�Ğ�BȞ������ѰGH8G����r�&���VC0�+w�r]���������̴H����Rq-&����4ugfW�y����_m��@�ac�]ºY����,/v�U&�o6B���?��p(ӈ��(���so|-_���8Z����N���;+����2�nO��a����3m�7���%��;(swX*����&��?�	ݬs�WIgmq\ ŠZE!}Lt+��%�U�ǘ��]�����Ԇ;�%�C�����h�P)?��,��`s��$9�[U�q�����i�-	���A�:� Q�9<�飉�	:���@��O4LFU�Hh&��t����Y@�9$��0:�.��/�������[�8�?Bf$�>�}���@�P�r�#�P })':�\D s��Qg��U�u=�Ϻ�� P�8`� �nC�&�j6RX/�t|���
��$��1=�eO���:U��W�{-@��� �c�w�P<i����e�c�o�����#f���;�3��r�	�;���ڏ/�ev���0����2�
��Hq�s�T���12V�G��P7���D3'[��,E�7�����tt�e���D<f<�HQ:�rS܏�e	Cc.�u:����������z�"�':_��~��׷�e�enXo>���7Q���J�(��v��v���\rG����>&���Z��],�Â���[�<%�W԰��sv���˳��t3�����N�&w�l�z�gN��phRp��z#��n���ohG�lRf���&���>=�-T�s�g6�%Fe��Vݸ�g�2��B� �DO;a>�n����$�q���)�b��%CI�� �#��HJy����>V��P,��9���?�{10נ"�����읙`�t_�5����5]�eE���a 9��)܎ڱ�{��׽�;��w�益��������(�J�s1i-��U�v���܄�;d�B8��Q��z��:a��!PD&ù�yҴ�_��u� $�U�1)���'D����D�Ǆ�����o��L0`�mE&	��Z~'L�v�[�܄`�f�`
������P��uK�\U Jދ`=T�@� [<aQ�s�锗�8��^1�KW�"���j?�<4�i#e�ǦZQ��K�%.�����`�ZD��&}����ŉ��ˣ��F7���v��B鉺��}k��w��b��+���[��G�I����B
�b�Z�^���;�4p��f��d͵�UԺ���2��5H��Y����)3���&z��▝��!YؙL X�vM�g�C)j�v���ݕ�V���r9��?�É}��<��m�ѻ�N���ʂ0#:��\]BeB�[��s�+�)a��>��[ˣ�t8�3-�ſؕo�2͘�3fkut�/d�r�_��CRN�4;9���B�\����63����3�s�9���T;L���N�"��� '�G��z.��<��R�Q���yֵ��Ҟ1��:[Jߘ�c�f�W���ck2��h�K�%#4K�Ʈ
��y"	9��՘�ѾT�q!���3���J��6���k����}�z��{U���d�f.���F�{�?>O���'��A�!�|9�?y��	��Z�e�W��R�p±>*��c̏ب�ui���k�1x��)\��C�r�Jْ��.f߶!�t^���lE?�[�r��l�Eר�H$Z�6�kT��}n�s
�
��I.J����H_��>�����"f�`7�hD��P�9<�y����U�j���ߖ�]ፌ?�ő�凕w�sZ��zj�Jֈ�l������� ~���I2�3�iՙ^�1r�?i�*P��4Gވ��V�n�֎4C@��%�im�����r�\T�]��E�v���#>y'<�?�������y�\���{�o+.�g���"���JeI������##�M;K�s�[�m� ���ߔ�Uٳ�gj<�q�t0"6K��~6�=��Nj;x�1Q�Y%l��	m-��X��g	�Soi9��j�	E	��{M�g"�

5�_ �1��j��N�UO9ɘY%L���Mhɇl�.��{�w��<
�(��N�Q,��{}�����ȋ�m
Z0���T�Iq�9��.ٹy�p�k�ɹ*`u�J�!76�e]?���6M�d�7�p��c5b�I�ԀX�RJ��`�(:f���2
S�j![�K�4�ldUX��AX�Ba.U��G����H�`=G��4)
���9?0)c��0��Z�u�8ޚ�7�_Mm�YB5�v���΢i��_O���v]���P���\�z�X�v����Aq1Np������F\�����N	�����<��KA���8���P�a�g7�S��x��5�Xھ��*2=>j�7$���U��%_<��G@�|�ѝ�\WJ��`%�Q�+�|��M庮d������f6�w_�V"N)=wl����wU}<�Bd���T����R�l#�5V��q�=�?�}��+G;�l)O
uWc4��4��Ռ|�2�J�4n0�T�����&ǿ�W"���yȭ\4�4��3�,�
p�-���V������r�tm_Bڅh'<63+��+���$*iN�Qb�c&Ԃ��8n�ݣ`�J���+����T�j�C��h�P.�uF[G��>�S!9 �i�F�4�8����葓�Q��
0OK���1$36Ok -�a�z�~e�$L�tR�aݯ�Q�ԫ� �d�U#�%��dv��^aIu�LnU�kG�~���u��	|�f��_͟�l������7���ʜ�U1l��-�}����9ٙw^�񰧀z�ݹ�s0���[ca�G�_��Xc�y�ꇚr�,fяdR4A���ET;�����(�H����Ȓi=�K��w�e��q�=�npg��~t(HC�~�/^������h�X@�U�Fy��Q���I�+s�����ހЈ��,LvY��-&)�T	����|]�P#����"� G�HǞ�F�/�����ƖP�VD~Pߴ	���u?�:ʹ�'&PZ�D�Á�MZ|5S�P��\��_@��.�P&�u:�?z|��c��������Ak�k��4�_��W��;,�!�,{��랗�V��?~<a|�v���`�QR�8��4���5�Mp�'1����`V�o��g�f]j���PN�4��K���o�>� ��v�wFc����5� ��O�j#p	��E9_@���rH��)��uoj;�ߘKE����FEf�[��ԲYg�khuh�],^U�J3��$d�'�4#OƎ���W]F�$'lNߌ�Yv5"u��m@]:g�@���'��V9��U4*e)�)f�71�sG�t�Qg<,���~՗�6��{���Eo�;t(_����j�ϻ�1A���ugڬ���՛NJR豠*�����6�z�7s�[��E'P�:���V�4� ���%�<#�#�0�J�oy/�>a 9��3n�o֓Κ���3��WB��L#B�ݷ�Y{M�U2j��\��-;�T�-Z	�e��ݣ�;�Jjf�S&6 _������ ����LG;"bu�� �:,��Ɍ����My����ʞ��)�T�vQ�}�*��G�R��L�,�xou��H��o��~��sƬ^��rs���z��%W�+�k����Ww~$ ���I=̂&�w�5)�,�?٘���&Y[3�Y�^��8U�^��-R�6T̞w�3�gnq��q�������8�R��y<_9�z��Y��V�G�G}��`�4�4��z��EL�p���S���A�u ?��W2��%���֥_�%�:P�S�[@E�hFHb���3bv}�(��{�7z��9/����RH*#����~�Oۦ!��+�\�a�C�$�ݪ�7+U�+���(��F�	�}@�ɴ)q��t�,���0��3�b�0�-dc���$�@Z�F��X�NX�ͱ��60�[�eV7~S�f~�ʹ�؎b4El�����A�*���#@�����Ɏ��˷�h��샆m�m���R U^�t��KJR�3�)y��:��ݯȽz)s���.V�wf��'�z�aO!e1p���a,�e�v�ԬI����d���5�z�к�Z�x>}.:¹������Wm�,@�sÑ	��%��A@,�q�`Νԩ��1����VT�WN�3�������������>&l�s�b�#���^�{4Hqȳ����=�}�I�r�1� M�聇N��^�j�8X�A���cA�N�2D����)��`tQj�h��WI��[�p���E���LwE�9��=Ә0�puƪ�����������.  �7M�{p{	����<xfK�����)T�P��y���	�C��@3��j[p�-�"[�^G{Zg��5Մ4�~�B>>,/�+�����x&��$A G�qܷB�־Ѓ�*�t���z��3�r��d��1V� p�����GܡIj(O�ۆ�T�+J�ӦP�@Ln���k�&c�p�ͦ9%[�c��N�".�Yr���G�s����"������L�����D�|2�^% �J�V P�M���J�M�X/�ǲy-�!�!馈Y8�:�u���@��]�"��ơ�s��K��"Q������k�3�%�^��ߣ�_M ���ᢊ!��7�I21��9�_Aq���$�s�l�$��Kg����V-�dZ�$lK�1"���$f�S$X`��/�.W�M��~r��>2�	���!-���Z��T��0�|o+x�\�I=(�،�ء,F���EU�|��8MK%��"Ex��`�g�\ �D_˄�}Oö��E"����Ú�f���f NuB�9��i
�4�}�@�ή��`�#��H��Ѿ9�]�~/e0Z��;��h�s:�F�����\�2"vz�Rh�@�=�q��(��eL��,O x��S�� \Z���������jZ;��%�˛KB��j�à$������"�t�ڦ^iu�1��m9�ȭ�a/�.�fS�"#L�<�ɮ$����|rQ%K�nG�n��6rm����Ƕ�L�\S�)(��CN2ʒ��2zP�a����{����?CЅ�.��s�a�����e�~�`��>�3<�m֜�\�D��rM��<���`I��q��Dc�? �|�������yN1�dz�[���`D�H��q�2�h����Z���qqTl�q ��S5-B�I�|������<�.��F�e�݂$,��GR����[^�O*n������?eN;�P~I��U�G�0�������K-���aP�ӏf�ӭ�ii���S���:P�O�-��9}�r�SY鼸�%� s�:��@T��Lk���,��No�-}D�$� �ۅӞ��O:�	[��T�y�/�=���q��|����1