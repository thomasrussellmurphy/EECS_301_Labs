��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\���V�fnvx��ÍG_;�ȅe�~�>���9�>��Y;�0GT��}��ExjXd	E�2�W S��5f�l�1�=7j�:Li�d>�$�����e��i�����+@� Ɖ�b����úR"N��xWd���̃-�jU����B"b����zg+���d��h�/Q9CC-����L�]�>�����l0��xj<*�"��	�I93in^����=Io'�X��T�A̸�~�x/���*��w��p�$��/�`�z�藹$dr�t����s�6����n�k�Ey�D�vm~)��B���{��I*�6!.!��������k���G�z����mB�����i�I]�ͻ��q`<\:��B�+��0�b���Q�0GA�fѫ��}��	����A�-<�ħ���;�����ܘ6�]�ӒU'�P+{�C�7vb�qT��T>���Ik�+O#�w��GP���ܡ�O�|M�ܝ=3��:�"�Ņ��n@
:Kߪ~mA~��
@����5	�����zQ��_r���`a�#���Cq&��;�c	�,g���O�$~��BB -ž`X�y�`f�>R����_�Uc�k�\��s�ƚ|:{7��[G�!{���F�E�f��D�������L�y��w�*�4]ÅD~
G7;�W�Uց S�3��d!��
�.l�Fx�Ҏ��Ze]��Ek�D�^�*#9{%�g�p	Me��I)�e �7/*- Ti�;4,�_0��Y���֊��qx=`�f�� [wռ
�r���6�M>�A�إT��h{�sNyƢ�b #J�vGm]l���ܘ���4��
X���y�è?���ɲ��]�{nGci�N��<-�(o�bg)�n�*�����f���Ә��i��`�V�B�r�Zz�TF�kR�c�Б=Е/ 6��|�C`��Z%V)�+�ٝ$|'L���
e8~D��ѿ���Cn�9�9��hKS��͍�2K?�]U܌��塚')`Aw`7^��Q����qī�D� ��pχ^P��8���t����?_�R{v�x����5x+�%��Ө?�P)O*S���As��hy�Q�q�}��D�X00�[Z����*U>��q"��0YJob�?�RF���D���='��D��?��] 6D�2�#	�7�Wd����Ҧ;��D4��AP�H ��xp�N�YFC[m%/���h��W������9Kv|L\�:�����{S�kϳ�ѓ6%%*G���V��c3s�qd�t�`�����N�%<���+0� )z*W=gk�n���_�DgS+�Xv�+���9E;��VFԪ��(�ʠ�Ԑ)��`� ld',�-��rYAPQ��[���v�:c�M�5-NG���NF�i�3�rok�p9S���ή��]8�x2�&��ŻUY�@�u�`���"eWN.�G��c��u�6�+S��@��T�˙{��G��.
-�}e�7Y�C���Y	G4�hx#z�0uq�0Q�9��s�Z>Yմq[Xe֨NSi#���E�wpί:�Ȫ3�_jv�w%�
5��s�c9�%S7͔ě4)42�ѻW��MT��� )N�j��hN y�q,)�'i�T��>�]N�	
��_��ʏ5E���wV���E�
t��=	3f�*eK�|��)��k�������EKl0��l�d'ɻ_�r�������F9�qI(�F��1���7��}%xT���N��H�F+N����!��K��~A��V\��y���t�5�����
�Y�~`��`�$�����TZ�1�vkь{~,�8�'�)�_9(̛��zf�dzt�E4[�x/Lw�P�ଽuA�۟��|����l��A��41t�c�H��G�O>�A�|�-=�:�1����^�Uf޿+Ü*^(�+�"+���%S�2m.ŶS�N���G�Ö-l���)ZO�uz����>����BJ���2{_��4�e��mS`,k�a"�=����}��U���)�%8��؟#����5��	���ߕ���������VpA¹@#l=?Q���`�i�r����9WC���14s�����{\׊����+�)5�Ỳ
C<�IXO�V���Z �3�D�~��2�l셎a+d�:�KF���CA���TrS�lC�*�-���A���
�o"���^��?�B��:�C㘾w�CC���eҗX�Qse$���x�^���Ҏ�m-���M+J��1�ۡ_V5X1��l��)AZ���xؿJ��s�-���d�؅n��8Ԋ7��=��@it��z� �lJ�:��K�A�M��K��2%栈�R��2��)O���N�>0�4$�i�Zl��Ds�Ox@Ƚ�i�iq���Z�Je���`in��E�7d}V��ټ�l�$�4J��va�t�zz��U�T6�L��P���)6��H&O�NJ�J�5�2%�>�ǮZ�7��ޒ��Sː]A+�r�
���ĉ?U��D��r������S ڪ���Hh�5�#C�����㕩2o���B�sY>�N2��J�����������M��y�GiGvٶ,[^�^?�:˥zj늾�y��Ff��q6ߐ��5�LV/l�������^w�w��A��&&>K�cîY;1�8���{M�
1Z^0oS�x��%1(�� e;�u�\���tw��b2pOn��F�6�=�H�S}ֺ(����땝�][��WGݶ�Ӛ��W��	=
�*e��s3�^���ĕh�����;�u�#��T�Ig�Wq;Mj�6򽰱d�'\{��,ֽ��96�
���B�����/2nw�]�U&|H���ժ����gT�*�l>Q;�z7��gxZ̪Y��X`=~I��J�Li�¿b���h24\6�h�rM��L���*���<����W���&�}�9RW=$��g���H�;x�X��g?$z�� ��,����2掌���C̞���|sUW�����6���a��T�d��i��d��s��U|�`w���X�-�Q�f�����`n)���$� �\&X��M���Wu�v��҈S��:�A���ƲI�ɻ�Ƈ�� ���.�gڜ@��D'��N%j��9���L�I	b��Y��&ĵ���ɛ�M�cg���N�m�"�{y���s]l�"�vr$����$$���X�K���a�#f8Z��y�~O�m�)����u�x��+�ݪ���Æ!����ؓ��4�f���_-�����z/��*��d�M�	��\w֖�2��ʫ���3�A����:|7 9�@&
���{��`��u`�8�'��
NZ�J�)� ���h��ũ֟^������Y��t�ND%�{"�&[� @�s#��͛��P�D�Ӈ55���~��Ђ�ap"tzmؽ�~��Ҏ5����H�l��r����8 ��Yw�+8̀R��aFr�0�Ԩ:�/���O�����̨���]{v|i����U���(��'*Y���� �~z97�S�YJ�SD8�&zv+7�� �ro��Y1�u�=�N(�f
?�Q�;�}"����	�_���Q�:^��+�[y��݇l��{�����7���H�L���X�z�jX������=
F��A��#�8�r��ڴ$.���Y���n�/k�(�Hq�"��j�}��.Kg���J�@!��_u�΁����F�(S��S���3r�?�s5b����σ�Π}��Wvđ$��P�ҥ��ĩ�
�B�r���i��Yw&�+E���hK|�\����gU�J����i W��Vܺ3G�9�K~��Sԑiȋ��!Ɋs�j׃0Պ��&���R�_�XK��&�zH~�ǖy� �"1�#)�%�1AVʒ�?�.�[Q�}�gr���M�����z;�����w|��@[��p�4n ���N����C��.;�0LX��:�Sh�4�wj��/��Ȭ���4 p �<�Ia�!K]Y���!h:f�c�R��Ku��ia���<I���_^ 4�P�QvZY��l�ۜ�����J�ʨq���2Geu.��L߅bd6q�P ր��b	ǅ{��F�����0�ѡ���R���-q��2^M��;����lm��XR����qY36��%ud�t��L��h	7�|ZT; E��4֥�Ѷ��̟��*�n�WZ�[��+񛋯���6��6"Ԙ������V���'�$����!��{c�PW#�Iiǝ	
y�B���"�i�S���������g}����_?B�%46n�<~� B�eV���L�>��NbPNl:v��ז8��NE6����l �Y�b8 J�T�κq���69	^�$O��k�V���	S�F�����c��s�����#�{��G_gK�&�tR#��� 	cT��&�x@"�����L\ ���&�h�ž1d�q�R��E�ѧ��!z�Fw^gfی�V�����C�-��}�Z�)��Y��[�3������SVLma��(Lf,g�1�<���6�㔀��$NC��#_�zY�h�B���::^.ם��{��d�y��r��na��o�=�v��Q�1�9@Qi#�����H��em
,-!*d<���.��	hF؁��wka����$��-_Q>�,�o0�3�'S
7�L�䇵8��� �x� ~Ng��.�J����5�[=�J�8;7�y�I���BOXqU���q�dL�����{��K���f|pdª���g���9�C�BO�J*�^� Η)D=��(ݽY9T\R+2�g���ҥ��9ϪXG5��Z`GJ����%Mi�
(]ﶰ���p�G-�l/.�Ν�֖�����3��="P
�=����beC�S'��;�9��#;�{��M�ג�P|�Az���YY3��7ζ�Œ����S���ZH���f�ٹe	���ٗ3��J4u���M������`P��0���\����|�t�U�U'e�8�����ZW��������&i��e���{�h��5�2������ԫ��t/2�J`��
�ڶ��^�n�YG����#�x����bv��V�0�?��ܦ4���@��C?Y��Y��Z�V�����u�J��\�n�|0Z-Nj�nG��hF��[l