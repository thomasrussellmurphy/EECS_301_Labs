��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>hs�*�U��Q���qh%ws�[d8����ݪV#P�.Bec�]���N��:�pیvB�&���C�pwg�헞�*f^�p��}�$��.������ub���X?���9{��x�
����!��!Hw�	�v������\�L02*���Bq�l��KrP��հ��y�I����p�x��~#�D�g(� A�O��iQ'�;�f�� >)����?s�%]oO��a\��f
�{���f/�<�V9���4!���h����B�o���/L9V�,���K �'NJׅ�X�.ՙP˰��_bȀ����X���d��PN���V!I�C����	*��H�(No2�]'&��<�8I�+��+�y?7������%����ZR��	�5F���ݾ̗�r?A����[�ؕi�i��be�y}��r��'6�t�;�!���=N�~z�]?��*���C��­��c����@I�Q�vOg��ۍ�q��BǶp��RῆUG�D�*��[�Tf���$��ys���У1�k�WP���d�f�Tֺ�nC͌�>�g2��������Isq��4�!��5����"%fT�r�����8��<ͺ�&�|u��R�j��{d��Q�I��/��f]O�dpE��7s�rAGŮN'������]��ɭ�F�ȑ�%/�,e��3�+LU*��{$Cp��7��r�R�h^���8�a�(��jș�S�#�����˿�d��l缥�dԱ��By��/��b�g@���2~���BS�j�hZ��=�ҡ�99+.��Z@�#o���wx���Q���:���#B����q��$H��|���N���7p�lX3ڽ8[���}�}���n�1����,���;�c�/��X��l�ZE�}e�����Gēa�~~�k��m�+o1!���!�8,D��S���aw���{~�;�
��u�.E[�/�˄��:7M<c��6�70WX������6�4[����iC�3{
��5--��`86z���X��B����p&�K��6t��"�����2�����]�O�k�,�ɬb�]���/�|f?v#růh]!�!!��|[(K�e*u=F�Ꮥ d�>@�R���~t���$C���b5�v��ʝ�������eoih�ѥ��6�ˋ������_�r��!�k�U���8W"]u6H6 �*�6�Ĝ|���C��mw���c������(�\FY�PI꼯VMh(����V�<N�Rԏu=;��ǴhJ��9��3l������m�i��e7&�h�!�~��G�ӂ�For���"#�� p>��]�o_�U�"��X��n1�Uq mҹ�i}��S*.Ŏࠟ����bI�"�ҿF䎈�-?;j��,�/;���17���&�"���ּ��QT�E�Xe��H��pǨ��c��oc4����*$S�O��04�t-�P�k�gȬk:�Q�p~k%ۡ��m�r�����=��8�ٌx`�%�_Ao@h$}t�;��桁1��P���^>��C�<R�s(G�_��'Zp�Ks`lK��=U�����
A�0Xk?B'%�A>�Nz���R�
@	�1�����[A]�z�^��v�/��Ī�ԧ�����?�
����@��	���9�vWH8�}��!�8oΓ�3�%b3�JY�Q9��*(o9g&�o�l��ݲ;|�\��E�3�E�y�"Zn,�Ե������y�[o(^&�Qͫ��S4R\�,u��m�glH�9�g�F�0 �X?�(On4�8�*רA#�ҳE[�P�ʰ	�:��B��n\|ڍu�ηu\�%���X�,��v*����Y�C^d��8^�T�Z�����iⷝ`�t ��G~ϯH��OE�h�RV��i���T1��,�}G����"!��d_�� J�Z�U�U��Cj�>.���3�V��� ���_�-<�@Uc��I���`l4L
ca��}���#������	�\K,�uJM16���Ca)=�Ѽ��k��M�Lg�>$�Cʱ��߫��ܞ
jx�~<�I'i�ɱ�'�C_����D�Ly)����I5��"�ώ�p�GP����U��T�1�z��ɫ!�V`������KȊ����ad��T?!>v[�XTZb��Jx�y�N��R����u����!I�������5��!�J�z��lo63�R�]�HU��n�o����,Q���Χ�5��7ʑ����y>�3e�����"�����j���f�doC[�A5z�6�=�I�+9֨[z�W�ӕ]�J�����=kW{����א��a��f��E�u��н���@�w�%띰 �O�d5�zh�rKFQ��b'�q�:��Y&@=iu1�3�m�G�G��ՕF3��n��� 
I�UfC�_��@���m�_+�jmN�=!�S����38���$�EC:��.ёT�C�����2��"��>,x��a�\W�K3HI^�eB\̝#I-�"3���wa6��z^��c]�W��\�%�a�.�&ܗp-P���>�C�t2A 2FT��� ��߾�w^�u�F$-�D�}׹C� d�hg�+�Q���I�ǲ��Ý�`]G)��ND��Y��1J��b�u�2�D����(N�����K��������`��#:<Qn*נW�b�n��X�e��gV�g��O��5 d����<��u��(\L��x��}gܭ�/�Tl�r|Xs��V>�� �N�*[�-�J���aw �[UD;M�?��%���~�Ă����m0`�z�>&��ш�8��̍�"\��fזZ9C�~釈%���+���1t���䗣T�T~���8����j\	�_�r��(��(\9��|����+�5�"%��s�Y4h���5��g���c��ڧw�LT&�}�`�=�J?Yy��<	5�Z[��NU=�֟	�QS�o5�����
3�~Z�&��G��4��e�⅋��	b������n�[|��6g��!�=�	�"��wR�~�r�6�pIQ��>��	��^r�DF<#T
�pYJ�vt�y�2�'���H#�)�r���1=�Ls֞*V>�r�Ҧc,�9�em�*A�l��Ѥ�<GB�j28�\�zN�1�ǗT�4Z���Ǳ.Ø����T���L9�G���_Pb�S�c:uǇ���_I���	AN2� �A2ԍ��+�v� ���և�8�ޞw\�R�O����<�O�9rAf޴�}�^Y�|�\O�xo���v�|��x]vKnIY'2*��'׶�a;[eK
f��_��˓�4�D���/�4��*�e_A`����3e����xHKt�Փ����	��&��%-�s���s��=V�n,��}���{38��	+��6}�+>�AKe����s�� z�5f֤cѴh_��YC��.J&����ߛd��[YgU>C�oǭg�g� �j�J5�G���Ÿ��>	����E�-�%�v�8q��Qm��G��9��YP��4�n Cn����/�π��㼁�O��,�0 �\�g�4�,�>SNԞ�$ۼ'�%����h�4����j�[V�m�#�v�-)o���q��z~#���'8[���ag����%ȼ��W�%q��'����?�?
�wN�0`��݈�^"0<�P�'9�y7���y��:�$�`�kV�n���Ѹ�~;��;��û�E��!I 
�\�!�����=:�3��r��Ƨ*��8���X��J������L����Afܞ�`�
�%�S�WQGk8'1;�\b5�s�A�S�$��ºp�c���3(�(yLہ:�����'-�X�6_� a+���EZ��]����yAo<)pa��Iދ�A��=���5�U��CO���;�F4��ܷt0��j�r��퉹�!��@���������a�0����0�ь��4-!iwq=�Bx �U�v5�z�_��![ ��{O�!<�����%8{��q˓�k;}�|�vB�ǳ'I�!C_}ݨ+Qm��1Vs>&�ay�&��ڏ�U2:#�9� ̝����'stirI�[�È�!�6���l��Vt"��M���v����>�� �g��U;xb&�Y\��a���Ii]�{�\�v��"�]P!J7_�n��)����)�Hu�^>���0�I82ZB����Z�X���4�.8�f8_�Y3s3���Λi�|I3͈
�Z|jQ9d|a{�ؘćj�Q����4�A0��'*�Cn�%�� ���4��9<U�삊�§?%F�{�DA�x�q�{�x'Fb�u蕨�E�9CvĤ����:I�}��p��V�%����N��ڼ���_��&AsԐ߭~d�U��C�/mè����4��i���q����7{[�Oj�Gg �����h U�7 B��8�bk~k� ���]3�n[���@��4/�0�Њ�4�8�oe�C�2<�a;;PL֘�`����Y��|rᣋ��H�����$-]3G:�Q�c���RwKN$%�JwG��SFw�x]���gGVy�d�k[��Q���q�iG��I��g���|t>��60G�)�$�j��m��Q=\��-����7w���q ����5O�~j��z�n�f��֏%y�;B����IO��>�Ӵ�"���H�'#3�jj�!v�TSy�O!�^y��)�Txv��_�J^�/Z��{��啾d�u~�x���R�|�{��~yE՟�w=IL1����/��Pf�`�OT���Xj�/IM����Qk���V5���������7�'��|��U>|�")���ۘLX���I��+�E���mpl�:X	17�tDTq+�;M��XŞ��IN��^R��A������7�����t�*i����ڭ�О����1 �
��kŐhi�����_N�F^��XӾ?���sS~g��D�f�UN�đ����s
�tr~e��5`���{2A�}H�M��L��if�jN(tϖ��0�*H:�l%^��KS8�� [�ʺP`bg����[;���&�f����ۛG!-����9<uW�� %$���mS�y��E���[�	1
|��,w���ǦMp9��������ڜ�o69b�_m{�y���&�r�h�_{����*�8���$�`Z��\�FA�����|�N��nM��5g��7��	E9Z�u�4�(	`�y�E�D:��^#�(�w�/9�|b\�X�'ͯ�����ƯU+�\�����>"?
9���(D0}�� <��yB��'j�ݻ��X���Q��Ǘ.Y�^�\����S}8p�)����*yl&��v��U2��36/Q�p�f��$�a��i�Rp��ƣ��Wz�fk���z�z4]�~q�Jz�2�����Z
 ��rR-l [�9u���$Rsě?U��ح��BoiW7�B��=����%KI%c�h b� =![�Ú_ʔ4��qR�X\�����sa#^��;KA���j�(�f�E2�02`範RN�� ~�+&����`<dQ�-Y���7;�Ҹ;氷rP�st���Ay�V��]��������H���੤lzQ�U�J��M�=�ԣ6q���BGKQ����W������~3�%�'�B��q�'����[�h�߂���G9 8)ɹțP�q�k�	�/YQD/u�U�D����A��tȅ<7;�G��!�ۓ�&��K�6b�!��˹v�������L��Č��i��#P&-��YU����nQ�D��=OF'�2�)�W1t�u���	�8�_�j�l$�eI!�_�nS�m;�$��S�X�{6>�
��Y:���*d�ѽ{�����ۂ<,�[ϻ�6Х�#.�V���	�%%U7j	>��Jc��@�#�R��(0Mbx?7*2��]�$�~�?�#�=��N�v�M����/� ��T!�Y�.2�w��)*�[(����!3���������Bth��")G�>�G@�	���},�x��4��D&\�����dƤv
���� �_�Q?�-�7�mx�;iӘQ��{5�qY�
�w�:��������lw8	 �l8��vb�ތ}�m}��y%��߾�	�ק�R"?�@q]9.��6����TW�)��|�iF��	Q�w�H
]��jx�Ғf{��R���i����ӰQ��v~���=6W}\Ǩ?]Ao��1�r ��%���$��-u�_rh�ae�4`�ԤM�V	�b��p�� �{Hor��:��3J{�bF���_��D���V�vF-T���A���p}���d����1�T��Q0���nKff'>o��~����d��� 9���R�7�c�0��3��,퇑�t���� {�ѐ��z5}�6�e���e�㽿�|�k*�z�q�C)I2�R+�������vM�j��X t�F��h�8Q,7f�J�զ�*9wO"[)�� 80�{��B=+�W�2-�w}�� ���V�3�j�s3���i�	|��k����5�*�'��Ʌ�,���{!V���D G�"\�L!`H�g�T_�l�g�Zev!�&�vIQ%�\@1p�܇=��7�E]�T25w���wE��M�����4��1���Z��ź�@%�1B��&W���Ϳ�G���]+�J8�t�9,�j1�O?%��?�Ŭ+���]�����}�"�k����˹�i�>�Vuu��ȃ��%r���˛K���v�� ��nf7V΁ر���ifC\}�C�������yl1��bX�x��1���*�O�L�MQ�
4��~<���N􎊢Kr�!�D�E>�'��{k�����JnBR�	wE����Kǿ��	sy�qC����2�� �#)�K�(��D�cΆ�rj��^k!��v\�R 3�=���鏯K���-���Ɨ�,\��.7 ^�~�$���J��2���eT]?-4�,ַx�e��X��_���c��؂����& C�Ƚ0f6<���s��,zO��$��z�-&�Q{3��AŠ�o�;�[{�ĭ��?�@��hx�>6SZ��%��:) 9`ZO����Iя?�K��]�`xF�i3%4jۆ�>'��4%2��;d�����Vd�q��=xs�]��&M�i}�����+� �&�U&!)�8N�¶b����dP2U��������}�g�y�&�U���mw�"T���x�!t�H������l��q��A���џeDF�O��@g	_������Lb�
}�H�8f��Z����(̏;���<0�2�R-��ć~.�F�[�t�l�BK���ސ ��&Y�}��1��O�񣏩��vF��
�21��e��7*��X6q�e��pG��s��6�ưE,�� �(P�(M��I�tC:�ar&T&HI�7��*���&ڛ5l�'+R���Ϳ�=��<�}��k�	qG���>S$6��ɧ�p}�&pf�5k����i��Qͼ&�N��>�5��QRx�I=]bi�S�Z}?_mї'�I^u.qP��*��J�$�{�t%�a^���:؂h1B��s����2��7�)�I�`��-��Z���ù	�ϛ�1���(�ꙟ��n�ͳ]�7il<����!/�Μ��e$� �B���Sڼ2�aSL�r����k셐��I�'��G]���g?l.PRr�t%4j�J���.�����g�U��x�T�����P*XYA�~�ue��p�{�j��V�T�š�F�`���=k���