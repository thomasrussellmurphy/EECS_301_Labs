��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\���V�fnvx��ÍG_;�ȅe�~�>���9�>��Y;�0G+��{�d"��sJ���z�JH�t��	c�jI$����߀�':�����}��	�jC˕O)�F������	:+��E�<�Q�8���Ǐ(���dT<�p�as���]=6��yDl�`Y6��+�,(Q�b�B�v5��f��q,�ѩ6S1��o��[���+��>j"�[ Qd���y��a;� �7�Qj`r	P��Y�N�5E���Rr�Ie��B��Κ���L�%{���'&9�I�0��{bH�>�ʎ��`�,��97�h=�L�}�t����Q�*�K/i�TBG ��
��� ��@ҋ�97+0�C~��tn/%���~8�O]�Bͦv��Q��9�Q�;lʵ�:��ڙσ�� c�zgR[�uQ��w�^����ђ���n4�j�����A췤�&_�����S@b̓�kg��WIۃ�<������hu�p�hRO�d�"|<Nmf��_%A���xa���WF=��\H�Tm!�A�l51,QǺ�,m�_�jpG�6�hj��C��E:�<��BVo�Xp#@%�v�3�n�0�V��$T������kN�!�fSLqgUZ�l`�͋:ng�va��Z)�t [R��b�-�|��c�Л�h��zEQ���u��Y��QG�w��U7�k3��V�EX;a UB���Qt��s��k��:;sf޽�u��Z�Xhܢ-�v7Ssg���J��:�y,�ǽLz?�NR<�EA�x�Τ��g,���CF��u�c
v1�-���k��I�^�>�?0dި���9�.� B� ��f�xA�������=��`q!�x��ɞE;�-�(~ XB�+Z��S��P�MFvL�"���וֹ�	�^	,x���u� ��r���t�r����a<h�����n��M�X1!m	(�4�K�-�U�lg����vw���j,���fF@���� ���ؒr�G,��4}�*��ݨ��\�ʋF#=����B�� �X[�s\8�V(��������̀.Yנ�Ci�\�
F��!M�ة,0����p_�YՖ(d�7|�	�¸�hV��H}%X׷T�c�\���H�Z��F}�	�oOn���M�(p����,d��B�Τ6:�|��n�~�i^|΢$��.�Qjz�R>3[r�r�!2�ݕ�p�h
�����C�h�<����Y/j8��ub6���$�D����}��D��4?�tn��H%��c�����8�}�3�f���ܭ5JTVP.�<I#B����3.��,��|��e�,��x:��B�3j��Q4�6��U��ʏ���fI������)�� �3��	 ��T����s>~r&v��3��X��^��u3����1d�)�a�>�8�*k�o������C4�eV�8T��6(f"r������=�ʶ���Tp��5�2?��4���NJA����+�ێͤ�=��G��Y��I&�I�+�Idk�ɥ/oOG���/�in+a�V�PRkx���ٍ����<M�K�j?u�n�sġ�����+_�~T��+�7�`
Musn3��i�nQ�ϊb}.��dJ|ޞ�w�P7$�]R��-��lVm'աG}w7��"(��g!ˆO�k}��X<R�?W��~� [,W[S�cG���H�%b�QԌ��Jb|&��Q��J*@U�h��4G���HHZ�C a��pkn2��j����Oet��O�gdoB��"#}�",A������qi�Gc!�)���JkM�Q3���ѣٻ:��I=0<>�(�̛��朇��s�������Y�%"�dJN݄���G��ز4�7�5�D��O���6h9f����,�+l#�ty�f6lԦm	�"* Q��{'��F�'AU�2����zs�f����̪b4�[�*�)�H�̂(t��d