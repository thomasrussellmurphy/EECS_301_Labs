��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��S>q��}���C_[��\�O?&�;�/o�X�'���V��Q<&ma�>���ի\AQ��R�1��PY�8v�g-��]��KZ�CZ��D$_��خ�6kFa���f�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�i��a
Α1S%� �uj?�L�3��TLei-3^5]E�$���,�;�^���Y����.(��A����ص^���G3Z�����q��8��.��9�|���fK<s��2KzW7$:�'�u���dF�8(��-����yVU)s�˭G��2b׌m>JF7\ �ݵ?*��`(�0��8/y��*���@svĤH0��B>���'>�uHu��m���U���Nf�7�bz4V�q�؉�'
�+����
����%X��܂#^Y?@�gXY����B$e���Q�;�+�|u���Mt�x�02t-�l{ܠS���9�atV�w��t�Mj���Yb]�;OƉL	랿6U[׵��F�ݭz��w%�N^����i��b��+��i��m꠿�ݍ>�΂'�����jGOߎ؄{����u�c�s�q��hv������$��!}��G� ���J;��avd�Gq!�P��!�CJǹk��pU7����eku�W�'�wD(�G���{�O�9Jт
�W�*����$���n�Ntj��'�C!5)�-a=��@7<�y0`Yʶk"�a|�b�)�����gp��j~h�:���F �YJ4ޕ���v�#J�	hE9�V�hg��l��n}]���D)�у�D<��P����Ō�1>�[v\������� v/W����.C"6��Va���ײ�;X}D�����BU�d����m���������@:3^��iJw#Շ�C\8% e����C��C �>�ؠF�<��~]9�s��/':9Bb]�6��u�.�x�SeD	k&dT�t��B��[�EJr��{Ek!/%h��e���i��R�aH�Kĵ�HA2�趄ޟw�1ћq���҆�eJ,�Pũs'�.�� ե>(�nn�����*l��Y�1EP�����Y���P0Զ�!���>��p���y*�6r��$�ά-��]�4�1��<A��	�ȕ��R�BZ��.������Y�g;�H��!��ְsƗ�炦L�Mɗw�px�L�D&�:�u����x�W�?v'#��p����e��s��1����+n�N]_㬶�pG�F��Ϡ�F^}D��R�D��uP,�?p!�"+_��c�K��rES|�l�N��aLl��^�-�n�%0�@m�)}:�#���p<��;r��uU������lFj��;<�n*����!�(��������d��X�����
"����5��d��ו|n�#2�fe��"14e}zz1���8����F���.QK�z�i��l�����ZB��E����a��Qy��˺�h�'�N|3i^?�.����	�~)�u`�?�yz'k!�>��Gp��]r��0� ����!z;N}�8V��S/���1��R�PTB����� MS���Z��'�:���3�"E4%��?�E���f�9��Z�x��Q�P������<�zX^��H8#vE��HyWU�/�A�?z������V.��R]o�"�_Dۨ3�&��#*3�~�K[�L��D�|��!�)sW�f�r�����;�:֛Uұ�do���m�/���x|��eK#����$A1!!����paJ���ӡ�)!��b�_IqpDh�"������j��"lE�f��
�]�w�����j�ݛr^�H������QW��佧!��Bl���R��4��ZR��D(��@�=�RV�٦@���fM��v�ǆ�G�hP�Ս�I�#�,�����������9��VJ�^��)ٚL�WTr��>X��	1.�ilں�B�LZ�O�,;*E�s����0�VJ��u,�mOt�H����D�W�ҋ�Jϑw>͉'���:��J�'
/��G&�"�������\ ��w�F�z��vD��-$�F5I��/����U���IuH#|�q��ьa_�Fd�^���CC
��UƜL�n1�{>�&��;b͢�HC!�:���|��$X���9�h�z��MS�{=��j�`B!���[�I�w�MI"��9�}/G�4�1�n�i�*�5gl��h��0Y#]$	�����e2��:�홏q���G������{��!B�ҪVp �X��'y���mQ�L苑�nU�e������䥶A%,�pNm2�~�O�qT6;�������RTٺ�+�v��b�7���;$�y4<�y�mam/^h��,v+�0IkI/Չ�=_�b�15��t��	����u��Y�M���"��B�j�	*S��ŗҧ�UE��"��������>�w&�l�B- 7)-|�o�5]@p㹼i���w���;t^�p(H�	�g�W��Ch�չ�6qu�T<f��4���k`f�st�ۯQ)���v��.�SU[<YS�K��JHi�E:
�	�`=÷�Y�;�6s�FgB�����T��D�z�,!3"l�y�}�2�w_��c#{��x�}�����wGȋ?��"��ӷ�8~Fm�+g����۱]�|Og�k�^�䅃�j�x&7e�*w��{��lV�J�^�M@N�6�;��cG,�(�K�y�Uf%
y���J���Q�l�N���\ٞ����J�y����ɨ��Dt����A?��~s`y�I���*�z��~@qc��7�����4/Vh�U�9]�bV�#BOӮg-k׷�_U&�m������%�V�����3.8�g�"J9�s|�'y5�[�C�ֺ�+�wm������2� �������oK�s��+��[��X�C�tlJ8�ł��e'5�@�3~ŵ0kT]�A�΃:�@M�f�p�+^���T����q&vG1��~B���em�9R���PsD�l$#L+�=�@'7�Y#�������d�H�jhes|�M�����ĲJǷ����z�r��x�=$2i
����`�u�׾�'C����xǠ��B�����l��ﭗ�3�p�в�l��?�U��� Q]3L���a!K2���\����rc�J��5�3xR�M�+����h�N^�����:?""4�=+P W%�ct�^�ѽ>�vAY�_T�i�3e�~��0P����S��⋳��D����J��z8*V/b��������5�F��"��j���>"�L��Ѳ�ɐ���]�pݙglOJ�4���K�.K�i�j���A�?u�Y��C��O��P���n�[b��1G1��;��Ã�TL�f�W"%1e5�i����-����t��f?��e'7���� ����}�v������j����x�U3�����a�Ҳ�_Ȕ�
�gؿ*S��P��əI���Z�o�Z��?9I�D��d�fu����jp_0��͚fn/\.NV���-ql��͓ۈQ�炩���}ypu�՚q)��L�ek��t�V�k��u@f��xYIM�e��N\64
[C\�C��H܍�;$V��Bj�&@��B�s5�2���a�����;���@���i��}T�,f���Z����2,��7��f�����j���W5�ę��~�n}K�|�+Y	h1jތILKPn\?��lV(Q�N�^"�ѪYM��ŵ�`����V�馃#��wI����AHD�F}0�@e6��h�����������u��P..Nf7�i��~,*���@�اj=�9 �M�jT�T|���A�͇ސ��E�����-j�c�:,�4C�g8K#{VTe�v��/�`� ��N[��dAM&�0���z���oC��� ��}�s3�<(v�>�Z�F����04�M�~����2��!��:�����#s��-##'�"�C��ѻ�GMyFK�I�>�D�fnI��P�b;U���*̀��ԋl3
pg���70�K�[����rٵm4[��Fb�������l�;�fb����d�w�ꯦ��;$�N4Z��2m�h�{�5�?9���J��/Ď��z7�1���
`�&�}�Y�r�� ��T�
�m�W;��7��Jh�W�vn�x�
�w,M��R��Dc��#���D��
��]�Ed�9���ҋ#�ѕZ�U�Y�p�t�����!8��2���Dn_�}\x��yo�Kz�2_4�����0������.�q��o�*�T2����== �ǮٵGPY�s�J>9�v?�� Ӛ�-�BUp�r_XJ�����0$֣��W?A��XӀ-�C�^�AҷP1�3"��B{z*K�?{vK�`����t����	���i���'*_��ĕL!߽��`�hs$'_xJq�DЂf�Ép�MŪV��,�Qs�t7�z�P�!��a���^��#�!�@7U��o ��F;�h�tt�\M�.;�p���Q�M��c~��d����pv�;]��Q���L����Ykh� -����{MI���$Mc�6S�i�̦ ��� ���#7�������"�2c���|�rul�]%?�?_M0]͊o{07[����w|�����̚�D��t
�/�Ӣ�����r��K�A��&��:����̣%��7����y����O`d�D�'��:�
f����㯉�$_�K�t�Q�'<@{����.�Ň�ʜe>}n1�"�dS.x�kd�0v���~0�x$�k��W���ZƄ�����|Xk>RNT�Z.�蓚�PL�j�h��0��v��ĝZM[(�_o���Z���k ��%�����q�Kրe�d`'ŗ
"���N��l���1I��4lˈzTf�u�-B��$rf+c��(@�M�g6��ɜ�q	��b ]���f$�h���a��4Gt�[j�V5	�T��DtGts� N}��@�J�*�ZK�����f{�`�2�^�:QG�>@eIM�������;����K�G�1��AUM�Rq����b�FBK������y�Q�H�M5uB����(Af�?���ۚf�d�e $��s�`^SXs��Qݨ�_t��oK�C�k�f�ӱ��Ӯ�^�[^�@a�r��ڐM-]�o��OFzCe��S���^��t,0eyĐQ8װ9��R����ږ�ޜ�M�%��/�͉͑�׎δN�lHC�����zer�������,׶Q��u`^�AF�O��,9�����-�����6����UZ��-�������,׫�!=����~���Cp��E�E�t�8��zr������$�W�=_/Qb��1@�r�("�`����9��?a�pA�^�Ӄ�^�?("��']ñ6
前}�YT@�㛩aR(��1�&���l���F���%�,UMH����8�0�I�C��;�:�O`�@�0Lh����.���l-dئ�e����;��� *'	9B�*鼍e?�Z��*v�?�z;q�k�H��\aL�|�OH�H�Oy�Ƚ�1���u)� ���͇��gc�ԏ���(�S����B?���~�"�2 }WG�B:p��D��XG��@O#�����IL�����j����n^�������'I �.���??� U�&��	��h��#�����܉���=��Q�%;�E:z�����%��&���#y���.z��/�H�3�k~ a!�ڗK�
l��
i�փ�c���uiZ5Z�J��d8�Cz?ے�av��A�Y�!B,�:]>�n:�GXq�����yiS��=��h��E-0�^�ف�D.��5�gQ�&)�����9)2b�X��Z�ڬ�U�o���F�0�'�U�ƂR<$a�V���OQ:���C�8(�n�F�KW����ŋ_禃�:r�Wo���2\z4[�[*���A���}^�]�� G��
�
�y!�?y��W]���K�bt|]�Y����a�2]�����<���Iq-��A�oaC��f�"��یaF)^��7A�E��Υ�q�D�@���g7�_C�qH�۴k�v9\X��9���	$�����=����0�\�����&=���4� dC!�:�����L`,�p� �L�5f� ?���4�8�����3��q�:�F�z���u�PK�QG[0�F4H�nz#�,:vp5'�F�n�Ñ�v���g�
&��I�U�*����1�I�m�Km�o4��w��b�P0c��F_=�ݗ���Z�D�,�+�/|)^Ґ#/,���pz�[�X!��e�z��^�}�q}�L5�-�1O�X"OÝt�SL�(U�y�%<`\Va_q�XA����c�,��U���)�c,��1]/"[9�|�� ���z�lSJ�Ox$,�Q}u��v�g�G�[;�hc��1�}��oP�fU:�#�%qd�L��MN9�xh6K#��h݃|��!v�?�{I�5�=�)]�@����G�����0�S�}�$)I��v�_����n#6���K�\�V#w��f}M���7E���|�^g?�{����R�'�s_��fb}H���L,G��v����h	B�-{8&����J'<T��K2�_L)�"0Qc��:]b���v���&a�Gt0������`W��r�.+p��}��	B6|�Noӻ� �qIe}���Ȗ�K���.7���8�����m�I^<Q����M��IMȈy�ܻgr`�47�h�C��Z'����|ӆ����'��h9���F��_s�n��GF��3�s]���3u�އ
��/P�Z���M�9���������n9u4t�]�/����%��p:��`� ��vv����K�^�� �N��h]	����� ���QB�J^���y��'s\����<��W��D����+�J��v�y�PA�����n;���'O���>Z�:Eᚽ�6���@���V�Tk��!l�_����;���³�=A�,��q��-�� F�[�kJ�gflH�3�"���_����%�9j���V�9���|7������&�/R�9���>ɀ�V,�z* ���%�T��HMa�lV����-+��a���ec]�C���S�L=�_x��Nj�o�֚r{�m��'� �Mr%�`��o���1��jT��e/��5�Ь`X�Y�:T�
s�����Lp�n�f�%MpѢh,����y$��p�Y? w��4/K@*
ThV�*���2�D��ֿ[�Ez��|+�j��w�Ka��x��� ��\�����h�V��S�M=��W�ط� H��C�����	�n����=L�h�L�/�<�V����F��س/�gwv�[˜i��o}6N��︬ڵZ���1�6��pĳȤ�������m�W�0X�ݮ�:�7 ���˗##J����i;E�*tt$k�5Xx� �c����ycsz*�6�"�|F����� ���b�w�-r�@�K��.�_4��a1�����T���RY��W�?�����V1�w�_m=5����R������K���b�VHܾ^6n%����w-�s��»S�P���y��c��ԭ��MH��;�hmw�ϝ�e���@����V�,\�60^5_p��ЊJ�P���WL.ף�����-��W+��˕~��5��n��}��u�O�o���		iQ�r�%�ph�.��3ժ(S���?i�[�<�>�r;坞E�X�g��*!zK���-������f^��l��q��O�J��bc����OC2_c�Hdh<� z�lE0x< p�(��D��R"� 6���$��d�1hwX�^Ο�.A5���J3ﴵ+��;~��Nwg�$���KM�ߡk5M5�
�s̻�BI�n=�E�@�flz��ǹ�4˜��y���n}8o�L\���D�"�4��Vy��lI#�^���EÄ�;�D�N�_�K��B��d���Df�t	$��Zz!xH:�}�+w_����&�+�w���9N�{3@�)
T�V���<�}S�Z�=k��f~")�{�s��BP~>io�R���8�>�l��h�
 ��Mt��_@��^gգ;�g��B'R%fqo�η��+Ŏ-u�<G����{�8)v�y�����Q�[�zGN�z�7����\+�!�=d�� �̼�pV�-�&��LR�
 c����d��D̊W��/ 3b[0jMΘÖDfs������|�C0�S`'��S����c*E�oA��j��1$�.*XsI�J��N9�I�m��d��b�|���_�?�t��|�����C�e�0t��Oo��U��b=�2p�������`�/����i@ŋU����e8L��'5��|�_7 ��Sg�I��^i�i�nl�,P<�P:�{$l��в�a��1I�(]��E�.�Ԟ���E4GN?l{�A�F����	��	�J������RRE=��2hD@GL�B�9/��A`Sq@��h/N>Yy�b�Q�P���ݱ�>�V
�D,��?��6�Z�SڎI��öx)C!�;�B�>	U2�Vu�R	�N��b� J�/W��Y���wc�m�����!u=�:�ą���'Y�2ݜӠ�n
�X1�Xj-:�6���������4HeX������;�9�I�;-P)5� �{�jV���&ڋ~:&��5b�nt�[h���"�k�����j����`[2|��恥$��ǯr�Ce�j���@�0����n�	��`'�(�J)���@;^y�@��9u��gD���J�x��0	�QW"�su��d�tbb<�M���T�aQ�IfA��ju�p Pb�*^D7���>����V9]5{�S'-ğ��FP[�n�#{�PF?Uߝ�xթ�+��/6�~��)r٩�x��{v��d�c�Lx|	�_ݽZ�>cT��|X���:���]�_j��V��ގk�ST�����
�ȄZ��&@��k2�&@'9�gPb�,e�-"n#�G�; ןELQ�8c튿���h��=>ќ�56]�2r#�nL��[��\}���[]���f�"��j]eؚj��㣤�#�ɿg�jb�t_�&��ɽIz���r(�(�]yK*�o��u���ɿC�&`C�����
��]$-y����tJf�U���%�����!V���S�D��!�+�)5@1ۣfdc��A})0-��.=ԵU|�0Bh-������64]dƯ���
�5ޑ4��s��Q�澯gl�sLA�)Y��B���p�B�ie�\C� ����6>g����K���}��1v�&b��8��Я�k�� �#�x@�.��Ű��8��<�A�_G�Eи����No��	p�ٗ����a� �`�[v��`
9
+����*sZ�̺�ge0eu�5m�T�� ��m��\�4��*'�G,�J�^�f��� ���6�X�P��}�_�6�������K��iH�,m\ò_����a n�w>����?�]��1���+#J	Y�����7GZ��q[�-�-��u(�fN���L��_���"ў�P�!$��^4R-����fwײf��,�.�"#��?4���
+��%�s'�Vq[���R�:�'�f	�A��Bz=q�/�1�$^r��-�vM��
��"�p�"�va]��ݻ{F�H�O9$��g�����
�mGZ���O��6�_/'�e��.!�H�+`@�	���^vhn��#���z-}L��o>�����P�#��]�v�#��>b8��*��WO�H���FS���%��H�� s�W:���-�aݐo����.�etٹ"���Г��ޢ��X����@u@?)�^�
�Sfҵi�nS�;���Ϝ���*l"wz��8y:�%��a�dE��v�#���|̾���9��WΊv������c�~�׬����T�b�P��R'�AUr˖��}�X+���[+�N×��������"���VZ���n�*��t0,�]���B��KN4��y�w��=9�~�٢�"�PS�)���G��-��O�8�F�&p9�1�(�@
ǂ2���L���-qcW�s���������TP���YG2�ɯ��z�F�S��K9�0�^�3�<@l��A����B:�R+H+I�*"�$a����𧈙�s���|�z"ݥ�ܑ��E����Vb�m$�'`��(z�f�J��"B؍���ly��[6�ٍ�n���фC����5��vq@
	�`��L?H=D�$ݖ��Ks����f;-� �Hc������U�х��;;q\9�4s�R��_v8a?oJS���C~�1�iE^����B,�x�@�6rBS���s�a����9�5�gS"��	6�Z�>Qg�$�(=^t&�ZS�Z4�b(��sB�ّB���w������iJA���)+]� �3_�_i�a��Q��].t^ th�_�Q
��}��4j�`����o�^p��z�=�tIۂy�~�9��r�J�N�=���i�&0��QIGb�]|��UEӱ�I3�ψ/�,(�k�����)1R���qzՉ�'
�����:���S�aB�5n�{rlh��*���l��:��0�X�~級i��R��uZw" Bݢ��gчJz
�T7�U���Ev< ��SZk���v[�A�� "�f������@o7`�����P�ƋxX���� �8Ć�H8�����br@T�/z�=7�=�5�t����]_6��oq��W9`�Ǟ�}����?��b�٭s�7S��0�8/��<|�# ��&o����#���7,\&j�?(.�/T�g�7wN��屪#*Bۢ!VA���fj���L��6(>�̵��}��8HN��x}�mn׋�(�:: e�F���=&Taa@�������]o�y�- |P�s,\��q��S�������,��1���)M���n��'�y���QY"�����N��?c�U�����Pܓ<���8�U.ns�ȲM�dZ�%i�X�?�p�Z�#I?κ*�t���ި���$�6�EZK��J�@|aX3"�$54�R㴞%�����J��g���z��ptf}�ȜCg��<� qX�{��I�ު��e��G���I���&v�%oO?��J����9����5��~:#��1�p_Ѵ�w�T�I~���+D����8�s~�,�Q$;6�6�.Z.%T��C�\����~�s ��ѥ/�L�j��WbDW�0K���]�e $x��O�������/���ݓ����]'�P�X��	�,���>Í��T�}�H;9�9��M��!I\B�P�.S�Đ���6lz@o�E�>��򉈑­���̳�WCF�1�w�f4|����L/��M�=�.p1��e�?W.v�Ap�W]��.Sw���3nN�Z��
c�h=�&)
�P���[�ZkC~wzd���W[�E\���F,+;C�|�s�.�pA+���]~;I�<xؓ������*ˉ��B���U�OH���]���/�sS:I窯��Ѷ	����֧ߎ?�.�B��p���4㏻�n$��9��tԟR�F:��T�m���( ���z�M>�^��4����|�;&�C�,�׾z��r��0Jd�jew�L���ʗÆx��������'���IEс��)�3/�Q\�i_��Z��Rӓ(��u�"��U�*w��˼|kF�*��$�,e޽�{��}�h�|�7�tB�C���X@����w���~r��Is:N���K�C�OCf=$�2�_�{�j���P=��Ѕ(�<��6������}vMo�c)S��?�R$+����en�L����]'�@
2�֡�a�M@��~U�j]��	��޳�(:b���
�.��yx!v��������X8������Ȳ<���i�8ݾ��Kv��U���P\4G�'[��B}	:7X�9��jZPy�j�N���,� �Ǫ޲6N$���\��[��K��$�e��/v�p��d���D��~����4X7J��d���pU��������c<}��왶Gɋon�{������3���4�N9R����&pTw��C1J�$�nۂg�$���ߋ��b�.���Ix�6y�*�uZZ�������.J+Þv��F.Z��d97��[�Gw �S a��`q�.�U�:�����=�O��*��)S����ȂVCG�����Pz�Ճ(ω,Jk6~���� \Z��Zm~O�[��5�k�{'5��o��|sIh�F.i�MO�Mp�7�l�Kxc��i5���Rn�>3����]�gR���㳀�@�Kꠇ�i���KH���m<D..-�;B>J�PO���fp9��8(��Fp�v�4��n��/�ԁ��y9z��d<��)��wy�t�+P9�2a�~󞯔6��.��;�ƶ�,a��HL�7]�ŝ�l�ߣ]��sB�b���(7� !�l�hģ��ZWc�s��^���M�3�������Э,)qـ�1�G#I�,�1�o�	�c�zܚQ>��ρ��݄�݋����-,���
A1���˯��,CUl���U�y��8󓦵���hl�v0�q�$$3�ܘi۾��H5�T��i���������vH`UdQAdáY�xnA�%dJO��p^	���r�=�}���HV/���I��u������p	UG۪ib�z�a=��b�'b
x���g5����q��NԖh�����9'}�t*�y 6mo���S�m	mq3�eB��P庇_�׷ɴ|�(s�o�i�����a�<8�C��e)Hy>Sl�c�UXΐ��S9%�0j_��`�`�;w??aJk9	yy�M�*�(Ą)����S3�T�i�ts�-j���߰�"Pg��T�ꞬI�N���5:_�R���	Ǆ)��,���PN���ڔ��aT&�т2_����_-�ǋ� eQ>��ΥDD�_"���g/n�QB���r	ZΟ��]��=�>N�Q"bI�B���3w�B����ώ�#H@��D�^v!3���
}l2�a#�MKH`��B[���`)�W(}�ky�3�u��[7��.���ˍ��o�(c'\�L( �k���q��u4�1áQ4XSe#Y�(Q�K�F���]6+z�e�j�>��ۚСD:��60P�É��Tݕi��e����a����Y:�b���I��j�ԭ��:��FN�x��C����p����������]��%��hkj����QQ�wf�%����0�0Z���S�#��;�! H,�$�b.�'$́�r�1 #+g��Ϡ)ˀ'?�*������^���_�r�Oe�/Y_L_aq����i�,�Z(.l�|V�����v���/���"������z���w_C�W�׍���Ϋ.`0�<<о`���p<E6�a0S�n�yľ��k�����+��k�θx�;���6�i�7���b�~Q�-&G�����5�r�#�h�Q���m<y�j�^}�#Ր��s�?�a�喳R���V��.�$��ڭ�
07���k��퇶��l���H�7���>�=�p��D�p:�b�'$�� ���E��ϮkZ�3.!��4�����_�5#XW�3�j�Oě?5�*��n��&��~�6w���R���BK�{ܠ����8Ԕ�w%SWSV�u�vM�f���A��x�$�e0��A(�K���fѳ�H�g���u"��r�'���p��g��n������������+�;���o��j=�ْ�F4�ε�I�5�:��⿃�����Y!%�} �ex���ȧgO���B̅���U�k��3�j"*��XB��djcE�z�In{<G��ҫR��u��%mI(R7�7Z?��Qل˹���d�qV�/Y�*�� >PLaef�Z�<�;>VK�p|r�F[-���G1GP&�uGaT����)I:��;b��^(�������^��qN�_��9˹ ̱DOcDնG���Ʊ=��刅k
�?Ҍ�)m������h��pU�[ގ�G��bs^�:9D�Yt��I�圠E�Ա�3!�c3ߠH<!\b>O�N���8i!�I::	C�E"Fήs�E�$�8�j�@�ޕ��P��1w����1�B3�k�x�Ȅi�=XA0�a }l"ꤛZN���*��3�F�B���z���)���vS��:�H��w@���l=���i�� _q�,�]��f�"��ur(��0�}�����k\�����O{�g' �6��ȎB�"R��LCI��>|�;�*���c6����Q|銕��z���$���UF�,r`8jD����;�[��x�_C������2/�R�Lͬ�^x�cK�N�	��+��t�s6O ��b4ՁJ��2�3�7[_F������"�\�fxd^�3����P�6jT�M�c�t<��p#	`�U/��=��qcA5��u�4��G~��g�^4�����9�uִ �=vJ�j귧�d�·U(ݸ~{�BR[�a�H���e���0+-�J'�1"p#U	�;���iK�K� m5A'߃h��P�i�x��X�a� ����`��)�ٜP��;�s�җ����`^���w�o�ۯ�@���N1#G=QVf�*�� ��6=���_�ܦ_1�Ѐ���G?���H�GjeY��:�v�q��yH6��w7�?�K$פ
����b��#|�N$ክc�.}���G]#،<��6�`lL6�ŃL�\���541����D![?�XF_8��v�� g��Rӄ�nAZ�����-�m���V:����l�0�K��y��-�j�٤�g��{J"�,�r.���?K�,�%ڄ��V<Z%��Zu(�z��!����8PS���������M��s��[ɪv�Y���˅��˗w(��A��7}���)q�l��LTp-�4���X	��x��� ub�6}&L�����b+�O�Ɗ����'&t_axE�e�6$�AL]R欑�8�S��W�N�8T9���-�Uq��辞D�*z�����|*����~Lm��$0�W��}�WϷz�5�aL���/��놱{���>�o�֎��R�V���=P�#�r��Oo6��𒫤��|"�j����̓�	å޶tW�8������@]k0�(��SO�ʨ���3�5����Spa���ܬ�K�6|�i�Y܄9r}�)�kf�����yd����\��L�9��˽^�������n���9�8\�QP�E��7i�1�2|���kT=�7�Q��R�����
����D��r�W.�>\�z5dz�;���u<�!)���{R85�6dt��n䡇�I݃��vi˒a��CD�xRC�����&�P+7-�ka��S�{��{��(�a�nh���u8�L�Yz�'\$*@�0�mI3U����"Xx�s��ڈ�]��` (�Rr�#> W��S4�{���8&q�'l)Ã��Ϣ�i+b��fǻ�@�u�n-@�XƧP��-������u��M�8!;�O1��+����wW�1�ubm3��K���KzK{}x�RgY����Sq}9T^�b��ֻ��d��M���t��O�_����q�s�{l;��p��v�!3��n#\'O���I��t��7�Z��4	�/ɵ�x���&��e�դT¸>��榑��D[��{�=��^��/�D��labLV��q�9��ә>5%���Y�����,���"GW�N�(��� �����G�bi���~/͟�!s�\s
�^#�*2!0�3SU0��"�-4�U
߱�l>Nh�rl�x�5b�$�O�O.�8`�����$Ұ�10�͒Wf�9-��;�G��RQ�;�Z�05�i�"n��c�]h�
�.,->Kz}3f�E�p]+@F���i�c�v7��H���F��!A���T�n̕�~��*j�F�� \t�X���]�)��V�{!(�ei�f�tǨ�9_5��S �Ѩ,�X�o��~mK	)���
4GVA����|���YPfDe����C[���==��n�깝.�|M�{x�*#w�|�+���7�
}:͗,�[�$o��yg:-ph����ve2S�=�rX5�'�@��{�v�2@�a��$�LDC����	������<s|�Ax\�ˇ�靟U��O�R5����$���󶎈�aNkv���w̄>����~_��������Y\����=&�i˓�f_H镩Q�Q>�7�r�-�Q��n��`[���]������{Hl�Phb���=�L��Ycv�j, �@���]�K9I#���V'���&Z�?#�f� X���-��M��+V��ةNB(��� �<�T��e�vT��Z�Yn��:(�ч^fJ%mZ$K�	*���U��9��C-a0��3����>y�5՚Ԥ;��E�X]�V�q^Ǡ%���c�m ��J���|xTëp�֠-cq{s �A�G;!.�Z#Ь��G��
GW����4�F��_�D�"Ol�lB��v��t �q���nw��R,��~{Jp�p�+�� ������*�X�EѮ͖����bY�pG��'�tsꪈ��OX��*r&G� �~�@�����\���lX$��
�4��N��ۃ���zޤ����e�q-�ߏ�s��&6�l�-��˭���E��"|��mo!D��N�9��wnhÆ�r6��_N�͵盖{��J��8����OHż��MH3���/E�~��lJ[��a �aج�1�{�lsQ_^��	�sm#���l��p��jJ�߾lk��_��K�ԢR�ɚqY�T���X��e���`�(/���x� ����RՓE��8ʖ�k0���i!8.n| K�c7͎��緣�Q�(����e�O�*����~(��D�M2#�Cv�T ���O��ϝ�"��~��~g�wک@�~�j"j ��=�^v=�f�b&��w��R@���ߊ~���Fh����#��4�ƿ=�,���"��Q��Nv˻i�PZ�)�'���}�����$6C�X���̨b\]I���˨CL�O��:ш����X`L�RjY@)?�f�g��k����X h���$��G�Ȅ���v[��g�U��I
�樇Zz��L�%��k�xw�,R�Y2}^'�S<y�*?m��?;��;���M1�C{�f1 ���@��6��9
&�RҎ�}�!9�B7�D����:�jo� 1����L��p���3|� 1�`�&⊣���9i�cS�)���fw.���=��q��s���:v+s�-EG���9"yq6(A7+˧����f�l�o�u���"�2�M�-lmsʩZ6�c,j����T�洜-�*L����oYl�����1�0�+P�_
*�xJ�_)��ɹ|N��݈q\��f��W�h��Md^+�"G�Ax\�������>��v�U��W�!����֪"��n0���dL�lf��w0^�_�n�\2h`�n��SH�B�UM͒_�Ǝh�2���5�xd?#�P���g�f]��ִlҹt�{^����͞�|a_���.�w�.H����By�_{q-|U�{�̋ja�=u����ռ�F�L�p��j�3^�P�	cUQ gii$,6�Z�1W�0��Й���[�G}�fb�K�a�hn:
� �=�E������YW��Җ����q��0 �Qf��zp����nj����(w{��ː_�d�,_��]yÆ8by���ƽ�Ŭ���[͓�Ҍt�05x�M��\!3X2�2�!���s�4Y��P@�5&�)R0���S�Ib�>��8�r\��B۔�[�y�L*�;(zwC*�cAӄ�.�h6�`���,T$��
�.����s	6ӹݏ���{��bX�e3��'J�r՘U}��/T>����[�;�`!�}�M��g������BΒ�v����+tC�g	;��'Z^q�H�T��B����9e�E#�K�&Fa�"�Λ���N��U#�|If�;�e�:.8{``�#[�*��mؓ�C���܅-γO�J�`�:��r�0Hk)�+�F��ok8ճ��m>�;���[��bLZ�L���䋷P_l�M��N=]
� ��x�@m�5�t��v_���X�>Lλ-'!�j\+ق�3܏6�w\H��{�4.\��+W�|B,�=��Ԕ�� o�� m@$�Y�+OP�Rf�7��M�����T}zl�K��"ː�����{�X^7�*��}���&~o�+�V��|/y�%�?X-�a��5��cr:����1@ȹ��m'6� ��N�zߜ�AW+X�c��a�F	,�{x͉���z� �q�dw��2e���R�T���r�%}�X��p�{XS(R�ؿ;-2��b+4��Tv���?G��V#"@���S�Y@`<f�Gkg����1�ƹ�X�CФ����!���D�;�t�@�.�aEl?џ����E�=�Y���|:�:sv�\��L #Nl+M�v:#��/-�|o)�����^��+J�_˼��ʆaȁ��ܚ,6sq��w]@���?�[ol� �/�4�9M�|�^��`S�=wU˱[�H��yaid:�6cw����A�������� >�o=_�j�F�^����=��u;I�E%�b��|�e��!.�~�(�G#/�qѬ. <�&�h���$�h��tՏc#�C�O:�^q9�� ���v���DH���Є��DI���Cd�e*��9��p4"νa�4���\6�~��g0t�kPwl�{G��d�f,%��m��0�6�j�p�΍`�{QŊSsϽ�}�'�ۻg�M��VWLկ{�B@>�0D�h���q��@��q�����Y}-T�0y�ǩ[�0��"��3�ūpں�)`���oy�j����}3͞�"M��V����=���n]���r��*|��qC�Vވ�>��Oȵ[��3�G�B>!���el	p�D9�4����f��lCM�>p%l9��^��[��\�,I��m ���L9��&��0�p5� ���M�`���k��t�+��0^+58.q}PFA0�&��H�-^�<�#Q���`��T��o�|�l ��k@�L�R��4�W�$H%9��]�iz w���+��M�Ҷ��Z�d?�8����+vyw��{�V{9��D9���j���=��E�R��b����>H��VN?��(pP"B��^���`U��sA�
b�!���8fe���i�v�@�O�gKu���eL�v�$�A]��h�JtBe���.��7�}K�1ѕ�M�W{�8�7�����3��-� dQ���;�Mc=.k�#�@S���n���G.+��u�/��X�~��1�1֒)V]��jU
Vp� �d��`�2v���P��h��!�WԔ���)���+�7��C��$E�"�)�= }�a���k',��p�Gotw�.\n\�F�D��4N��O�Uܒ��]�F�����w���8_�f����b�%��fk���A?��T���^�9V��ݏNxxU�p�&:$v���E��S�ھ�
ߡ�| ��W���ņ�vYӇM��At�EF\|*S,�}�E�����"��S�<k���$8�/�ՙ~�m��)�y�x���/3 ?ȁ����7:Ja,�R/�%��0����wlӭ�i�[����IlU�-�	^����1��g;?�Sd!�g��=�R�[y��+/�-g����i�x��o�us�'���絖z1�#� ����	e��,�?9UF�4�6���IOQԤ�'�a����&�Z�&o��!-X�/4�~�^F�sh^��',H�ꬳ�r�떹|��:���X[� ͵�Ь�³�-"�Qm�y ���p𥳐�$�Ȥ���ԹT0��C�6�yΈ�zX2w����.��c���@C�@lx���{�!��KR�%x(0�VU���eWA�~@{���ғ
ς�c�g��^S����b�	f��E�Ӄ_����17����(��f���̏�A��ָs����f��_�,ӹӔG�"��t��y��?H�zQ�;TC����і���:�%��z�ߊ�~cPel��n��qw�����Ы$[�%_��H8��<��+�.�7It /L��ATA�2G�3$��$����x���z#_��@��c�>eލ��38Gg$а�B��!���0JW���u���$Q10���g�O�4�p?�U�-����� ����[��"�ט���4�.�K[J�]�Y�n���
�g�Һx���I�b��R��Z=�RDJ7������՜,ײ鮼-�adMU��hva��r̵��Z�Z[!?i`E=�����Rk��A����Ɍک�K0k�̘�	! ��d�H�����O�c[	�����^2pʣN�1ӑ�s���ݜy^�W([j�E�>Q���E`m��)$�W��˧�Tڃ"�?n_ٻ(M��%�c���E�5Z�z�,b���ЋlkH���G�L������ny�	\�#a�W),�&F�l�
�6��cP�Q���|;J;�@�!�Qq��Q������ͅ�	6ˡgz$�^L�뺽���(����?��B��]+>Pсz�Uy����⭯��YhݠG�h���e6��鍑,[e�p�dݹ���f@&��^^NA�'(e�X��4Կ+M@��AHa��^TÖS�}�]�[����i�WuuY!Im�MyvQ��Xo���j��ag�0�, ɚ�\���[f�j��c�����m��5�s�������Z�F��i� �R�r4ˊ����1r�h.IL�5{��t��.�G�4�
�XD!!q����9
�k
�V�� �C��`�voy�[��I		���}r:�������K�$�--���@����?�ץDJ��V�%N��T�	*V�3&������h'6��%�r���$�$.vz1v���|���"�H��=�I����\�ߴ�ݮkt�A���t�8�dD�Q{�=!�ŬJ��aNCf���R���:�����Js�J�I�U/�7u�4�#]��'��c���	�^�U� c�	LՂ���2�)�
X�DQ�[f�{�������?�r>>.5��.��h�hHS�K�.,"�?ng*���]>>�CJM�Ш��֌7�b`���Gy>�/��qf�9~#�0Q��ָot�B`v�"��������T�������K<v����j�_	Nu�9F&;�)4���K:�K��M�S����#��o6G����o�:�C�rt���7�����C~%=:w*uhD����4�f���JH�=�oH�	�����Ǯ��j�b���i��`s������AD�ux�.�|��P4⾪�6R�uC�E��r��O��iO�����fDƴ1p7�Z��h~ݾ��dqCE�ˉ�2eQ5���_1b�T����S��Cn%?�0MI�==���i�$��I���'Dz�SszW�j��h�n�ai3�"��層&�`��rL����r]�2#	��m'h���~�����Y���}��zu8��}�j�s4��Y-��Z��������]��B��L^�l/��[�C��㍠C��ԙ t���1r}~�1�@�c�F�X�"tO�U���-z$wE=����0$biNy��v�,~����P���vAn!8�<ρ�'�ЎӼ�SLm������9����c7�MY�?$YEt�Q�Dϖ��F4> LYEF������R�sf&��z��'aG��w	�����L���	ܻ��US��P����&5�o�Ž3v
�a\���.����M��P'�+��PK�ܘ| A:��>��p��e"i�j�4<�f���S�)�m����#�m���p�p� ����[̎�0 ���b��8��<c�i�3	�kg<s�Q�vR״��p��MV`�mM��T  ������8P����s-`Ԥzʿ:�zbօ4���ɵ�K�H�}�Z��țJE.=��U���l�-�ߊj�	�^tB&��̝���n���/k�|�U ���l�j���5��~��*�B�e��&��D��1GV�Q�.pLڎ��d�:���V�9f�5@�����PZ�X�G��Q�fߞMZy���v�FwP1�ч�q��HP�����ħfU8�	CDvT�[�7���8\�k�]�xj(!hʢS����5���]��6���M˯\6݀�W�H�UgǺ����EhU}�p���6
�,�4�n�U}'��s�|f�Z+� Me���^�!���m��v0��Uʺi�ݭ+c�eKJZ��ѼLߡ�8̆�
�y�m�Ui5&e�������Sg�1��>O��LsC�$>ې��M���1Ҕ���P����f�R�J;�fB����á��Č�kt6��"����	>��:���^)~���}�.�귒@-9K���j��gJo�]�s��m<п-�㣏�P�k�ݼ������|��t:mQ��o����H� '�/�
�Tz�EXUd͇�����G:y������2�,"`|�l�-�%� �O���� #oS���
�g	/|��R6z�֐ð��]+p�2� Ay�J�+ }�-T< ���q�)��N]J~ށ"���aW(�s
э��6X����oj��
-
���������0�ł�B��hjJ�Ɓ2�\���y�b7�z��_1�|���!����cI���Օ�S�w�M�y�Vݟ�F�2z�ϫ�9����ϣxj�J�ZG�����֗b��r��xvE��al���,�8�B�bK�����%E�J9�F<+��֭:x9M�k;�#������%�n���\&�W�7X��*����G�ͻ�5Aʨ���|�}�����4�|vEL:�?��k��^��:>�5~P�Z� �"�Q���Z�~�}C��(|lT�-�AI�@��tD�~/"z�d-N.o-%���%��@���~�[�=�C���S����
��Y�r�ZWG;aJ˃�[P#������%���- f}���0���b�����Ж�dA�?n��O��a?��N>1�ʀp���7�Y>	�𕒳T#9�d�Xw��DD`;�s[�6֙ .�s�Y�d8���Rв����;b�GP����A�A�'�y�<���{-��.k��t r�4<-�W�pK���9��P�܁�D���E������1�+��Xw�r��tT���#M�+hѪ2���:�$b�r�(��N*NOmL�iA>��>�����ּcd�_��M��gn_�m�}&K_<�70ց�N��H�P[9q�$�������O��]��Ñ�{y�'�+-�Sō��wF8<�����a��
��i�4#���yD��/Z>�s���	N���!M�莗2����Zeq�oo���d��/T�A;�EQ����|��Bb$��/m?�y�sw�;lvV���w�r�~������Kn]mFaX�x#fhee�\>�-�tO�x7�vd�0�@ta�h�/B���j����Z�N��T�tt�S^���x��R�Fhq�H�W��T��U͇��\�\L_�2>���η~h������'d���V ��~����|��2x���D��M��b5�6�0���Hu.
��!�_�+�%]N_�=�w��L[��a�@���f·�$�6dd�����>$1 ���A�җZ��p��P�箃��:=��J�Ե6»��5y��P�aJ[�۾Mo�נEB�������x�����8���P�0�r��L=���&	w�CH�J$�����G9�+2�F��x�����K�c�q$+	�~�7�������/�B5fG�w>f�������ʈ���}��e8��P�m�ŌB�K�㺌3��q�2�^���s�7���1���xȓ�ڱ,�]zQ7{QBU�8���Ģ����%��t�NI�S��m)װ1EP_��bm�t��q����1o��}4Mƾ܏�zمT]���I��	�Β�͜��PK����V��I���!p�~���fwI�!O����;��g�>���g��)�������,7��Q�����=�7,0S�����- |�<���3�*r��3��Wqz)�vj�h�d>�#l,F3�^��+������ě
�F�f��@aD?�dxJ��&��0�,X���e�b����Z�@��Q�����	�V�ҽ�3ķGfU��I��|D�;�:2�E�Ԭ����qH�P1��=ƚq[��&��-��[�u�����˗�+x��2!c�>t�e<15eRP~�لJ`��sv����0��Lvz�q`iգ=e#��z_x�ƥFä��P!�=���FM���v]�9�E��o��g�YXtJ/9D����M�SW�V�Q=���ס �-�����d�w���X.v��k~�翑�
�UQ�XP�U�t1�8m��:ǤY7&��Nr[�{�w2\��mm�{�Z2�G_ݱ��Z��Lڤ���CCx�d�W7�6Wc����;+����^��Hj�z�0S}$$��?	nE������*���7�N ���-�Ȍq�ꤴq|�o�����>�`�Ɯ�eҸm�ΒF!���T���&��S��5�&�c F�k#\���a0������q�����P����V����ݲ�(������n՗�\p�d.��0�-j����`���}�ҚL���M��\�/�r4�zr�C	f���G�6e�p&�uuC�K9���2:��Z*����}W��2�M��%j�=�
0l.��$tY�����$��M$�X������r��IT�PlɇS�(F/c&�Qn����f��Inܯ�K�)���̝U^�\͝L�EO"iNW���ĠxUi#Cͅf���^_��H��!t��W�$hçA���[��>;+*�� S���$����G�u[hs�J2^I�������3Lb��O�/@��J�U(�2~�F8�0t�곭j��7�>:�A:��F��nH]ʞs�	���F	�B��^���x#���m#�YuԸ}N�
�mm��{��]I�Xe��µ�|s�G���c@UjT�i�������z���T�n���zh wD��e�w���&(�d}'Z��Vd���60��-��ؒ�wjt[�u�
�>+b5R���߾"'Ͱ�;"��HO��C��ʟ��'ɓ[77(b�A�%$�3�c~���e��Ӊ����U҃�5|Q�u�^n����a���S]�rr@�c�Ï>�H��[�b[�&M���15{H&�)�|��e���B�t��sY��.�=�pK^p�2-]������J���5��""͗�(_����T�����&Ilɽ
�P����o��D����BJ�m>��;����Zoi�~�E��A^w��
1�ԃo�����Ņ���,v�Ex�Ur/����O$�1|���:�"�s�+�v1X����CXﺥY�ЪnF��L��vZ~�Ȧ���s���G\`��EO�hH�����7$��hGk5�{�'��]�w��S_%Ϲ�w����f�
�K�\��ꂥH���S[ ����L��t`!���]��]�Kn�˺�Ic]B��Y�W�k��<�t�J,
s��i>����t�uܺ��R�+8�8"��0��g�@�UT(bZ��AE�3U�
����=�>�P(ӁLћ��+|
F=��ʦ���*��'��ՍϬ?G�����Y�#ߏ�����JtT�V*�A���=S���y{ ����H��2g�:��k��݌�c���i*����A���`]��1b�c@��ca���J�;�����H��O�-w��`bM%fw7��d4����o������hG6ܥj��, �B����N>��Ӵ��t���3��C�pop}�"��L��5#��U����D9��gKT�^�\��17��ߋ���ʹsa�����C꺰](tj�"�L�i��\	yV��M�%"n�k"���){��;̲��T�o�t�j�k�%/���9�'p� K��0�.���JL�[���b��V�o!t�^j���w��v'N)d��6$#P]���r�y�n��c���o+�F{�P}Z*�}'�`	yU�e��ͤ�P�G/5i�1Ø �T����uU�tm�B61�Й���?9	p�������{t�o\��k��l#�k��mԽ-�K��֕�?M�ֱHgB�űt�jlp�{��>�.W����R��6�~>�LSE�q�hZQ�|�x6V�Т7�R��q��b�<�	wf�nu{'t����5Z�Xn
}��X_[��*QߞP��(�࿔��xé���!G���es5ƺ�.D ��߶&�yP��GH���C�!��<��[�����l�l,�Q�DMY�E𑺶E>���� ��7V�˩�NC���,D��P/m3B!N�̂Ø��Ay��&ԊX@�߀�"!ǌ��O�H/�B�}�j����)��%a�H@�tV 1��t��A�;�ls�۵%�P&*n��J��V�*�F�x ���86�-��3y��D�e��^�cK�u�-�F>�f�t][�0�q��<F�2\{}�sZm�{���@c�ۖ'�{*�)o.жhO�S����a�o�����'T�x�>��PguV�Dl��s��R���Ȕ��@�*�[��Y{�o��%��/�5����,b�.�`JH�-*�뗘vZ��J�Ln�36`�ŏ>��^�b��5�|>&p��D�ۗ#�S�Jk%q�!	�g@Ņ[��τ ���
�*��Y-��x�1o�9Z}����*�}�C�Ȉ��&p;\ua<Gk�a�����K5(#Vk#����Pl��|=��~�U8������3�&�����F^,W��`&otT'p>���d4_KY�k��/h�x��{�pb5q7/��wH�n
�H�J|���j�����+bi��[�>�~��'H�5x�q��<3W[3S/Qk�m�c��'S��|����I�o���ˤ6���MT'	�\=*=�o�_uc���Nb6~��)���y��;��w��鋳�en�q�S4�Ѱ$�o�PA.���%�|�[X@��{�{�zԀ��N����0��u�����"����0A�v���<�Dm>��#��u�N�K��O?]J'~>"D�E�o_�4��3�x�x�ZܼՁ�&z�G� 1Ml]�C��Bs�6Q:�F6������rG�{�.勦�,w(�����hV*M�QN�I�c��Jƥ0�Q
3�cnh���p������\h3�s��x��SUE��2�?����@@�>gʳ��Y"�J@Uqb��'g����ؽ���/����I�Z��;Y; �ſ#
��Yނ٣戀�z�(L�;���B��n�#�I[�Wauj�&3��L2�"�(�p	��1+���i�&�Bf�ld�v�������[��q[q�s�{���0b�VV6��k-
n��A�~���������F8A%ô�,�����^BXJܴ�qx�5�:��FU=�~�/�T*?�ܱ�z�ϑH(�i���G��50��v}O�#(���u�Џ�����7j4|��|�[��-do��vU�I�U����)�{a���y�/��C_�<�-�^���I����k��^8�$��!��!��9])➟\��uq���FX������d����_�����2��h�Wl	��V�g�r��g��Pu�(t�L�GSF�R���:_^�l���F�%�^��-+�X���xEhb9�r}݌�I�n{0qqXi����u�-*�/%]X�g��?�+��1j�8d���t:���
���>���6<�2}`���7�ṓf�)*Uk���2a^�y �܏�b��mof
�9��5�$�s\��ټ�rm�i�u@Z��C ��sa�/��P5�:.��>�������pn	0O��9�묰$���4�>�v��qI3�\�ԏ&�q�R1Y]ܔ�w&���:FK����4��65�-_�&R�\���H�wiIB��[�+K����8�K[��@o�)���^x����)r�`^�}�r>'>�����69��v�òS=4H��=� ~�iGax�@��,�/�
z��~�t��͈�ڻ# ��6?</}}��v@b�����U1�k��aV+�[����ٰ_[�'��k5N�y�/�6�U��h.�+���G�"cRW���2	E���ZVY��7��t�5�|wl�rܫ>*���п���\Yozf6�
����i�Qy�� (92��/\vJ�)4V:�'���W�������{��I5B,X��2BK�5�}}lz�����q��5�G�iM�ܥ�Fd��1�@��溛���ӗ�F��#.��ǂ4/A�hO�3�W����86N�[k)�6��6)�wMC-�&:��L��#���\�P���:&E�g\���*j�W���q��n�����sh�f]�W�ad�d�q'������<�F4�~
7�8yh�2��xk�mw�S��E������k�3���H�=`�6!���C��Ooh�u��d�F��
(`�|�`��s1��G�R9���� 7I4\���Pԉc�q,��#�=夭ƀ?��d�s��2��ϡ�ܟ�2!���F���9�KxWG�/�  %��O���(�X���F���x��\6^mb�.��qӄM̡���Qt~0^�~WU�3O8 Gc�"��BV�Km
����}����)�mƔEQl���	�H�{/����s�ۘ#��>s��b��9i��Ta�_ҕ!�H�*���V���tݡ�Z�n4��<�G�?Y��3_�(Zma��s��U������+HdQur1�vvսf~��4�cqo�_y�/�}����6A�׹$k�Qbv�53q��pA�9�� 4�g�q������"�>������5b՗ $4���^�	�����R�yOY<���0jt�.�AҼi�!|s��?��$�H�0�5k
T�#$��B��~�>ή#Ty���?�(���zS=4�ln%-��̫��Ǟ�0�ow|��[���P/<
��Ǥ�驍)��6n��xߠ��/��It2�}�;Y�!� ��g�g���s�@���#6֚�|��ș�`���Op��!��nh�?ny5����uʺ�h6be�]o*���Z'H��I����!5�X�����(���3K(� ���A���l����t��N����m�%8��t�������E=���]bU�n�R^ZS8��W�O���؄��.�� �C}���4Du�td���T-�%�����e�a�90r�c���G�UV(}����>�� M�Eg����t�/�>]���Ƃ�~ �Vw$c�¤��?�{k
0h��;�p& ~&�Ȧ���X�������|�	�a�O��ux�[��Hx�8��0�g���3�[�Ն- ��x E��m��ݥ=�9�u"8� f�5U4���X��:��Ҳ�����������.֩vkU�j�-ה)mx��??��uO�I�{/�
�NFԋ��{��O\jq`t��`�� ¡��E�w�T��{E	�Q(���Ҫ����$�����G����M���x�P�f֪1�Ac�**X�H6 -�w��=���h0i.�����Z�	K2||��5}��|V�kK�a�-6�8����ʛ�$���z�ɰQ�pw����:��p
j�%��e@?*�$@͊;�e��i� �!����s`p: ��x@]�!���O᥀-zA\bUJ����m����MN�QNN(����yK*����\敪2ȋ��l�c�̀Ý��C��a��A�P���6/7@a���,���c�0W���\X�S�`�ne��eCV7���$��S�I�]���`��=�͈��N��C���5�3��j�����v��A+��Ncp�<>C@J���WeB£����2Rx
e;k���sE�
l��Y.�R_�	�f�MP?`�����w�����p9Z�������I+_�a�*�����2y'N+�����cp@�1��~�Kh1��^n[t��(>Q��:�����qll��"�e`/�&0���
qE��Մ��`1�N���	ɱ�;1�r(�^��U����hQ����:�G5z���i���ד7D��o�q��/o$_�6��0����>��u���S��s_�
�����\����\���0��[��8k^5���E��Y��6 0|ej�J:��}[���57�'���HI}P�lߧ9@M��҅`^�5�ŴIT��t��%��Y.�D�{?�����7U{qm�kڳԿB�e�&"��Sz���G'��uD�_���Xx������5���%^R�)�l��y?X'�>��ynd�i/�W&�������l' Ƃ��X����X�ߪ���d�[u��,�DFs!뜛�q@1 _տ{ԩޘ����k��]M��oV*��p,�W�&��jX�N����{�T����䙟._��W=�Bn��0V�4G(�|$��=�K���?�&G�>����Y,�z�*���	G��	
K*�~:�F�25&���B��vk��DE��04O�����#�(m���3=K�i~�;���Pl�Xh�x��$��E�	������ɹ�a���y��>]��𩖫¼�!r�����"%�r0*z�]Ã��*�#�M�n�X���O�e��g��a��_��qc�J}5�����c�h�OzV
'� W�J�:R��&F͝��8vW��;դ���tP�W읈ʔ0}��!�������8��!z��F�i6H�>L�5����Y}1��vz/���1�9�B�1�؈-��_(���7K��sp�!h��Bᐭ��^Z'�W���9{6��bjM�|B��8ՆЙ���[v�W�ܔD�T�w�����οw�����h��S�i�L&�:
+�!�?���$�Oؖ{��a�A�&>�*;��flɯ�[O�V�����E�0�+-ͥ_�]u�@�t,�9�g���Ӡ���7���k�m�dd�J�#��Mј�W�T�'����F�uЃ�T�~R�S�ͷ��Ja��}��g�
n���h1�7"��H���,��^��MzcvF���;,N4��U�ΐ�q�rŘϭ�o�#��eS�?vwTm�ֳ����k���;\	p����j���C1�'���J�[��iW� 
v���s�y�F�D< ���[����&)��'���>gv�4ŧ��#�j=��\�74�(���q�[L9L��I&�LS��;��n�#�� ���5Y�������K�(���E@�X�ҙ�,k����d�3�Nn�� <O�9x/�l��<I�ݟ 9�nۿP�!q�QbS~&�,UN�!�=y}��b�W`��櫱�T�������.�FQm�G����%/�71xf�����(���õ��Ep�MѶpN�]f��`�����j��z>�{��tp]zIZ���t�cgbHI��!���q�መwe�,�B��1l���3�F�m��?��n�y+����
�;\q���2䭾s�I����N�>4�Ҹ\�s?���f3ًܵ�^�X�U��L�E�;���)E��47}��˝Lo����\Z�w��1z����:EQ�C�����vrT��	�g�;���e�j/�?|<\l-A���z�U�Չ���M�נ+x�J�;����:�V�O�I�	�?nz�Q��!�0�BI���+d�a��d�eiP�<jA"����|ϻԯ��	v�-�d�ʢ,?��|�o4u���S{�b�7ٶP���r'ltz� 0V�]�6~K=dWRj�!C5��
����a*-�D����vcaN]:4�-�0
�����`���g�
�ag�x�K^�:���;(����䲚V�L�:iѺ������F�xQ�- ���_!��ȩI� �H���v��X�<�@<��S^�������5)����I8"��D#�8�5�[^I0󳑺�rV#g��&����[G扦sR�/ɮ`jV�P,%?O��L	)o�$�1;;�&��il�����	���хS��D�Dm�L�a3{]����E���J���{0ӈ0�\��[���\�d�g{�z{Zc3�`��,��v��C:Q�*a��i����8�}�r0sd�#5ּz���!R��`
cM��� ���/� �t��	2~M��&0�2��kI�q��xy�E�]�n��$���}Z��sF��źa+Q��M3��;��A��.0ȏ��LY�;xe�s�q��e��!N�I�7ږWophT��@��U���K���� ��6)�D�O;*׮-���B4\Tt�Ў*h>��ȹ�$U�Γ���'�ҍ��\�WO u�����ªz��N_���N��XWƣ)�p���ip�\��H��ZcvspS���U��gJ��X2Ni^Al�鵆\Z$�>Fc��y�Y�"d[�E��T��ڐ�89�,(Do���޼n���jG�,�YA"D����*�Fj8$z$/Vdr`���5^����m�DǬ�Y���@=cxfL~<r��n$4ct�0����wn��L<nrg���N2��J�9]�9Լy��~~j��G-��04��]�A�v�t��#�=�z�ξia]2ާ����.o�1�f�����ؚ0ٙ���`{8噠+jL�S�*Ƀ��=�%|@����Lc�9ހ6x�6|���#aʘl�d�2>�I\mB�`v|�"�\͸m�昪.)�ͩ�ca&W q���3@*�& ����yT�F��fǃxc�t���j2�A�b 0���pGF�;�?�� c����5�����.��{�a�b?��E<�Ѥ�;�h�%(�ξ5c��
�t_a�)!�d��
i��r��B�܎�~x�H�5lb��Dr��j��������i��}��[HB��OSi8r� ώ��t΃y��>��A���א<�ό#��gV�nj�
�3��R鋥,�[�	^9(m��d6t�J~8�Hn��X[[� �],�	K<�6zk!ܻ�ة%��g�OX�����6��^�t�Y4��(F��������2�+{zi�m�=q���z���z9�$#��R�6��u�L6*���u�iM5��Jܪ�]�F�r[��L�y�����դ�D��]���=uͦ��s`:��n�<�g>����Xa͵F:���诩�d�[Ҝ�Pą���U��ϯ!�o�E`�+�%c���بvg��0����~9�~��^ֿ1�v�'m �h��'�SG-{W�l^t#=����K*�dp�0���d	Qמ�Y�b
�旹_>2[�>��|���D�t�K�A�H0d���3g�E�f�H�'O���&Q�[�%��� 5g��&]�)�@`^��
u?K��U�[��'8�t]�ק�#��s��!��H���Ij����Ē�mV�����O�s���״R<2D9��*8'�t��|��&e$r0��1���k�4Pz��Zpc����Y��mR�+�"Tx��/���A�&�;E�ۇk���.:ޢ�C���2�PpA����	��*���k��'��Ri͕W�T�.��|ͳ��Y�A��i�%v�Ŀ,<��9t��$�/�>�h(p��企P[>��1�B���M�Nx���󶛿�|b:���>F���L����#�%A:����"y�q��Gu���@�xP�?��d�rz�E�%{]֓@+��8C�U}���5��2�:��]r��:Ʋ���'�4ù�#�|	�{�q�4��vR�6-��`�^g/�c��\)���Ű$��b>���A�t�UD��bW4�<�*uAz�b	��#	7T`Uk��P�F��o��0Kᆠ�[��<}��аݍ��J���Ag>�.B<��lA�Zs�'j�s�5�/0�GHkt�Ì���5��ۘN#�K���Q��2s�F�Vh��&>V�5�1��\�TYƒDM���jه䥯	����m�ɑ,�{7 O4i�����_��K����D�ĕE$���⊢�D0,b�|�5��7����yR�(^���/�4��h0��H��Jȿ:=�o�ۇ6X��>sv��T�U7�X���~��s�Oچ�!l���9��g���#��%�7e��g+��{K��?Sh�so=�w ��d��ȱ�� w�v����E�Yb�R����PVơ	�O���{8&I��#���^V�P�-Q]i���E�w~~�i�+hu�y�\�V6}�Q`�(2���3]�c�@ɸ7�ǀY����WC�)[=')+=ޭ)�X_5ϖ��^�ŇR0+�b����]�$/<҇a����	���]�Hq���%��G���X}-\�qQ�0  �������K��Й���Lh�:I��!�.9f��p\j1���L���rT��*i�,�@q
�uΐ�|�trSW����BpV�<����7|�"�5��@�f�vq���M�UM�4�6VbW2j��n#���q�{VL��+.?gN4���EM�Ymq �V�� 2�������1W����������\X�ԟ/�^~
������.���F�	)GF�`��~�����8�;���8=Qt*WfFN�a}Eg���dx�+;̪��Y�:�	V���a<��=� ʦLy���D��Q���T(�2$��;%���\�h(,�G��8�0�Q}��|�-zKq����<��> !v�_�����KXK9K�9�X�]�	�WRI��:TGw��6.��r�0g�,���I�j 8--��Þ��5�\�B�N����S�����9M��:���5`��#j* rO"ଳ^G?z�?՘3��ae5w�p�v~�m��uNnm'P�Z�X�����P�:?���׭��Q�j��qe�*pJ���K��aoi�h�E��/�r�{>pМ�hu���*n�Y�FkAt!�rv����9�Z�E�ъI���&�*�Y<�@���v&�c�A�]h�+���Le=�x*����g�^�M�+�%�7]�7�bw��GXB���URh�a(z���3��ݝC�#��K����~�V �����w��˴��Xo*'��AZ�uע��{5Dqo�6��̶�,$g��) �W,9��º��x1�a��}�c�	�4&�E�=`��X?<�rQç�4�s�p��s��e��i+��;`�O��R�d�*ϵx���'�y}��*�c�dvư� �_B��v��T�9������a�`7{j�p�DtX��2����kXf���gt���T�Aj���`A���pL����qMq�F�p1
����\h��W/X:hޮ�ŻSk�J�ضpckҏ�O�WQ��WQ�5^�;����CD����NhM������P�cIe����Um��v\���L��z�O�2���-�������<�	������&��^�\��Ec�PK�g���)�J?Ft�^��3p#RP������ˬ}�R�fwߔP���KR�^�����Q'kZڛ�{1��*`Q���K�3��4��Ӛ,��~�h,�_'��BR�r��ο������1ĒʕX�A%��SaI&����ȕ�|��48�x�ۊ�9%�1Zc�"����k{��!�����t���`d��iO%��>z�7	U����WנdS�&\|�"?�;gV�^��A�{��?�:~>;&a�I����<��RX�˩�K�?��l�ܑWq��Hg�v�p��ɐ^�֒��V%��ZQ:c��~��㬡����fM��� �w�7\� �,Bܴ��B�9�r���ł{#���;o�Qf��n�[}]���OG9k[���+R?y�r*���2ȁa�fڤ���0
X4^�.eIU�4���&;��_�aX%��*yc���0A����H��pѵ�;�ԕ���ex��х�0��P]c(�"S\�l��G譲�|Bt�9$kR�i�9ݦ��Mȟ�]�訩�L~H�L�}��nZZ��[(����k��d�����烆QT^��?&B��_�8���V���L[ 0<?7���8��%0���p㎿`�(�4�Q����4`��1`����%a`=���a8�� �Z�0~�C-@-x�9�_!���҄�Y��������`'�
�\k�N">u�+`lt{$�$�y��*<������8�Ǆ�����s�*u,�*8�͵�\�ξ�]����޽���/�J���G�U��]?�2�ǆY5�Ӏ�n�]d��.�yД��Ĳ��B�;7�����g�77���x�B�C|�.ΔV0�"��.�瀮�eS����=��r�,��#!����14�j��.�o�+�o6X;wjF�m��a� ڜu�E3��/e ��P3���n[�F;GD��c+�%���$4�!��y��:��T�<�^�#C
L�+Gf���V�d�J-83��O<��ۿ������� ��Z"G�;�We�&�H�������٪�f$ @9��e��?i�G�0���=��|�'���i9'���^ͣ"�z��3`����k�(�{���VϨ:7���,�rg^v��{�[7����d��"�ӝ}s� �NUJ(\ XֶWz��5��C����%��pT���d�O�.4�������J��J�&:�|���qЅ�#�)
ȭ
���3��6�MH�Ƞ�6��)�4�/!��*�^_G�h�Woy��dѪ@�֥`�:*�g�f2�Y�� � &NR^�#�5>��k�s�o�ܺ�߁v�}%~�Q�j~��b����Pq���z�ϒ��̾,̊ɗ�u�WS���vpBd2�81�N�z8̆6�����̭X\3�/I�]��@y��\%�׏��h�8C�}R���-�.M��dg�ڌ��h(��^�W�������Q�Z$�ͻu�j*�ӌN�+��=��>����i���
h�8U��,�}��?)���q'//��ZK"4Z�L��8rBe]��q%kwJ����g^�V�� ���:�X��b�\�2�"�qT@���^�v�����=�p��.S��a�@=����,�_z��)�v���VQ��e�����&L^�:��[1i�]S��i���⳯BxS2��Jq��B��RV��7�%�C�ȫ� �!�	pk�(Vj�R�jh1F�k�.���?� �HzΪ6&�h������y��Z���o�s��?�[���m ��m^�%�:\-���q����/��Z�#�V��n���{��:��P��uo+I@��T�5|[B��޴��ON9������p-7fr��'��v�sO�?�,>��.Ou�g�Q$�*ٔ�~��zy�����&?��%�j5�p��N�zl��6�\�B��L�^��#�x*���_��q8u�d}�y-PU�g��U� �������FeS#�?ן�6Yݣ�]g�{&�Ie�aBKn�'n�MN�I΅6�[���/�C{ʬ##!�;]�����/�+E�F��L9��-j�\.��}�c#����c��]���>7�"���a�u���Glñ\��H��=�d�Oe���e��b��@��V�0a��
��R$��P�-���.b���2>��6*ee}����'�F6+c�n�hA��(�߸��.WJ֜������iv�j�/	=ڊO1��|{��5G�xfh*J>潲�º3�����o�%bf����$���E��O�~�멢Db��f�ܤ�όJ��5�{>S�מ��e���6)��di��D���֍�<2��n/�`[r#g󐼿`?�䮨p{Lb��*/�F�M�pM����_��|��3����e]-���]��d�����Y�'tڶ�D���z�X�1�
! �m�?׶D��FG�\F�Ohlfu��KFY��]o+��S����d�Ge�F;\g��#u�:�cqħ;}��6���-@�t�I*#q�Zw��^B��Do�3XDM��9Y�V��8.��W�0�kױ&�Q� �F$���\R�3�u}	��Џ��'�r�Qp��2V�Fn��u:b����H�+�B�m�X%�s�~�v��_pi&P�A`�N`��=|��Ew��"�6mV�9L�xlTfF:Y��_#�д���
X�{t�3�Xك��}��u� 觹��N�9�h5J�Gs��W�%{	���P�**H�%�lvsW��Ê~����t�� ��-C����{p���6Z<�Np�!#:G�u^����JP�`~I�p¤�%���ьX�\�����S�p/�Eu�i��[,��3?��W��%&�b �����.85t�V���ߑ�w�V��#��-����
�$�r�[��%�5��.����kR����TH�?}d�� ;���Ff�� U£vS�Q��l�g7��Vz���]�͖̘Q�di����%��i��1�9���e�u(�zPp���,f�%n{���Mnl;C����ō�	�J��
��p��X��i�`�`3˜�\�~*X-���L�$k~eI�.n����G���P������  9��-_�7q���.b�������-�=Dr��mB�Ɩ�lwQ�k8�u�;C{bڛ�ϐ+� dý������o�F_�3��[��L�fh )�vxď��{� �V8;�@^Kå�:k�j�:d��g�]���bDJ���>��: ���a�s��{qS��ة�I�����&�y�ш�N����D�uˀ'���*K�{,^�����@���8��H�������d'��=�&�=���#��qnpx�sF��Iԉ?�����A���(ar�mV����</]/���魶�t��*���y�x�^��U�"����pm~ ��Oi��0��o���Y��p ��c"��f�]o�=�QkK�6P�������uB�t�I�w���mw1z��x��/����:x��j{D�y�x�:�E��OŗB]2�o��+���L;P��x�m���z�F�����V��dФ�ʲţ�ҍ���l�^�V�Ds,�<F�ہ���}�]�
��^�&�`�H'��u���%8�qr3AsAb��� ���F	���A� ��r)��R�&�H���Bk[]�_��
�����̨-�y/����핰K���!���2F�ȼ�^@զ�M�]L���g� �X+�7��5��ȟA����SL�j2���B<����M��_�x'oB��-�y� ޫ�V�҄�&�,�c	YRZ�<?7�e��r��~��&��7q���q������^v�x��樯��b� S�E��ԑw�?�ކe��2ۘe����UX3��%�~��4��ֻ�K�=;G����������*]q([��/���^�P0u���CZ��h4�U'7��Z[R.�������%_ӫ�(@���ν���<���_<����q�$\�{�)�z����En	Rgfm}�˶Xv�֭vA(��Q��v�.�ny?dG�Nk|������0��{�+Oώ�Y��z;IS��8�2`n�ui����4i��\k���@8�|'�̭�L�H��?�����H�&N�	{9.�lR��cq8⧋)m����Lzbiy?��z�S���u���8v������H�:��{�	u���2�ft���ڮE;�^�gT{�DN���N��J�Ңղ�$������'�ڀ���CN��HnX��&?�O�-�o*�4y��u%\<�6�����oqX��wc�ܒ��M�,�2�b]���Uz�;����h�
A�D�@���<Gm��Ɓ�M<*o���3Ȼ���������zQ+�@7C�}�NR�1��f�@K{ipz�a�-j͚wu3	W�admANwf�rg{�݇E�*��=Z�p%�	���2WG�KW0]Q	p=,�M��+��`���f}U��9����VC��{���9_���SmկV�|YEg���#F�Kz<cY�:r�G�cJ�8��������]��:� ��o<T[ �4>��$Ct�[�F� }
��մjj�����R��{U�:�Y,�����>|�=�i�- X�~���!1�D:u�QJL�c��A���l̑�~(�-L�BxN�f@���~�)��V�)&����-��7yh%Ρ-:tTۅ.��ɝc�%U���l�g�g��Kh�t3���*�/8J�j^�;_�.?3�P/�P�k'�P��q��|���h�%{�:'0W��_^LK[��[���8C����E5��a�ua�y%y}*֖�k�je�<Lq���$�Z������r9F�qN�j�e��}�0�S!|�\�6���kQ�;���N�	��$���M�a����i��r�:�oa�#�+�S:�I��X��d���K���^�yc�r�G�r�#��j�����4�R�0�H�B�V�%s����H|oV��ߏ��� '��աRD��&d�t�)4U�H��I_ѭ�2S����p(S3j[��
KR�+Dia*�	�Wj�fa�u�-�vc����0?�A&t֥d��Vb�؞}Y�FF"3�8���ꣅ�`�������0�tZ�7�~*���J���:����!�X��u3�.Q��y��U��TO�Ʌ�!M��,�* ,�B�$!o@�xpԶ�;���e7�&�Z��{=�����#��U�(���Rb7��R���,56Wn�Gp8,Õ�Ļ.���7�5̭V��y�n�C@7�y|��R&{m%Ս�$;*�#,y<#�"��+�@X�$Pi�8��գ~�8�o��>b��1���������s�V8A�y'�*��X�HN�0X���;�ƣ���e,h�/�Pz`݁S_ThDU���0�wB�ط5H��?�7BM�?��]2��T$L�7��\�<9�Ǭ|�$��<��s�����AY񄿋5�	h
Aj=���[��|������&7�8GR~�$t�����}f�Z�EF����c��?иT��J����|0�h,�}�J��Wrpy�x�TX�n�oB�^�e&j�?}c����
��T�u��}��I((x�;o��{V9�oe=<c��$b����81֓C����]G4����b�f������&�~���)!X!EJ�&f$�"\=:O�z��� zw��R�C宝�R3T]6��3@����Z�9c�$�0��[�Z�kO�wa+/����۵;aT_@:|`hD��r��a)6�^���X�[MWbX_2Կ���|�����B�4A� �Q,E��9E��
,e疡������A���r���W^؎�k�a�@ͮ�e$C�xjų��\�F��+�Y���E�S��y����a�
dlf��A�t3�RY>K�)�!�#�f�mf�Uk֞lu�`������6���Gi�>V�;��E������eu�������{V&���-��Պ�O0|�.�[d����_�]!ҩ��?ջ�=)�{��MW��*�����&��Ɨ�t��WeJ�axxs�:���}�g�Ϩ
��́"��M\ò��I�5��U-�^2�6E��LP��MlӾf�)^���T�j:��'�̟b
�����`�57�]��!�N&��p�T�����1�fj�F�s�X �$ʷ�S��$�R��̀I4�Qm��.����X��O|�����ބ�QL�~�08%���y5�s�0c�$���`��F�f���XO�/N��ZM�-\�/!EɈ$Pp��52�h��vΕD�_��arZ.<I{�
���D����Rҏ��F�A����d&���t<5�%�=�3fƅ��43`ɭ�^Tn|�
���A����bf%u�,�db�)e��۩��!�E�9�FZ��i_��L�1��@8��3.���_�e�_��e�u���H;����PI�KΓQY���U��%�$�F����J��}�j���E������D�i#G�Ȓ;���R�}ڠy����������ĕ�;��W���BP}Ã�P�_�v�R��6�0b�Vl{��o�>�_p	�3���hF2Η����^7:���F��`8H1��W
_+������Ȍ7.�6�D����7�t�W��<x?�J�f;�N��=뙙��ym��}]>+ߤV�t}��Z�P���:,b��y Ux^E@�/u��"��N�/:�(�8���M�X,5�O�w�L@rA`Ϡ��������,�93�D���4�Hy�`?����o]1��@��������n����o1�ʪv�ǝ4�f�K_&���=+p��9���U�M;Y�6ԓ/Tb�œ��9h�<���:Y� �*�UJ�_EJ�]�8���N��?+<`��O%/?��U7o]�&rό�Nk�DZ��_u�
����:�`v�Kx�.��ڂ��,��L�Gf�'�]��p���v�l#µ�B�Z���e}ٿ�����ř�T�|�K���k�x��?Q���b�:<�����l��Zk���F��%p���Ď���������f�<�`츤7�v3�\�`9F�_�l��К�ʭ��e�/&�1R�0�t5
��8�,�����R�����̾Qd���a}��-p¶�D�׹hA��LqM�w�v9s	U���f��EぬzU��c��Ъ���/e�J|/#op��$��'��CL��3yx��������C (u�-f.��Wݎ�-e�-����ɻf|��s���S�z��f(1������S���'D��n�Tj�U�����4���ze�ŕ�j�Ln��h|��_����҈:&�;��n�Ŝ¿"�T�{����a�$��.������um�;R�hm�E��5��&ak�М��ߛ�[_o�승hxxz	�<�3�����F�M7rLCN���8��$$O݋��M��pK[�`ȄƆ #���e�UB*�F�";��z$�qw۳��SRC���8L��mI�r��ݸ�whU����\���Y�e����"?9e��;C��X�'��l��>�� K��`�!o5+��'1ʂ�#1��_j2?��Mn5񄂋���^�l��ZsrMH%�šrL�x��ݭU��t�t�Z���P8���݇1p���@�r֔�k�}�B߬��v�S����������\��}���>3zR��۪�+f���S�]�;Btfq���_�������S�ʺCg-�Q��B�����q�r��ىↃ̇O�gN�2Ȇ�9�����ē1Q���E2<Y���&q+�5��U
%㦥�Z�2���K8�E��u�ɫ����c����e��H�P�/I��g��뚸�!��m�Uڄ�2�I�_����5��ʌ���5���m*oTl#�2&;n���3�h\����_{�|��}����	�,����^uzs8�[� �����2	,�pxZE��n��h�82�0B�p��`�]����z�\p���55a�ʞ
�M��B�K��zLz�܂h��AKg{���f�l)�ZfS忑���`��-���LC�,}�yD_*Vwn9��Q�eS����� ����t'�,���ڄ���'���Y���Uǧ����Ї&E[ͳH����d�� o
���O���G(�\��S��%d�R����g����U:DMK�#n�掩��� G�>�O���(v�(FI�\wJb��R� ��h�
�~p-~�4�ϻ���sT�.a U?�8n�b8�8�4���R��P��ހ�μ��O�7y}��i^&"w��ʯR,i�@�%l9?I���dW��`��A�������2D�G7�����+͝#_�혧�mPd�����eH�ߎg�������5���%
�jt28$��ziR�a"���K&�\7J�wD�դU��Jp�����$Iױ���Y���T<��{�\�M�w�4�k4� K��$��%�S[��b�Q|�����H�K3��T�j���W/��~f�lE9��-�ðH�z�#�Rٔ
�AO�a�r��̪|�Ƴ�Q�$u�^oɂ�yk
"uF����/���}k�INTP�p=xIQ٢}H�v��l��1��{��G|[��1�����|�l�>� ���M~�OQc�u�^}z}FB�8�z�3��q}��M�8C	X�h��%�:8�!$-a�\��qCc���%��\��q����1�����׽xj��R�8-(n�lŝ�(|���c�L3i���hӺы���/l�ѡ�^���r%������S�q$Mܼ���&4���б<�����PG�9��lSs�:/3�r�[����u�0���LP�jF���j�ܟ��͢��K��+��
���N�^ő'[�^��"F0��_V��C�B�6*�'.8�[����f�+�|.��a	�[��;T>oD
7��d�#���������~b�Q�^�p��B�/������"l���������9[7և�뢯§]�9KZ�s秇�.�����-pl�n�z���:M=bCK�QKn�9��s��aDS�(�i���*fz��fp��:���ș�eV*'Z`��P�9杢�"5�8L��y[�W�b�cg]�t��.BѼ��L4P���K5{3�W��Z,�h^����>X%4ۉuDI�ԅ[=�ATIP״O��C����>�ߍ��Yy]g]f�GZ}��4���F�SyV&)%~�Ν��n���ZI�ȺC%$�'k��1+~SZn������g���H<�+TAwS<��i <�T��AV{QT�S�Q�e��õ�*�_R8Z�~� b>c����5k���3��aS&'��B�&����լ�V/�w�������A�ǥxw
�9�T�_��t��1�A �L֚)	�.��z"ȃ�ƾ�����zm2�^��t��Zu��ғ�x]'X>���vQ�����	P�TU�=�á� ���F�D����bta7*���:�����v�Կ��G%S��~;�_�D7�������G��n�g X"��T=,^\�⠖U���Ii�kM�������O4�X���L���������T�~�;B�H��]�G��K��Q�D7��|[_��|��C�[�{�����Du�=�@�1�e����jOn�h�Djٗ��#i�0�b�ы|�z)��϶x)7Hd��]��_��F��T^*-=C.t�k{
x3����NY)#�}8����lL��>K��R��'{�` ����ߨ'�m�����Yq�JL��}.+�Z)s�K�X���3��oLޣ��G!�吧��U�f�!����+DK{������.p]� ��ΩKN��Z3�y����S2S�����
-fz�����{mm �3�S�pm\� ށS�qղ�SSh��8!����Mj'g�v��s����s����+�[�q��z���b�J@{N𗙋p8���FǾd��>���Pr�-b8�m��(޻�zO�Ԅ�jB�L�;`�q�w���#��$��ȲWRFqt5w{��9���3'I��U���)7�[����WŒ��Sѫi��|y�����?�۟�_�>�J�����|Nm��xU�8�wHHf};f�����:�*$�A�t)�S ��D��YU-[6M���*0���J-_`�]z���W�f`8]_��p ��'G��~�w�zc\���4���N Ң&������#�����5��\PՁPq�Dqd,�}�\�Q�2�&ّ�����NJ~3�e��me���Y���X2��}�ٓ��6���;�l�(~�o��Gԭ��L�PaףȭmY�SVs>�K]��"a�&V�b��=��q��,�J���qB^z�w���� mq�C��0 �;���I G�y�!�#Ja�~N_��9qŃ�O%�9~ �4�4rgjԩZL������1'�!�[I�6]�KMam<P�kIKׇ��n:��o�*~�%�sY��֚!g��h�W%x�6�f�oRԠ� _p�C�b�/X�(p�R�-�Md�G{�x�[�`��;�m��{�aȘb�ܖ�^QX��tBQvp��j?<0z�*���B���X�J���7p�}On�T�Q=�ʢ5F��^�Qh��_/��s����}�˅Nfԙ펢p�VQ�+�|2T�^�Z���%�
��(�	A�`���7�NA��w��~�%R]{,B-t�(L�Қ��ې�V<�-]�-D��1�T�8sj\*U���-h��fvO=�����%_�*Kp�����R���0�1�%"�w)d}�t�.=$Q�*��qG.��N�>&]��J� �Q<E�L�����N�D����z�1:u�=����>�z0��,���^���u���m����b&�qs������������ޓ��	C~%Q7)�b'�؏�����_��{�ZL����D��QZF�P�����7W��U��]���z�L-բ��;����8�f?l���@%c�s������5P3sh�s5E������b�lyW܈}�4��A^B�� ���Q}�f�v~-�B�ʼ���@�����f5�IE$���������'�7��V�ƪ7},�&9�8����*qL��|K_<��n���}�QY��Iuee����_���T�ǣ�;�VӨ3�'��;:i���K�|��?k���w�&V�	(r�
���OP� �K
l޵��ڝ�4�vRs���ǨiV�{ �QCk9m��%�wخ�	�l�ߙ��7ND�+ ��R$�	�P������l��M�P=�6��K'0o��L�ߡڼ-����j�1�{ً�ٖ��7R0]�8rݡu�9�#�4Ԥ
1���)��O����^/�T��E2������\u]R�����^�vf����Ɓ�Z����X��Rm�jk++e�1�8�[�����(�vhBy����1�-4>��8�p����d��(��j�+��N�1�->,:X�����(��.�Ş���I�$�zc�*�)�v1�r|���vb��>�+�ၖ��F��q훜ر����rs�ʧ�d�~-j��<�����F��q?=B>_���g\Tk!ʣ%)��V�;*Zh�[$ G�,�ے�M]}F�uր=��Â�A)���
$ߠ(��p.��D�t۰5#��D��J`���b;g7Yc܂́��,����y����-���9 ��o�`^���Mx2H�,@��#��p�Id���A�ړyYl�\d R>�0���%>�\3բ+�i)���.X�0�Vس��T[� ;������.�)o���&^+v#�U�%4&� d�$w�rI��҉�F�Eݺ��	�x5�����kg^**fF��G4���RS��jq��v?'��yG�[�XH����<��P��>�qƆo��7?8Mz�]#>�؆-E��Zn�"
��#sg���$�r�_����kMO)�v'��ջH9�"�
�o{�b�2�
�X4�|�n�/�Mm����-��.����,V^`Ŋ���U�Uw��}@.�c\��%;lQ���
���YPR�y�v/e\������:Ё}���Eud��~V]�J+�Z�ޭ��(W�x��
5&x����%��鉩5�?##��&v�Yl�*}��a���ɣ�K�М����"l������j`G{}z�����:	���ux����l{\u(8�pP�ͣo ��)tb��T{j�W3�T���@v�VԞUpw���z��\�׈|Rقx3�&��6�_�c�N�������ʬxq?x��}��_����O�I�)��Np�e2%���*���G[��e�U�ƙ�s,"茙�5
U��J�Oe�c\���å��ZR99��~$'���R<�e���~;��/�8Wߩ�S��	c��S���q��w)��M�A���Mt��	��4L���ڋ��cs|v����V�"mLQ�;ʁW�L�=����.�0͢%gi9��E��{�!M�)v�@�_�k25\Y���?;�rFN�?��M����ҍ�mp��]F��蜶AUc�����K���@�/�J��{ö��`����:��Vp5��T�	�c�E�b=|���<��x��Pg��:��>a��.O`QD�Uh)3u�"�H��B�fa��8p>j�C����&��QOא� ��=ҊM{	'��>{��J�eD'�!�R��nX$�	nߣ��]�Q� ������)hN�,�V1�� �!��Ƭ"��-��Ȃ�?�%G�`v6����ę���f���̥Ed�U�������a �cA��b�a���s�;j�n���y^�� �)��
@<�<�)���g��qZ� Y�kf��<@v�6��|kIm��wL?on�4�����ddc�qd��+�έ3y�!F�h/�r��6m�{x�
p�^-Bx�tb�C1��g�m��Ÿ�t� 5xհ�EH���tV�	:_�W@x���(D��ݱ>���(�g�v$��}����x�;,�[��=����t.���
��Tﱹ�4Z;�����y�,�#ϯ��ц����7����})�H�k��M��m�j�� �Zj�B{��Eu�m�o]�;(K�DY-�������7�ђ� ��3O�-��[�Z{�*�֘�Û⩰!��|w�G݂!cC�&��lDa�9��I�%����8���UMG��"z�Hm�[��I�ӠÛ%#S��X�l����TLA��.WV��2���OR0�tA��֏�8�9ܶ��#����w�W;��>�Ё�?��Ab�ϴq,X��ԥ��:F^|{._E@L'=��W�3��e�GqH
����oARL�>�%*I�r2зk���Q	�����+c8��"zh�v��#�(���m4L�Dxۈ	�)�[F���<�v���A 9z��e$�&������5�����M ��K�P��j����m݋9�e��UƔ�d�����R�ȗw��=��8�cD�)N�{7��E�/	C6��Md>5�z�V(��_~ᾄ���UR�1'l��Ջf�B`+Svl��%D�S
Ꮂ�d���^�L�����6;�A�e2�iE����I�Fؖ�K�h�3��<��3��U+�r�R��5��
�\�`�k�o�N&-�^r��Q+f��S�r1L��~LY�Zy��;gG�Y�鶁&̿�s�+���w1��iz��WH���WR'&��1��zȄ�]5����U�μ�4N�]�JfQ걉�1�=T{J�f�;��#ε�Q�C/o�Jm�RE�?�TP;���6�
�ʱ3ʇ�M��r��|pN5�ymx���m�`f�XL|Y�T��qx7�N�C^,h�{|�"U᫸RVT|�4d7G3����Mx{�wNo��ۃ=cU�����Hr���T��%A\�e�#X��E�՞'(��^ R̊4�E�#$��tҎ�=r`�P�O--��rl��2��aj;c��F�к恲���>�utF ���(ҬP �٨���?K�zHLS5��Ï�B�!o��%I
_���ʼ����M ���ƅ����}�GmEl��Xt��aߍ�Koڥ�_R�sa��#���|?.�2�NXmۤ�X\�`���w0�ཋ�n�@���F 9�>�bՐ7�+���pl�e���wA̍a4��
��V���i!-%O�_QĢ�W{Ҵ}&���2�#��p�G�݂%E�s�/�t�ժ�����B,�����~+���Na������1�8ӹ��c�nZH�1U9�y�T�(%6`��}���U�*Ά����+_� � \�L
�Y耣Y|޸D��_ɺ]���t_;�/���r:�Y�>��f)��/IDL���w���ꚣ߇(J�M>$����*�~ұ�_��t"
~쐜RV����>�:��`.av��e_���!�SI݇fP�];,���A�6۝A.���-�gv��n����a
*y�ksԠ�MDɬ�����zr1��3v+m��O�yuY�I(��� ���A��O�!�eڌ��N�\��������M��k_f�dVo�k�X �P������%�uuT0�	�_�l��	�ʯ��1�٭Wy���}�+swm�����]1�G�M�"GB�XF��6c�6_�e���st����C��6ݖݡ4+,#S�Z�F�w ��;Y`r7q~����K��E�!����0�5F�8��?-�Q��y)N�z@��\���\P������]j�I��eb$�<�yj��^?2S�t�ey��A�����|w`����t����*@sʽ����D��8?���;P�Iۯ�Ǟ~"N�l��?���GSɻ�`-���qXZ��5f�vh��COn,��0�:pÆ���s����}�އ}\��QŶ,��<�t'Q3~��D	fO�Ӫ����%7�'p0'ظ�!c�P#��P@��2yo��Ļ|⸠�H�ϲ5[m*5���[�Rt�E>��y�r�~%�s@V��7UTL��9��r��47�Ő�sݑH���Fp-���}7�r���LD�U���C�L�O�2E��v��n����Z.ɸ? %x��̄��F��R�~�G[��*���v#��h*	�C'nJ���0��quD����U~Y�`�c����RMu�|pz+�#j�Z��c�������B�fC�?��|  t���f�2M%�O��_-s�t�c�����`y�i��s.�o}�4��0����1��G���>�6*��4��\�y�� 1�שn!c��S�N?W��I�z\I��iX��<�0��@��ri�6ɖM��N��1�:_aY��s���C��;��H-���!`n�Y��	�PKHV������*ε�֔��挝��N��K'�N����B�@!pW������=ZO�=/;ʞ� [�����Z�C�2�q��c *3F��"����",���Xܔ�������.O�-���P8����^���B�?
��0� �_o:�NY�So�ȷ�H�P��,qa�o����z�q���k��y�a{����q6A��T��7v��Oi�0Y��S��?(oY1B����P��@��F1�U�������4� c��$��]�7˴��M�a����� ��D�`&�V#n~.H,d�]-M�䑏O_�	��d�W9��G����,��Zf
�#Brx�<�����haW�]!tc�� ӴȀ0!ג[}���>�O����v��y|L��b��ۊ��60����A65!�Hٶ#Oh�v_����#��"�FU�T��-(,��1����g��yb�X�$g���I�]�W��pV0�r䓿�j��oRʡ�����3)˚l~I!��@4h�6�{w��'����ԗ�Y,�v��/���c�»��#�_\ ���[�>��XV	u��+f	�W_�h�‸=����8Ɗ�/&��D�&��>�Ś^��:��{Ш���WJjtw㔜õ���A��?�+�5tj+�[Kga8�W���0��0q��"	����+�`�̦��g���О7�;i��ȫ./�7aT�'�$�ʡ����i��1�����x��0_���p�V����ё���d�8/�Ξ�'����P|/}���v.��h��uz���V����hKy؆���iػs��zk�J]�v��S� �ޖ�wld$(��f�����[��G�w��%",)XA�޺�-z:��Jb����f��g����Z��
D!���J���WДLLQ�e�<�YRɝ4���ê�K��0�c�e"I����\����,�+r���t�z0��6֎�S�b�{�>]�bZ3���>��qk-������-����Z���F�2�[���<��	����ʄ9�V�E�!(r���I:�;�D�� �~'n@
��n��q�"gn֨����+t)��7��x޼�c��tM��(7ZCށ��Dw�������J��.�F�b�-�
��-kQ��p��J�D/����� ��(��:����s����*h�2Y������M��۶�� 3��l�t4�۬\>(�ʶ:9�	~*�����\�e��Qs	~P2�O����`@�x'�u��;a��z�$��D_�C[P�=mAq�*Mrw�$����P���U��j����ge���[n���]���#�`��A��#iK<y���)t0�f}�ABɡ�͓w�u�w�b�eb�5�?3 T6X�W5�M��1��q������\|~{Z������%�qVf֋	,��Uv�ob�,��Z�MvW�x*n�dIrGn��\zqA��W�����"��n�ڡf�n)ñ3BGme0���A����<�2@X#���ð�tk�:��\���V	���w֝��X��!�Ҵ���f�̃�!�N�J
з/2T#��t�2+J\Jߑͨ0���+���%N�L��ZC������.F�@�X�9B��!����^iT0�]-h�����N��/-l��z�gAB͸Q�q�e�`��I��$ԱX*�C�q-/�L���"8җ�T�R�"�}�j�
G��V�6�_H'����20
�ʶ�{q���a��]������9�1�_�R�͉ 2�SX���ˈ�8��˰���;����UwH-Ȅ����s�&t9���g�?s�'QFi�i�v��eR��cIz�s�c�~��u+E&�j���Ş˾©��E���l'���XNc�U+��}'�󘑮���f`�6C�u'#'���*�s))QJؒt�ڐ�ņ��.gY�wӘ���8�� �@ʖ~A�0ɑ��!�^�5�S0�K,�~1�ސ�m��8s� ����'}�!i�F���j�gT�����k�8�-�fx��5��2� (f��ڈ�B��;\�l�̐����9$4�ұ�mΊ��H�]x�8�m�z�؝�ɻ� 	�����Cܙ��y�x>��r��B��zǈ���@�&�1�	`�7F��sw7��((��b C榾�<��+]���0#�R|���� h��sCV.)��g�Kj�b���\���Y�Z"���B����� ��H�Gɉ�	����ϑ���/������e� ���c�G�'�>�L�F)�!�Qz�;$������lF��e&<�S�kgK���I�{���hb��}�g�V���p�ݢ�g2�j��������􄸖{��!Z��%.���)*�2�܋�<ߨrN#|����[h�%K��7��ɑ����+��#�\ò0CЗ|�6K@���}�Z��{�D�/_����l�l�ɽ���J+��6 �����H���|��<�:���D�*�iާB�|�	XFm��B�I<�ӫwIź���wG�8��e��ԇ�L�F�kߘ�X��T��ތ���U��/�W�bg)�}T)(�c������n��U�:������N-�V+L����t
��Nڋ���r @�hxĂ�B�N-!���3��*y`O�x@>L&R�n��K��s�A6G�65��B���`�s<�� TSl�(ALj���
tN.������GQ�!�]��<߶��:�����Z����1@�8c'�����R��qW���E�R��Ws�D��|�J�{�L��`�l �fQ7�O8١uSh���&uk�FP�|į�E��@~Z�CH�8t����-���$rV�8��{sY�_��J������a������pxF��R��u)_�M~���AQ���~qb�H�s%Z��,1�Eo;����ZQTJ�a�`�CGbV4��|V>�VNkpc��$>,�z q�}s��a�y���9)eS�W�SQA�S����(�Sw���Bb�z���Fe��� ��jzhQR�6;�	�bXD��#%Ş�#�n�mM�x�D�	�����Vo�c�s�;6��nL�³-���K����n� 7yJ�_|Ϋ�Ý�nDl��'�C��>ڕP�؆O��!K�I`Xc&����H�&B)A�%�Y�31�������v��!��>5�fl���L�{���5�;�Oέ����ӯ57i�n�U@�TNM��?ɱ`ΤOT�)���g��(��j�UC3O�tp�Ҿ��5 QXQ�a�9����"�)ZV�H�5p���G��f��g�����S�H|��t�|J���H}��EA����v��&U�{b;Gk?�[�m�v��V�K|G:��Z��:��Gd��;S�:��r��}lo�D �����W��#z���GHs@09s��h;9 ��Q�5�u|F8+�V�_�Mp�uY�������'�i�(��5�C�&�s��MC��V�u%稛h��T�Ɏm�Nx��w������������6��n� 	�wU�0���0%p| ���v�6e<�"�g��H\i]G����2���'��v;�L����Uz'�&K���0!Վ�C�Z��Ы�U֞�g�Hd\p����"��z�s0�u�4g�z����S�ßV���� ��D�J��1dxqQ�ӳ���փ®���j�b�wT<0Ñ�9+hLt($9h�O��N�0��(]<���9kZ=.�H��j�+���x}�%FW@c��Z��5�A� r�َ�s�y�=N�%�/B�r�qZ�fU Ui/Q�s�6g�Ij
�V�@'�d�k! �L0��h�N;�٦OM�OL,����b�\���x�8��Ԟb�I��B�:���ݡyp/7��Pӫ�9nw�et��o�����`Yd�v����m�Z�LC�����W]k����7�� #3xK��Cs�v!�I���,��>A�����-���������m�� ��U\vg��W\2�['�k��3Ӛ
�0��P	�43ny�`T��9:�4���IQ���E	��&&��I$��"7���<��.A��?nŊY���؂�Ȃ����r�Y��{$c}�=�}�[��u ��D���y��bA'S�,V�e��}^PKm��܄�cON'�����������& P�����Q�Ճ���{�WFu���yr�x�_sm#,����QF!�ѭOǫ�@�u49�J�!��hI�0����}�e#;A�fh5&2ח-�ȕ�Gκ��� $6l��0��Bi��l��>��{��z�(����h3ٹ��#�Pp3�ZzX9�\}��h-������:,F����[��x���M��㋍!��W:J1�%↵�=I�z��TM`ڑ�^B��a�@���t����A����J��&a�>��%���h��B�?�`R�!����]Y�I���ۿ�|g:X�����u�}�n7�D1�V�$xH��-cFF%f�%��:�EB\�||�i��n���R;���l��������"�8�|�_n*v�|q�#xı1˜c}�|/׎���T�fx����7)��M�p0�����x$!�@ܜ������+�|�MBB�X|�+�"b�����_-	�Ը��/�wgh3)*�a	2��}��JMoZp>�
DG@���X X�s����4��@��� 	�I�-E�x1ϊ^�c����N��I|��o(#3�ꊷ&;�RTc��~�����ݙ6���X�ѠG�N�ت�m�E��w��s��`���K|� �]�v���(<�5���`/�H��tA],Kf%�"'(%̑9�r2#�!�~	��ʸ�i���L�#	mޒ.<$>��@�!\ˍ�r;_��0�9Vu�/�]�?�?2�$�p�m�x�H ��vX�8Vܯ_�9���/ ��Fc�A{�}w�������1�m��.
�H��GV�0�X�5n	�ԩ��^�d;�p�Z�Jv ��
@�#O�v��ug��!��닾X-��r�kַ�n�g��cd�Hu[ܭ��������?��r�Ƨ*L��#ac����<��⡣x�]e���%Ak�N	�g+�9:/���C <D�L�{�������Y�	A-�q�墯�.�,y� ��Iq.;����{��� ��Qh;k�Q���a��v�`�(�[�3}�u��	��}�h�"��0�,�}�B�~:�
b[>K����(dl+"�h��R������r9&+^T%�����(4��W���<5��`h�Hl��Iޫ�o?��xpѹ�>�Ǽw0c�(�7HT�~�֑�s� ��L��z{��bf#s���"y�F��:޾�)\��6��Q_z�(
f�eI&"6�n\����ߑ�c�_>�Ǭ��~L$���酝�����hJC���)(�e8B�-�A�#�������"��p�.�,<I�s��϶�]��i�x��G*�X,�Lت�O�����A��6��%n���O��0��������R߽��4��<Ft13~�&7�4�{�����@� t�MF�1e��b7��7!D�Һ��!D���"X��ID�h�|g�ĕmk�C��r\�%&K�Sى�d�+�$wu[�P�K� �z����*�5FWI�Je�߹Xta�$����� �N��_N��^�E{J
��N'5I�iC
T��^�.�4��)ۢ،�h}��a��3u���g���pV�_����'gzۍA�h�8o�:]�\�T�����5�֯s�g��(!?J�wr���U��Ǯ&x=���d�LN��lF��i^/������M��8�[��c¾���: q8�B�����b?��7���.t`�+���q]1)`c����18[hn;��^�����ЫS��NU�q���;��N\����G���X�D/�8���KcAɕYC����E�Y��JM��ˮ�9*�8�z��=W�T�7�����4ܙ�I��w�%�ׇy�O¹�QoB��6n��p��=A�����mY��5<�z]�'��,�c���Ee>r��+�ԙ�z�~�ͬ����#�ƨ�*'�Qr�U�.X���@��p��Z;�nAk���B��|�S��p�Ҕ��(,6W ��~�lD8$E{�;��R�!f'��3����	5^T����wa�H�P��oE�{i)c�н��Dw�:����զ&G� rq�� �[@�R��G��ߨ�ޓT�Y��v�!��F�`Z�)��1]v׮�G�c�^:���6z)���K��v4��<��ߙw�Bú��3����Vn�g�n_l؋������x�׎ ��i��27�\��*`6j�'A�h|�q�����H�[��4�V�UBL��L0�\���؆����3uz� xY�yxz�DD�N:{�nF6�sB��^������У� )�&G&��\	�nL��~ 1�����2<O��A<R����">&�i_5���,�t����%AWW��Ey�Bp��6�a����A�3B�&�dP<h7xy����
�37H��3`@߄�{7���AZp����I���}�Ю����7�!����*��½|�3�@������nJ���(��f��7`����X�K��LE�� `�g7%��Ќ����4i=+� ��-(�}YaVGSKH�Δxr�@u���g�_^�Y�ի��!Ͳ[+�P��A���
ǵ��l��
kǆ�d��ַ T�A��{$Z����ʓ5����\������^�A੆��l(ѵ���I��L�|hl2Շ��k#(���K1E��zjX��zU��:Ё��!WM?���	�f�� vW�����!�d��r G=tp���h�/@��;�o~_�QR�)#�	�}�T����h-X1&T�f��B(�N��Sҭ�R������_~C�Żߺ�ZF�����0��tf�I�#'�=H�la�{�"�d��>#�7X�o:K����^c#��;Y��_�����9 (r��>/D��\�B�����mIc����(8�d��J�lq�n;���X��������+�f,=F���=7$̤��jp��%��픯<���e�B�S"G�k_I���.?ֽ���byV�>h:�z�Ҁ�ٌ{�W���k��jY�eI�J�6��[��)��������5Rx���)�`����By�~%�&q�0m��+�H�R巿��S���ӟO?��0��_�0���k��W�[l~}��k+r�����*�U {�x�-]�=F�J�V�`��jp�/%�_�����D���J��3(z2�tX���8����^K.ކp�&/�{�J���M	��N�>�?,�6�(�x����H�H,۪m���aX۬��?F4ٖ��2���ֻ����
ηp��?`�R�n����2,@����1`x���UU��mmk' �R�+�.#T�ͷ!�Y�^�+P�
RO�J�����
,��Q�y��>,9����d*�*�yY�pK��p����oa8��H���W�g��4H�I�$����W�D��*�׼=�	�E�������{�z	�Xn�r���"� }^n�b�9���eP֪[���>�@8	��$Uf�D^��Ns?d���峤��50?�'6B}{@��9nv��H|eJ�	0�%����v,��M�#�`��J�%),��T�;�(uȿ���%�B��E�|�P�.�$Y����D�e&`�P�z)Y���#�P.u���7��k�����clG?�c�HS��zf��9�V#*�y��&�i ��l"_OK��� �`�ǯ����D�gH���Ý1�W��x�RNP�h�p/��B�A���2zDo�=8�o5N�cd�0P�49 ���8�#�b��р����G{�Y�nJoZ᢯����t�5�"� ��H)���"�,����vSb�Dd������g1���ΧV�$���(�00�L�c/�����+0��]�a�cL��F+ɔ�6#�q�T��B�A�X�O(�P�2� p��ߗ���U�쉆GC��@4m�T�:RWMc����eY~�ҫJ���y��#)�PM۽��ؠ#io7+dZD��8���/�,b��E@�oo�H-�E��G������P�Kq��F��|^��ӼO��@�l�-�/�Q}�a�~��	��[*�pK�q(d�pD1�ܝ���*�U�M� xe@�n�"��""���'Z~
d�cJ�:���6�`��^�� �׵nH<����J?��˖�$���ĵ8���ޤj�.��gd��)P|GrR}x�NM�;9i�{
g�Ig'�J��;M ���.SG�`�A��L�x�﫺s��� ?�	sm�2��YC��QYg7��@L�C�WB6#��z��a 7!B��C`�%D�:I�>{�X�JY��1��o��i�#+��"��= T������(��5�&z�W0 �t�e���Ǜ�w�/C�����x|�!��-I ���9���Y^_��lDY7ė�j�^ౖ���2��������c�咒�I��ob�t�Ȋ��&���6<#7̍�O�WK^�Z�Z�v�D���6Uชj]�{ٔw[ey)� B~��N���
~�}�hDkJ�h��T����гs8��wZ�8}Ή�O)b��mm?�b�H�V���;,f4\��x���&�p) �젮3l�e�U:�Q��yO�	-F����	�Z�v���wF���O;k�����hp6��(Hm��b���BYO�,&���T�c���4�hL���U�	�&Z�++Î�/k�s4���~ݲk�>ޥ��g�&��~r���%��#w{�RH�Q���S<������'Z�W����{�����dGM՞��0�)ܷ���|o�3շ�K+P��p9�}*s$�;U*�C..��DJ���'�[�U��J�]�x0��5zMϯ�ꦲ�m�	Ne�Ag���^����k���cR-����~z://U��,�41���S"�f�GH|�2m�Q�JMI�LՑ��� k\�QAd�͆:m w�v�:���C�������@�k�Y.�O�(��>]vf��	]��*$'�ꏓ{@�GJ��[�Ȇ��PBRϐ�f�`��쿀?������㛇m���ߦ����3Rpж ��|.�`�}U��e��	����7�s�[���]���L�<!�ěUx�ܿ�i�v�����ݢFX���#,a�]SV���(�p�Ǒܨ�:ǵ� ���C8m�R	Orak�������Y=����\K�^��fc���}��|܂�`R*(l����U�.�1��������Ǘ�κ(�|�0#�=��N�D���d�w�����PR�,o��ڈ���~�mr'����Ӊ�3+���Ƿ��Ϝv�;���}�s�lO3�8eo
�t��y����`����vrHS�!��r�����6/%��t���@ �@A��I��tu��>��z#96���[K��}�ud��l���wGL�:'��Y^��)o�͹�Ejt&׿�xeUK��B+F2�	���3$�qHE)����*c�3C��� ��X�:m�:�w�k��W���yn-�od�FTr�� B?0�$@�8���0�Zu�X|�H����""��I�<J���f���L�!kj)�w��M�8_^���	��*{��n��������ϫϱ-I�_���иiŚ�\���V���SȐ;C\��I�����w�-�.�ͷ��2l��W߆�Ov�������X"�ֱ�.���ST�C��I��]�Y�)��VEbb�[�ߠ>���A����H�V���V��%TzUr �HN`�{���?	S1?�P�~!�'lRI*Y+>��=^"�tf�*p^	�u��"���)Zf����|Ue#E�7�~�R��`��)� ?��c�K��-�q�M+�P=���,�9�'˷-�v�c�,r����Y�/'
�԰�o���������X�)�e����3��C��G��1)0S6��n����%�l˴��v�U�"�F-24#GL��
}�B�6�*��D�I]F���[�+6�8wG�"�"����!�:��wuu�/5Wv�I� c��s2}t��Q����WO`/&S�QN�:�v����2�N����=RBH�]��0��,c�.~��������C ��ӎ���kZ�����#knљ�\��.6ٸ�e[�H�ٯ�ɦY*�LuƮ���:����ӪR�5�~;fq:gt���X��L*p�+����D�!��]��P�J��p=�f�!��O�� �_�����X�g����S��6Y��j���XT]�/J��<��4�'p��o�s
��	N�W����*���R�Y�sF�|���c�}�Kd

Nf���n�\��%�Pr��Ҝ�RU�&v�+t�Z�1gm��Cu���i^���aK��-jarW ����R��q��k�T4�z�D���x�2 j/=Bm\�E�d���G�f�`��P�,��~�I�T�J%���y\�*;3�U��r��ji��BX�Ol�T6�	e�`/�E�T���ԯky�2��׬Q�t�}=��n�,mQ����M�� Y;2Z
�q���Y�����A�|sY�EM���iB����̖2�$�L��RX�4�Y&z�(�p�d�h$����21&��nv���r�k�y�!2Z��U����Ob�[wd@(W���N#O�T�6`�8�7�dk%��s��E!���<�8k�ky����'���"�X�!��O8c�Β��cJ���p�(6����J���ff�x5j{�]�,�.(��n�(7#!,�������!�/�玚Q���N�L��S#�+����`P����e���-�3ߝ�H�J쀾���iר��Oh�@���Pz�����g��,r4Q���<���r<�T���x�� ��N��j��z ��\���oU�����L�n~|4�$�*�x�{��|����i%��&�ZB���1��#��єͣ����ŋ�{<J�R�>	&�o�� �i"��u� �u����ѝ�څw^o��l�;r�?u�Xx��Gۍ�N��9I�>�8�r֑�Y�ܨ��,2�~���]3�ȅ�Y���y��}ZuKq��J�@7ɽ��a���;$�tZ�JkAPW��sټ���Z���,���ܶQaʾ�C2s#�e���Ic{��z�`[�z�G�����I����_m�^��K�tp�������X��Q�����LkǮB�)�B2��"�(����҅����_*�>���U��t^�{k�)�5M\�5��*�� %;��g��R:��ŋ��^�')5C�R�ލa|��
R��+2�>)�*��$�E�H��S��wH�%�͜�Z��MR=��>�a��C/�=h3���@��c���-�oXd��H��}M��'��.�Z��c�Ȓ� y�}�P�eO��� ���/�l�r(��+ؘ"�cgk��v�Cva�޹]}���>](�-S�7�a�e��8��i�)�>�b-H!R�gRx+�jӾ�7$4tW����	�*���pW3�s����� y؀�C8�1�E�X�l��_��P!}�b��-�㗆/���aSe������B�����V�a�uJ��G��Ě��ڹWb��l��^1��:��KVnۧ�Wֳ��Or����<��БomQ��j����ˤ@���~,�)\P��X���� �f�"��1�������I�8�C%
���Ҟ��o�6�7��3�#ռ�-�7� �=�cE�Z�$=?mzR�=ܫ":[��>��40�]���*Rc��
� =�W�M�aK�����MGB��&�M��ܿ��ln�����K&Q��<)҂��0e=�p��,-D,@u��{��ͻ3ӎ>��&��p=~����V��n@|4��'}t��W��)��#�^C8+�\ ����F7���~��jD�����ufǪ	����v�D7����{w0e\�BO-���u��d��dj�Ÿ�h!4������6u[X����Pg\,�5���l!_Mo�z��������o�-įڠ�o���a������dޛ'3�UE.8�L_�B2�PË�I=�lx�PB͔>� �S険d�T���,v���8��� ��Pt�����5'�����`\���p�0,����n=&��b��;rU-t�9k+��X/�X1���3<�	�&sp<H3���>pC�w~����eS����Q�e���𳿹F��]����υ�@4%ۦ?��L���0�9���oC�e'��O��^��}�aQ�X�d�cs+q!�D���Pn��u�BD�'��������}�Y?�Iq:~̤�5���c�\0��y��s:j �'�� ��9E�w¸iz���c���\���.ÏW�@@�qƻ�d�!)�,%�Pn��p8�|��W�@�(\������7�'�wZ�����e�l3��s���^f���%*[�MY���~+֤��.�O�y�M܄33�|�#�D���O���?�d;*�w3�늻�<D�p�	������]����MD)]nm
⿳��I�9쾒g�:e�K�v�(I%-S���3�5I��c"ݙ��W?�A�Q��['حz�b���A(?��P�io��_E�~�/Ƶ>�x��F,�c��hy�F	��M`5�1�cY`�J�	�Վ�u^K��E֎�a��ZX*����ulu7�y���q#C��.*'M����|whG�G}O>c�2|):�p��8�n���s=��Kv[�,@$��:�`��_F�l(02x8֋�8>)��;��_C�i�],�(I�'p}��iɦЗ�u�}��o��:��L����t�C��KI����+��L|�,���ЈV�F�C���9��l��^��A ����B��{	d*~sj�w�L�f���x���(�u�d~��6�5;M����M͘Z�,��&�Wy���{.�[U�ن���x��*���<���7�,-,: |OX���l`s�����x�[�� #��0�"ϟ�\����5p�^IaM&�c5᫇t$�u*�B�6���ȓ��� �:��+^�N�A���?���冈׬9���FH���O�.[t�R%BZ;1���"�A,�{�t3���k|��
"H�w�x6��5�Vu�~�g��H�Ȥ+'�m"�(���tF���B;4ҿ�j�0�e�����țVzc�P㨇��$���h��B��<h1{=��7�uU�i����鳒zG`�q�D(v6��ee��u�I��f���gB�2%�����3/�"���V�M��_�a`Q �x���Ф���r��j�]�>��gJ+�ӊ@��J���8���;s�R��<�V�<�����z��!�� �2�`X�M�J��6`:�ҟI������1�p�ԚrO����33���u�N�Lf����S�u]��i=�_xvv-hJO���#����$5��"�Jw��g_ck�	��wU�vo���^�^��x�?���[	���ة�,uG��N+xK�����56���#tw��#3�A^Ks�t�l�]�T�w�#�6�m�b�2"C�A��2j��y2Qɹ/,�+�_i���,)�t��!ʲP�=I)k��J����o���rtK��W���.m(�����V�Bc���DBf(x�ݮ�	��ՉɳF����8�sG@����s�r82��m*��Q>�j�G��2�)J.���W��M@�rlXM���v�5,��(�7��J|>�!�}�t���Bn��l(�0��w]#,P��8��ż�XCO|Cy����b���XmS�ϳ�a��v��]n��9����1�6�w+� cl�e�=�g�1�������15}[����O>j5�i����ů�|ñG��3_��鉡m��ˡ��~0QAO�0��fv-ޛ�om�W�Ϛ$x� |��9���+�p�H,;NZ�蛥��1�	�Y�~b�BE����j�1�~\�3"���������6\�)�����7��H�Bg���hS��l����E� $I�t=��Ջ���tf���ď�r��Md|Cco9���i�~Z�s6�qP�6LЇ���ú�<΃�x��k�<�f�O�������=�J0�Q입���k.�|أp%[�-Q�E���"��1��;� ��av��C�p�Q2��=�A�}��a:>\��i�UF��=B�.���G�rʻ�$z G�'�F =�[�X�.��~_I�n��+e԰O��;Sk��̚����2�F�p�\eP]a�$r&��8�^A��yPh�L�������G���d�v�m��=��5h��]�`qY�ձ��#�5�晜���+>���Y9���N���՚js�3��Kb:�IZ.�V�<�P#u�0�0����B6�V	9B-X�г1��L�*f���=(�j����T��pL]V�
Y�kX/&��Gp�ks���
�t�	ۣ� ��s/2B����O"��f���V�IfV��G��0��n�^!�@}���v���C�ݻȘ��Gt����a,*�����ቄ��b�}
�G��H�W ���\`�$��YE"��K��3���E�@�����5KR����Kz�h|c�.s��%�O�� ���"�Oi�t����E՞v��)�ܽ�@�".U.�0��Դ.�ל���Y��.�.2�	-#����2yf#�i�8��O�������X%�P����]�����wN[ۊH��$΍��f��a���d����Tvg��8Z�u����U�`h6��O۲��.�dτ��g��9UN�@X�+�D�,r烏�?MW����sDE?y����b��a���b����cO"_���@��Z�"��ʣܥ���(�y-bw�ڤ�wu _��8`R�!��ڼ.��gA��a��&d@�ߦv��F=��ѵ�y�d���Ŗ)ĥ:����2fI�'?#�bXU^�V]�+��K,�F
��&s5�9sk��܃���&��L���!�v.�  �Z
��	��2���'�U��G�̠�?(��r�'_��h�������=��0*�7,����-�p�w�O��5�Z��-��AO���D�L���p�"��G,�d�H�C���v�k:W�l-jD����>�U�ھr�>+��N�C�΁������X�7���$d{�s>�,n@�8�?���@Wrէ�,ܣU%�sE�F7�J
v��M܂��|�Š�t�뙌��~���Q�u�kC���;A-�q7m�p�.�	�tAs$C��O��m���IPaA���by�m��qfm�.�mP)��/w�k�41˓����SpM��V;��c�u����D]j��V���� �)��H&P���)� w_�q��{�������1�2��s��˟�E��o�f-��w)�bM�ֺW�%���5l-�~���a����������������_s�TY'�I%���p'`k6#MA���d�41�y�a�|�jN/2]�=�:unԨ7��Q��MAj���B�Qb�	߹�0�){Y �U|���[x>7��|dx�lo+�\�n���Y
GO)�34(�ط�c#�y��/�r3@жpL�X�����ͩ��BL\A�7 lB�̝�I��4iP��)��q�6s�D�ܢ2]{�4���j�y��0Q᳗��/tZķ�J0�-��|҄��!bUb��%�^�T{.~AQ^��m�lv(J����6	)��ke�j��4��6�j���7��F'bby/#�f����vR��!�����o�Y&�lfs~yãzl�K=�t|��	Kx�~��6�J�P��]�u_`%���H�t���YSi��:$yU�v��)孪�)�c�U_�.��Tz>ڝ���Tds�?x"n�q�4^�����/A�S�l���?w��>�+0�~���>&�n@�!���\�R~�r���f��P���HQ@�h������J�榛i�b���n�/�c3g^�>�'�����E������n�@i�ӒZ�j�VP}:�u*�������)��m�<G�[�.&$M^&��X��rck��.��s.����g�ފ$6�f$�-�j�5<[r�L),��0e{�
������e59�	����jy7�U���T���!k:��7�wr�%/%���"N< �;�:v`�$�ڂ ���$s���}���Gw94dl��Y\���6�z��+m��.¡��a�[���KB����d��1�fwJ��K��yv͸�J ����?0��z�������o�&�PD5�hϞN� w�0�࢘w�Is(V����m��"�검�
5�(�p���:�_��R��p���X��c"U��Ʀ"p{�Q��Ngo�}g��h �]n���N�-g	K���$$����g���)p�2�N���m9r���q��Su��+Y��?Άj\�tԻ���\ c��"���`���z��>���������1cD���ZI�����pu΁��o�
��c��5*vh�1��'����E�@"ƒgt�ԯ�*���"�iE����Yw]�+<�!"@P&����T���!i��.�,��6Ml�5���Q;�)��jŢ]>|Ē��Y��*��U����U�]7��֚}��+�V�묍HD��1����Lz4W�$0��J,C4�/]箛��ɝ��s[JǢ�&�.��S�65���)�b�	���>o�~��e�%&"BG�.Гץ&���j���P� ��سD\l�REf��p\Ŋ�����DQT�~�m\]?Dn��צ�Bp���ӈ�_�^}7]��>�+0���O����z��ڸ<�B"v3���	���4�BOk7�\`aĵ�J�����V}�y#�`��ad]cF�����/9�AN%�����u�������<¯�
��ٓ�v5}��y�w�+�����"�Z�R8�7��rՔ�}+~�O�ՑZ�QM�>�o},B2�7�:fuו��砑
�#~%W�x8�E�`V���rLm~w $�8��c�y��\����vOK�熭�M�0�S92N�)4����1�=߃�B�%�Mؘ�ߣ�Ȅ��D���n+|�5sw�,*��V���)q�$�]��7PO�͌4�l�A2�O�X�$��Uܧj�&���0�g���W-�ʂN��֡B��o�ҷ�U��	�M��u����+��,���V$zC�*r�$uyjpEs>bf�=��{�/{��t>��p�u窷�f�k%&��3��^�嘺�����u�̙D@f�:[�d:R�� �v~���	&F�4=�m �J�W-�^W�IT�v$w�^�Q��p�V��?F���=���\3��PW�������pg9��[�a+��4Wi4�u�6(OzB���o�uE�o(��=>�F9	�V&틲5��f�Y4��>���4^��S���"��2"0�VWOo�����T��f�W��OG0�OȂ�Pn7���<<�Ղ�)H����\��(~��#dD��
E�b;(���<_ؕ3��j�0'u o�����e9zc�$#@VR��(wz�@��n�?9`��56���@���N�UF�EM�N�����'�Ѭ�n�@����O�9�i7�ߤ�:�����bQ(o.�t5�%����'i��;�#Қ@�<�ݙ��ݘ�#�n���0N����9No��w5��������\�X4!�*�=<1`Y��4aK�ݮ
,"cZD�$4�|%���[O���[w#���
�og
}����檰�'('��]�h?y�!c�����Gr)��+`����Gn~D`�S%͜0��dOA֋Q⑂���%��,|�o�\Ta"ܛ�:cO{��� �)\��Q��k�	�nK9���ׯ�G�*���($��5ľ&�A��K��/���خEF����'X螵�7���U�P,'��ͬ3b|v@O^�(������oK�K)Y�H脺I��}M��� ��i89V��#��z�� �ioC�	��:(�#nL!�,��ߧs֩K@a���Ɗ��u֠��
Fڤ5C��������'L��1?C�|�ۓ�C�ù�ߒbw��a��ڰL�*f��a�'+�/����rn�
��@i�Qm���8b�>H�h���|�nOp�(�e���Q��w�c��7.�T�`4?E'x���rC���i��� w5fVYOH3��jp��e TƩ&,n���e�"*�4Ol}'FXd�� #��
 F%ԥK��&�'��_n���_>TΉm{lA�s����V�p4Wő�2�+B.��T_Z8�.�0/�*M���m��$�2��b�z�I)�_�x;�zw}"`�����3�u!�JQ��oN�]4�t���9��$�]�z����=Zx+�1{�^3ѽ�D�os�YE-�c4�m�Q#��W���a%���K�?��Y?h'�����X�L�*�fH^��Eo�]C5 n1h�nAt�}tSE���B��Cw�HR�l��{'�p�Q���ro,� )?`�Gv���o|��1�/]SQ�CQk��'d��?7D�~c W����v3_l�4��wM�i�x��ʷ�X��i������e,����(P�˘�'bkF��?Q&���P�)��؎�$�)���m��0��V$m��3EbM;����P�3�I��'X�A"}�*��T�����l6��)�
6J�������D�cB����rɈ���c+:��c����+)�����B�;0��nv�y�(�hj ����
k��G�F�R"�i��C��2\��#�9>���~b0�ՠUa7�����-i:�a�gX
$p#����)�@7'H+P �|���������<����}���d�K�!<�dD-/�l!���8��%v� ��U[�u����NY&#�I�7�lo0Z�&J���7^�͸���!��K����|�gs�'6p:�t�W�Aq<�[���r	��;�}����1�=�W6�A�CS,-��\�R�B��=����T����������"_��T��15���p���~4��V�E3/O'�%���p]��/��$xV�$%t�R������i5�6
���gr�d�jK�.9"2R�����P���Nz�5-Q��MD�w٬.�hs�>�nԬ�Q.�Z�<[&�Ε�O��qBS\��$�?�C���EDy�Y�X�0����&�2� ����p��C����t�+�~D�c.�k�w�9'T���XNs�}0�o���-�rG6�K�8�m V��V��\��>=�()/l�t��y�H3翷��#��%��P]�to�<#��Y�&M�V�}�	�֯Du=s��֠iԞ_��e�#���K�^Me�����띢L~��D�8S�I�?n�Y$�P5���"�͙;����������Hh�$��a6�"�K90����B���}�|�ysb!�7b\VoX���e�8�����.����M��8+JQ�~�����-���-�0qj6���(�q�SR�^n ����;���rx�wN�U�#K&��6='���L>�F!pm2��Q��V��A�漾x�V@[f���^Cq A:���|�5T����$tM�k�7Y��,?��?�&����h�{O��+��.���_�½kG�� \=Ш$����m d�Y��l����4�$�����X�P� a���&�*#u��[<�u5�����U��Ժb*gmڽ������n��|$�>�dlG7O��9������L�n���m��Vs��'���n�B�q�^���1Y|�!C�	��A=�p�=2T�;c0�Z˽�|&}u�f�R����
��
�� ��E��x��m%Q/�%'��f=COPV��F�ɇl����v��Ԅ?~%L��7���~l,�*��02�� ��L*Z�!�Іi���B$U�o�o� p�sO�F(`���o�41!���0����O�,������:�M��-E'�2���xH�r�2�p�4_r\b�s� �R]���B�]$sb/M�G00~/��edb��̥�2^Q�)1W��e�@�Q]v[���Q��h��-0Y���������Զ����N̎[Ǳ����߫�Y�������=%࡯m��۠Y�FˬOЎ}��
S�s�f��m���e�#���q�����ғ���`ԓIl����n�������H��b}0檆���"��{��s��o�
?��2��-����.^B�	g�������tC/Μ�{��"��|��E?��)�T{��Sϊ�m]��@B�
Qq
���:����Z4ԅ���i?:W/���~�I�5�=Z�+dT�H�� �#��2R������
�r<L�A(knӹ.s��VVShڸ����K��f���h;�HZE��!D�)U�'.C d6��B������f� �am��>y�AQ�0�!��L�����Rh�a�ݏ�:ċ*ƈ����~{ ��)r!B�5�
��=��0�A����5I�V���m.퇂�)x�fӽaC[��q	��%��at}�3�Ɯ�o������0\j}�p�-�X������0,&�n����ݘ�,���X�V�?G
D�<PG��&z����V�W��rGa�}e��'.\�_0�f�R����`#���M����\������Ťs����pu�+:�Z� b����v٫�`���W�U�oiF���:{~��щ"�D�X�s窄]���s��D �D���ەCE�C��;��ح��=��©u���K	���1f��D���$��"Z�t*�^h��^�Z2Bn/NU�G)�Ra*��:�6��������m����!b��B۾o䦂n��Uĵ���X6���:��ۃ��Av�o<��Iq�<��lٲ��g�ҭ,�-�}����ax�Ж?, �A$|�MQ�VIq����н���hcR�6���;��	i!DԒ�BYͅ}�>�p�iC�K�l�6§g�(��$��aDd4]5Ԓn[�{��9�שCk��`����ꉏq����hS�C��(Q{�K2�_(�X�� ��kUN��7�W5�O�ao�#WFf��՞�s*���ŰBL��<@�vҧ�`�j�/�w�2��Ӥ�Q�JQ����-l>���S�Q0���j�$��q����_;�O�'����jg��gɻw�_�Q�1qƪG���h ���T��'���cRT7E� #+G	�-���V��VQPD�պ�}�D:��im��}J)B�fka��E1s�t�Q��W5�DBL㩣�镰0�9��z8���A:�Tf�U��Ա`���HX�N?V f�!%�T����ǥ���kx%���0��,3��԰D/�S���Z�X����K[	t=q7W�I��̠P"nM2����o4� �����W?�e$c|Z4����UE��+Q�h�ֶ���ش�q���;�I��:v�~6��\�~_W�G�'/fX��X�116�&w���~�k�%���?3����Q��%6�����l=�7�v:xx�&�����uxb��9������RX'�/��3C�ޥ��:"�c�X�r���c��k�m�+�]-�a/��ҿ"����_*(i�~ǿ����M|��c����	�HW����Â�t�sq.���bBJ5̼i2Ta6�É3Ȅ؟^���n��P��61P�����a>V�j����+�'��U � n:!&K͹�*�s9��JD��K@�B!�:�x�W��yt��ɪR����z�H�ےL�ٳ�����씷`����84�z\�����XlF/Q~�w䧀��XaSV>Pwܲ��>(�e�>
�D.��dujS�6�ff)�G���<9%��[n�? �X�pg�}M���
&�u^F8�@�wց&�9����,�5J�vZ����IS���o'Ϗ�$�I�)�ݷoS��߾)�rE{���a,Y@ B��e�&+1�я�Z�2U����1�)����#�d닋��Y���I��9l�C[��d�d����pM��䌷�}f_*� ���5g
�'�;Uvfw�E�	���a�P(eFe&vOQ��,� %�/�}6�0D�55�onq�aМ�3������ʕ�Rbms��u���T�^*>�o�l����\�J���m��S
������9	�����'D�#��B�{����REQ�Pa���i����j�K���$x����M�s3!���Fȑ]
 �MqӿKd����
� �k�;u�p�mӬ�Y���������s��ʯW�Hƌl�bYŖ�V�{m�N^�N(���"[�/� �^��+���*sN�&e	�*'��T:B�d��+[�����S��i~�)�(��T
j��.3H�ڤXE[.�k��;�5�A;ށ��daYV.�%ؠ���1=�č�BDч��]������vR ħkv�2[	��8��d(]�a?�ir����5�A��{�Q�2��}6?��#�&��N��Ή�_G(-�at�����в��!,D���
�����fGw&6	��/�D��o'$���rͱ�kk�\y���۽`�C�3{k�3p�cGq�E9���n����ۭ��Qma?�MѲ���:���y����jI�jѱ��1?7j�����l���tn0],d�����-�o�&_F��+U�>�0�m~,�AF�<��s�%��IUz=X�+��"G$�V
:�f��$��1fI�W����
�]S ��Ѯ������/!ݱny�
fb��R����d�}���-�-m��s�T�6��7��$���W�C]�k������5����Yrs�� �\n���0���0��������׵]H;�Y����6|�k�z����(x�5�:ԁ=pi1�`*j�7Lx�1���� 6U�uZr"r4��x?�i�"SA�Bc���������I��r���Y6�� e�:�Ա�iջ���K�|���@7�
���3]���M�^7%�sI��fAHݗ�^ln�t�����
���R�.V4�\!��=������>���O;K"�3jΟ�a,�Z�@#�m$��7:�I��-�4��3FA� ���V8��E	�|S{��k ��j���s	s�>�p��~��9��� �1���ls�,�0�0�J�A����5Ui��]�=��vP۽�z�?=��eĨ>��>:L"Ou�Cr&�{�R�ޒ����V<�/oG�Q`���j��� �{u��
�D0kء�e9V�j�:Oۯ32�(��/�+|Ù��58�f�POB&�t��uVl+�K/�"�<X<=�$�$�������ר��Iҫf8zD�P2�ل�î��Lj˟���b�Χ؜>����_�������="��?J}�J��*��� Z���-����עD����� ��3U�M�����ܽ
<�6p����=�)�U֒ƭ.l���.s�����=�	�ni�g��N�?��AF2�Vm����	P�:4�ؗ�k�D2�P���[�xٔԟ�\�hf0��"�Otq� �38Ϥ�L"�h#U��b`��
����D{w��cp�A4��}��u��/7�^4)%♯7Vcp9���Do{G
�@y�@$�
��K7����;�6�x��})�6�'�p?�%�?9�F��0#߱�Y!̓��gl]4���2���CN6m�\c�#�`�5�E�4���v�٦D+t [Zy��w�������V|��4P��cR�z@���i�stA��i���>��w��P�q���ڤQ����j�(�c��!7���`u> K�mWx���+�t�1�P�<y�� 7��ޯ�����P�f��}�%�W��"�ʚ����6P0=�_��(���o���Ԫ��@���F=�7޶at,�춶���up��)dd�L�=�i��fOc	DH�z���_�(�
�����1#i���g��C����IG+��2;�ԛur��i��*�L�N'��<���~L�hy?���]���V��Ɵ�s��2Ft��5�#��t`��|��y�.�����p�+����v$��7�ۣ{�/�GŝՖ�@,�LAgG����d���M��0Yd�sP6�M9�On��]���rn�30m�v�Iq>�Vy�w7��'���0�\�}�M�8�z_�ӽb��K�Q����Tw�x�z�&�����2���M��l>� J���xi��h�)A�%�D�"���O����>�ۡi;�Q��s`��׀�G��4��C2�C��-i]נ
�.x�'<)��<��H��zl�禮@|�� ��=G��M�O�{�Ԥ7�R�W��2T3j@�T2^:������L�ne#t�Y��ov�6������㍬���]�D�*�wnV��.�; �\@	�մvc�)�������{�Qd1��Bm%x�,0����j�8�4=���uN��ESyo�Bg��QB�\is����Ⱥ��mpp�n�D�p~��Ibb��p��_O���%��JI�G�+�ɥ�rh�H��@���d�&��s�U�C]X�^�h�|iA�t�V�d��5���<��ާ$�s3H�<�)�+�ERе���S%��?PTH7?�X*�b$shm3�ٖ�� �.�븤��*�b�r �b�@�N�ϲ���8C=���.���4M)�మq��*V}��h:O �����A^P�@J_�{��!�NT��z6����jv�e�L,5-~A'k��v@_�UE	���dS�n�����	�<�H���X������|����R��>���Q��%}�jL�@�f�	2s^F��9������t�Qkʡ�/�^n�cxO.�1t��݂�:�A��%]�ͽD��`|��]�KȘlK6�	6J��v;�Na�a6��W��j\�!�Bjn�W'_W��&`r�EA:�}1У�1���*	,�3=�0���b3]g˕Ur��&�%n�Kh�븃K�s�j??}���e�2�1A�m�D�a�1������n$?�^�Y+��Ǽ��ᧈw@�JU&
�!ؾ�7���R�u�9=x��' �y٢�A.��W(�c�"^��S�4l��S����#�#Ūt�/_�m���X�U�/��9�v?-�)��qSyg�K�,�(����$e���s�!�*�&��[(s뵛nQ�Vd�C"� ���y���j�݊����\܅�%�Z�������
�Au]f�ˋ��;�U|�To�H D��W���9.wK#V�_-X��_M�k�0��)�3�v1cmy�C���[�qV��ۅ:��0�,�.^����� n�	�tg�9ihe�v�q&�r]c���7����|WN�������>�pn��Ү���;V�p�ϒ&�vto4�~*#����2���ab�5\sBǣ�_��]L�d��,3��b%����#٦M�]��>�h���,���$h���"��K��X���1����X�}�%��o����0�M��H�Le�y"VTj����|(����/Zs� ��=$��Rҽ��ʸ�x.顂���q� �K�������Ћ��h����V�M1�
��8n�G�0�m��Q"��
2 0���[��oi[(ּ�}��1^Sݠ��o�D-|h%�Z���0�fL/�Z�b*b��Ű~>����i�f�F%��p}�f�=�8P��M	��M����r\�ś�+�D�(V�@ⲿ��ɂ�t�$��;����Yt<5�d�e-2ħ �~1�?��W������*�]9-]���\»�?�r�a����P?�]�9]J��"�n7��ʋ���q-�K14���XT#�<����g��+Js�T|��K�	�9 -�h����[��;��`���0FJp�jw�w��c�H��J����
���r��3���Y>-��&ִ"!�,,R��A�Tc�Z�����2;�� 8M����D��	I)(�3v����"�s� b�I�۶��ޘ��sJ �ϯ�D-H`؏>��+�����r���YD�Wj�a���z�mRȰf�TZ_6ē
1�S 0�1��^����=!΃�~��J?~�+���_��#��NlH��Lp<�^ɎŒ`��_�CO������w�Х�`�.�o&��@��m$����O��~=�f�u��-�n<f��U�w	�	��5��n�����<�ʾ��K6���4�n�(ou��)'R����%��3��� ��	!�6a��R�v0�7
�O}�N`5�}�B�E��7�M�ɋC;�?�Y� �����4<C��t-��~m�=��,wh�~-���2"$����o��s�����C�jl,h�F�����`\�ݭ�>�|c�a�Uˠ����2�5�[���Ss�î�x 8{'U&2�"��=��u�ce����8��ѽ�ڨ_��� � t�����D-~g�X���~ǆ�J����Lʘ�v2�OsS��ҵ���n]hҷk��ϯ�r���Z�y+�V�}�}�Z38W�H~�	��3��}���QJR�g����~]��e��G����s��L�bRHC��Cl�PV��B�؄�QɬD�� ��q[�s����F&5�(R��b!�$G��W��7/شVO�.3Tpƕx��:12b)�@Ar�
���
ߗ��^�
Cl�c��Jm�j~fU���=�E�TftV.���ƹ�%''���6����R2�,��23���&En����Zk���xD!�
��i�v���#�lْ$t�Is 곅w�MZ����zޭY.�B
��{�r��-��~!W�$7�S@V�ŇDK�Т�wӃN��䴇]ֽVW�dC�H��?/,��I�8��ñ��=����:�J�>���P__��6�YS4
�}>��k����ڃt���fhUSQ��n���.���L>��@XlI�Х
��Fu�o1� i�[�3]H����0�Aċd"�#n��@4P�0Q� �'���q9���j�]�G��:v�ȷ�{D����F�G �Z��W ġ��!
�.��$�2VT�H��~��4\�y�ɼ�Y�ľ�l���Dߛ���!�uS���^.s�~���&�T�b;�.�����7�B�/ܐ���{S�����-3��p�{z�<���I�2�����xq�OyW��MT��c���*��b:��X��fΖ��,M�KV�鴫�H���N;拣t��U�a�Pt�a���h�)P	��	��x;�8@(����M��]��j�~��F�M��l+��i��� UA��0�����k��")[��s�*E�x����z]F�&B�wIY6]�x�3�$��ܛ�����!�\e&(Qe{���L������Q^K���!��6�u; ��d�"c�8�	��ܷ��\|��#X���[&��Y]	NA������ �ª%VZ2P��
J(OS�()yH��:�7���T��%���TcJ�F�H�&��v�AALiRƷ'Bڝ/�	���(٨˩�fҎ$��}�DKBq-	],�$�6���}?�2V����a�	���s,��:���C��R�cɹ��8�K[*a��2A��Ro\�C�N�'�8���?9�a�4���R��[�T�v�}s�y��
�)�'���[� 0�Jk�hei*���.�J�99�({�QC�c��}t��� ��V�%�|�,Yhj�ŶOq�k��fs�q�f�������*Eʏ���}X3!��T1��͂�K��z��{'`S8�[�#�q�\��DGr�<Eb�3c`��2��/�UAXP�$/|rn�C�}��0�);���M�Aem0�u��3k��Uã��������:��9�s�U����N9;�����~;l�!�����%��
Li�@5��1&��'�9�g��}\�i�A�����Fߝm���R��3p���r�^-�Hc�gat��M��^���>[UDMÒ����m�;�U9���iu�(�$��d�Vm|I��1���t�8����q��3�\��8L"��Ɣ�����@2O{ ��[p1"���o����qWr	.<!%j��R��F�K�����Жn������*gKW�2�\��X�
� �z�ĭ�ϸTw(=�CdO^Nb��
ʠԐ8�����/�2]�P<vֆ�S�1j\���(�������<3ii6�Jb��K�m]���
S1���p�Ď^u�I<�k�8<���:�u���#|ÏUX+���+6c�ʈ�s�'�<D=G�f�-Ot�����v�vF��jf s���i�h$�X�
����!~�5�c~��eu~Q��Qp6��\%ut��8[��&����F�^=�1�J���xS���W���V�܀-f<Cq�ۗ>��XN�]��˓�M������5,���Zj��עTe���o_��2���٪ռh��Ku�~R"}m��ez�G���n����t�˘� Nȹ[凑N��V-4��7��
��*1�G,m;WU�	ׯ��U���b����Pc�@
軑H*�������f6����Q�'�d���I��h���2�����ITeh��E�Gt�E	��>��W����M7��+t�	�lHC�RdOy|䛭q,z]exd���>���m ١��4=�>��2.>i���[��k?�;�C��ظ�U�V�"V��j��GҚ$���\���/�j����T�@�fz P��Vnޑ�Q1�iy�#6�G�>������k�ݿ:��\�ł ��F�l��&/<4��[oJ���&~��i��3���2��f��"h��V���~�������2��[J�X���d�.	��Z���s��O��X�A�����,L�v������m��V�-��ަx���s]��ݑ��:}�SP
��\$�o�m�P��+Q`d��^�cC3Vs2A�p0VOH�H�Տni���}�����U�`�Wx�-R 9�eVq��d���i��q�u�Jd�-��z|�(�C�A���5���Qq��Q�nk��Y��"����[4l/H��`��� �#Cנּ{:6*ȇ�{�b�4q�XU���/Uu+ۥ��fu\WܯK]��ş�+e��w�.��9-��a=�c�Ä���4є�qR�|�4N�LX1�4�Đ���>�;�Է��bA�u7�1h.�W�H%���JvJ�[X-u�D��#w��B�>.U��e߭�?���i?���
�$|-�ؠ{�ᨻ�0��*����KJ���z�9�{�x��>2=��[������5\�1�1fد�3�O�E�Jb����!�	��N�J"�k�>��w��n��y!�Pa��}d�r�<���۝�� Y^D"T��7�Z��?@��ޣV��±��3d�%=��raS���G�ᆖ���,7{R�ղ�[�1�t������0|�0<d���� L���p�+���6�0��E�9��怋b������_��h�����g��.�/O\�P6�]QoN�aU˵��\]�$g*�=Vk�B���O�{
(N����<�f	Pi��k�:�R�����4�YvO�� Zquu�8/G�e��y���MM�k�xǖ���3&���Wc)�!>��	;���xb#C���T��&*?�W�W#�������E�;���L6!�X۪+��5dPu�B���cY�v��xQ����L�����j���ȟ�s=zۈ��k�?!Q5m�᥋�o'gb��h�:z�(�aB��f	~������X�>c��h���i�F-�؟B3ز�we
�3�1���U�� �y�Rب\E�M�腝=#{y�ki+B�k\�I��; �*��#����e�_� �Y��'�P�?���Ֆ�S���'��xRo�/�bYbI.|����N�Ū�ă�3t���$D�P��^Mzj�c1�"�<k>��v���%{Z�XK�p��������h�T��/V �P��qNc�]H.�z�0µ�����y���܎�K:vޒE/=ۢH�2 @��Ԟv�f@к��wr�l�]g=M�4F즰��c��L�)���y��a[����L)�Y6��{���I|O��ޢ�w�7[n�=��@rT*
����!no!z���D�=⺚��o2�\t�b�#�j����!~t�t<�T��[�7�	�DP�n-�]<�i�e	h��|��?��U�ǠT�:;<�I�ԙa���Z:�q�oQ-��2oz�Y$�Cj����RZ�L�;'��г��e$Q1��.(X��|&�QvA ���=�0A�zgD�aA`%���p�˱�Y7�%�X�],1Jh}�'�[�oQ b�oA>�~:n��$t�)�cL�F}.�c?o���$[b�Gb�O4Q�"$e1�T��21�ʉ��O^��>��n�l��v�u{��xf�}4��<~�D�T(�i�W� ����뭫�;�';٭��̑�p���_h��$�'�R��)J�E�`B<��1}��䑆S�~`B����G=�fwoØq�l�4;���nAm���Ie<�)0A���c�U�!ƣ��������U���H��oqC�O��;��Hl"���]�w����\s���þN��,r5����ƵБ�1sV��p�Ɏ�낲��R0��XG��O�qy�q;��Gk[b?�u�;�E�bC2�ڤd)�_>��* �5�/,YB�eE��5����:W���� +� ��/�2_��$u���������\����e�+'y�n��R���2�߹�A/��K�����mNᒯ��-��M#+�킛��Z���S"� ��ݐOw5�}�@�bWBd�������-�]P�/AJ5�����O�Ī� �3<�{�4e|���-��d�S���3�f �*7?�����	 �VT�`��ӓ��ǂG���hIK@�67���9�{/]�/u ި'��Cyq�g^��-b�S�V�[#ӌv��=2\Ϡ��۟�(�@!�9�N��D`�#�.���&y�p�����WH�0���9���������Z�5��#�����c�s�nd�$��X��/��%�@ͅ�t[����a)���<�_���FǯW�&1���ǒd�%*"��S܈�̺�w=Y���Db��L��l��w�.pz���h����؞�㫬i�Id��}��h�ݭ$ �6��m�yvZ�|�����&͜���Ɉq*]?n:+�f��p�6��v��NŹ*�9��B�ynzhW�+E��_Lz���U�����B?�W���f�t���ѐ�/���0���~��wl3��40� �c�ŕ��,Ɣ+#Ev&���ݙ/���P�ap��b>{&�
�Fo�ؗ���F>3���X��6�u��uem9�t2�aR��cS.X��O')R%���ƫ���v�&n�]U!+:f��*�x�ɼB�GL�涢��